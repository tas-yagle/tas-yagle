* Spice description of ram8x256
* Spice driver version 700
* Date ( dd/mm/yyyy hh:mm:ss ): 12/09/2002 at 10:13:36

* INTERF write vss vdd en dout[7] dout[6] dout[5] dout[4] dout[3] dout[2] 
* INTERF dout[1] dout[0] ck adr[7] adr[6] adr[5] adr[4] adr[3] adr[2] adr[1] 
* INTERF adr[0] 


.subckt ram8x256 5181 5182 5183 5184 5185 5186 5187 5188 5189 5190 5191 5192 
+ 5193 5194 5195 5196 5197 5198 5199 5200 5201 
* net 1 = mbk_sig201 
* net 2 = mbk_sig211 
* net 3 = mbk_sig219 
* net 4 = mbk_sig220 
* net 5 = mbk_sig132 
* net 6 = mbk_sig157 
* net 7 = mbk_sig192 
* net 8 = mbk_sig1 
* net 9 = mbk_sig3 
* net 10 = mbk_sig204 
* net 11 = mbk_sig212 
* net 12 = mbk_sig222 
* net 13 = mbk_sig221 
* net 14 = mbk_sig135 
* net 15 = mbk_sig159 
* net 16 = mbk_sig193 
* net 17 = mbk_sig9 
* net 18 = mbk_sig10 
* net 19 = mbk_sig205 
* net 20 = mbk_sig213 
* net 21 = mbk_sig223 
* net 22 = mbk_sig224 
* net 23 = mbk_sig136 
* net 24 = mbk_sig161 
* net 25 = mbk_sig194 
* net 26 = mbk_sig13 
* net 27 = mbk_sig15 
* net 28 = mbk_sig206 
* net 29 = mbk_sig214 
* net 30 = mbk_sig226 
* net 31 = mbk_sig225 
* net 32 = mbk_sig139 
* net 33 = mbk_sig163 
* net 34 = mbk_sig195 
* net 35 = mbk_sig19 
* net 36 = mbk_sig21 
* net 37 = mbk_sig5200 
* net 38 = mbk_sig5197 
* net 39 = mbk_sig5084 
* net 40 = mbk_sig5083 
* net 41 = mbk_sig5082 
* net 42 = mbk_sig5081 
* net 43 = mbk_sig5140 
* net 44 = mbk_sig5139 
* net 45 = mbk_sig5177 
* net 46 = mbk_sig5176 
* net 47 = mbk_sig5137 
* net 48 = mbk_sig5077 
* net 49 = mbk_sig5076 
* net 50 = mbk_sig4904 
* net 51 = mbk_sig4905 
* net 52 = mbk_sig4945 
* net 53 = mbk_sig4946 
* net 54 = mbk_sig4985 
* net 55 = mbk_sig4986 
* net 56 = mbk_sig5022 
* net 57 = mbk_sig5021 
* net 58 = mbk_sig4983 
* net 59 = mbk_sig4941 
* net 60 = mbk_sig4943 
* net 61 = mbk_sig4750 
* net 62 = mbk_sig4751 
* net 63 = mbk_sig4791 
* net 64 = mbk_sig4792 
* net 65 = mbk_sig4848 
* net 66 = mbk_sig4847 
* net 67 = mbk_sig4903 
* net 68 = mbk_sig4849 
* net 69 = mbk_sig4845 
* net 70 = mbk_sig4788 
* net 71 = mbk_sig4789 
* net 72 = mbk_sig4617 
* net 73 = mbk_sig4615 
* net 74 = mbk_sig4675 
* net 75 = mbk_sig4616 
* net 76 = mbk_sig4674 
* net 77 = mbk_sig4673 
* net 78 = mbk_sig4711 
* net 79 = mbk_sig4712 
* net 80 = mbk_sig4670 
* net 81 = mbk_sig4671 
* net 82 = mbk_sig4611 
* net 83 = mbk_sig4438 
* net 84 = mbk_sig4481 
* net 85 = mbk_sig4480 
* net 86 = mbk_sig4479 
* net 87 = mbk_sig4521 
* net 88 = mbk_sig4520 
* net 89 = mbk_sig4556 
* net 90 = mbk_sig4557 
* net 91 = mbk_sig4518 
* net 92 = mbk_sig4475 
* net 93 = mbk_sig4477 
* net 94 = mbk_sig4285 
* net 95 = mbk_sig4284 
* net 96 = mbk_sig4326 
* net 97 = mbk_sig4327 
* net 98 = mbk_sig4382 
* net 99 = mbk_sig4381 
* net 100 = mbk_sig4437 
* net 101 = mbk_sig4436 
* net 102 = mbk_sig4379 
* net 103 = mbk_sig4322 
* net 104 = mbk_sig4324 
* net 105 = mbk_sig4133 
* net 106 = mbk_sig4132 
* net 107 = mbk_sig4189 
* net 108 = mbk_sig4188 
* net 109 = mbk_sig4245 
* net 110 = mbk_sig4190 
* net 111 = mbk_sig4246 
* net 112 = mbk_sig4247 
* net 113 = mbk_sig4243 
* net 114 = mbk_sig4186 
* net 115 = mbk_sig4187 
* net 116 = mbk_sig4015 
* net 117 = mbk_sig4016 
* net 118 = mbk_sig4013 
* net 119 = mbk_sig4014 
* net 120 = mbk_sig4055 
* net 121 = mbk_sig4054 
* net 122 = mbk_sig4092 
* net 123 = mbk_sig4091 
* net 124 = mbk_sig4052 
* net 125 = mbk_sig4009 
* net 126 = mbk_sig4011 
* net 127 = mbk_sig3820 
* net 128 = mbk_sig3819 
* net 129 = mbk_sig3861 
* net 130 = mbk_sig3860 
* net 131 = mbk_sig3901 
* net 132 = mbk_sig3900 
* net 133 = mbk_sig3956 
* net 134 = mbk_sig3955 
* net 135 = mbk_sig3898 
* net 136 = mbk_sig3856 
* net 137 = mbk_sig3858 
* net 138 = mbk_sig3666 
* net 139 = mbk_sig3667 
* net 140 = mbk_sig3724 
* net 141 = mbk_sig3723 
* net 142 = mbk_sig3781 
* net 143 = mbk_sig3780 
* net 144 = mbk_sig3779 
* net 145 = mbk_sig3782 
* net 146 = mbk_sig3777 
* net 147 = mbk_sig3721 
* net 148 = mbk_sig3722 
* net 149 = mbk_sig3535 
* net 150 = mbk_sig3534 
* net 151 = mbk_sig3533 
* net 152 = mbk_sig3532 
* net 153 = mbk_sig3589 
* net 154 = mbk_sig3590 
* net 155 = mbk_sig3627 
* net 156 = mbk_sig3626 
* net 157 = mbk_sig3587 
* net 158 = mbk_sig3529 
* net 159 = mbk_sig3528 
* net 160 = mbk_sig3354 
* net 161 = mbk_sig3355 
* net 162 = mbk_sig3395 
* net 163 = mbk_sig3396 
* net 164 = mbk_sig3435 
* net 165 = mbk_sig3436 
* net 166 = mbk_sig3474 
* net 167 = mbk_sig3473 
* net 168 = mbk_sig3433 
* net 169 = mbk_sig3391 
* net 170 = mbk_sig3393 
* net 171 = mbk_sig3200 
* net 172 = mbk_sig3201 
* net 173 = mbk_sig3241 
* net 174 = mbk_sig3242 
* net 175 = mbk_sig3298 
* net 176 = mbk_sig3297 
* net 177 = mbk_sig3353 
* net 178 = mbk_sig3299 
* net 179 = mbk_sig3295 
* net 180 = mbk_sig3238 
* net 181 = mbk_sig3239 
* net 182 = mbk_sig3067 
* net 183 = mbk_sig3065 
* net 184 = mbk_sig3125 
* net 185 = mbk_sig3066 
* net 186 = mbk_sig3124 
* net 187 = mbk_sig3123 
* net 188 = mbk_sig3161 
* net 189 = mbk_sig3162 
* net 190 = mbk_sig3120 
* net 191 = mbk_sig3121 
* net 192 = mbk_sig3061 
* net 193 = mbk_sig2889 
* net 194 = mbk_sig2931 
* net 195 = mbk_sig2929 
* net 196 = mbk_sig2930 
* net 197 = mbk_sig2971 
* net 198 = mbk_sig2970 
* net 199 = mbk_sig3006 
* net 200 = mbk_sig3007 
* net 201 = mbk_sig2968 
* net 202 = mbk_sig2925 
* net 203 = mbk_sig2927 
* net 204 = mbk_sig2735 
* net 205 = mbk_sig2734 
* net 206 = mbk_sig2776 
* net 207 = mbk_sig2777 
* net 208 = mbk_sig2833 
* net 209 = mbk_sig2832 
* net 210 = mbk_sig2888 
* net 211 = mbk_sig2887 
* net 212 = mbk_sig2830 
* net 213 = mbk_sig2772 
* net 214 = mbk_sig2774 
* net 215 = mbk_sig2583 
* net 216 = mbk_sig2582 
* net 217 = mbk_sig2639 
* net 218 = mbk_sig2638 
* net 219 = mbk_sig2695 
* net 220 = mbk_sig2640 
* net 221 = mbk_sig2696 
* net 222 = mbk_sig2697 
* net 223 = mbk_sig2693 
* net 224 = mbk_sig2637 
* net 225 = mbk_sig2636 
* net 226 = mbk_sig2465 
* net 227 = mbk_sig2466 
* net 228 = mbk_sig2464 
* net 229 = mbk_sig2463 
* net 230 = mbk_sig2505 
* net 231 = mbk_sig2504 
* net 232 = mbk_sig2541 
* net 233 = mbk_sig2542 
* net 234 = mbk_sig2502 
* net 235 = mbk_sig2459 
* net 236 = mbk_sig2461 
* net 237 = mbk_sig2270 
* net 238 = mbk_sig2269 
* net 239 = mbk_sig2311 
* net 240 = mbk_sig2310 
* net 241 = mbk_sig2351 
* net 242 = mbk_sig2350 
* net 243 = mbk_sig2406 
* net 244 = mbk_sig2405 
* net 245 = mbk_sig2348 
* net 246 = mbk_sig2306 
* net 247 = mbk_sig2308 
* net 248 = mbk_sig2116 
* net 249 = mbk_sig2117 
* net 250 = mbk_sig2174 
* net 251 = mbk_sig2173 
* net 252 = mbk_sig2231 
* net 253 = mbk_sig2230 
* net 254 = mbk_sig2229 
* net 255 = mbk_sig2232 
* net 256 = mbk_sig2227 
* net 257 = mbk_sig2172 
* net 258 = mbk_sig2171 
* net 259 = mbk_sig1985 
* net 260 = mbk_sig1984 
* net 261 = mbk_sig1983 
* net 262 = mbk_sig1982 
* net 263 = mbk_sig2039 
* net 264 = mbk_sig2040 
* net 265 = mbk_sig2077 
* net 266 = mbk_sig2076 
* net 267 = mbk_sig2037 
* net 268 = mbk_sig1979 
* net 269 = mbk_sig1978 
* net 270 = mbk_sig1804 
* net 271 = mbk_sig1805 
* net 272 = mbk_sig1845 
* net 273 = mbk_sig1846 
* net 274 = mbk_sig1885 
* net 275 = mbk_sig1886 
* net 276 = mbk_sig1924 
* net 277 = mbk_sig1923 
* net 278 = mbk_sig1883 
* net 279 = mbk_sig1841 
* net 280 = mbk_sig1843 
* net 281 = mbk_sig1650 
* net 282 = mbk_sig1651 
* net 283 = mbk_sig1692 
* net 284 = mbk_sig1691 
* net 285 = mbk_sig1748 
* net 286 = mbk_sig1747 
* net 287 = mbk_sig1803 
* net 288 = mbk_sig1749 
* net 289 = mbk_sig1745 
* net 290 = mbk_sig1688 
* net 291 = mbk_sig1689 
* net 292 = mbk_sig1517 
* net 293 = mbk_sig1515 
* net 294 = mbk_sig1575 
* net 295 = mbk_sig1516 
* net 296 = mbk_sig1574 
* net 297 = mbk_sig1573 
* net 298 = mbk_sig1611 
* net 299 = mbk_sig1612 
* net 300 = mbk_sig1570 
* net 301 = mbk_sig1571 
* net 302 = mbk_sig1511 
* net 303 = mbk_sig1339 
* net 304 = mbk_sig1340 
* net 305 = mbk_sig1380 
* net 306 = mbk_sig1381 
* net 307 = mbk_sig1420 
* net 308 = mbk_sig1421 
* net 309 = mbk_sig1456 
* net 310 = mbk_sig1457 
* net 311 = mbk_sig1418 
* net 312 = mbk_sig1376 
* net 313 = mbk_sig1378 
* net 314 = mbk_sig1185 
* net 315 = mbk_sig1184 
* net 316 = mbk_sig1226 
* net 317 = mbk_sig1227 
* net 318 = mbk_sig1283 
* net 319 = mbk_sig1282 
* net 320 = mbk_sig1338 
* net 321 = mbk_sig1337 
* net 322 = mbk_sig1280 
* net 323 = mbk_sig1222 
* net 324 = mbk_sig1224 
* net 325 = mbk_sig1033 
* net 326 = mbk_sig1032 
* net 327 = mbk_sig1089 
* net 328 = mbk_sig1088 
* net 329 = mbk_sig1145 
* net 330 = mbk_sig1090 
* net 331 = mbk_sig1146 
* net 332 = mbk_sig1147 
* net 333 = mbk_sig1143 
* net 334 = mbk_sig1087 
* net 335 = mbk_sig1086 
* net 336 = mbk_sig857 
* net 337 = mbk_sig916 
* net 338 = mbk_sig915 
* net 339 = mbk_sig914 
* net 340 = mbk_sig955 
* net 341 = mbk_sig954 
* net 342 = mbk_sig991 
* net 343 = mbk_sig992 
* net 344 = mbk_sig952 
* net 345 = mbk_sig910 
* net 346 = mbk_sig912 
* net 347 = mbk_sig720 
* net 348 = mbk_sig719 
* net 349 = mbk_sig762 
* net 350 = mbk_sig761 
* net 351 = mbk_sig801 
* net 352 = mbk_sig800 
* net 353 = mbk_sig855 
* net 354 = mbk_sig856 
* net 355 = mbk_sig798 
* net 356 = mbk_sig757 
* net 357 = mbk_sig759 
* net 358 = mbk_sig567 
* net 359 = mbk_sig566 
* net 360 = mbk_sig624 
* net 361 = mbk_sig623 
* net 362 = mbk_sig681 
* net 363 = mbk_sig682 
* net 364 = mbk_sig680 
* net 365 = mbk_sig679 
* net 366 = mbk_sig677 
* net 367 = mbk_sig622 
* net 368 = mbk_sig621 
* net 369 = mbk_sig451 
* net 370 = mbk_sig450 
* net 371 = mbk_sig449 
* net 372 = mbk_sig448 
* net 373 = mbk_sig489 
* net 374 = mbk_sig490 
* net 375 = mbk_sig527 
* net 376 = mbk_sig526 
* net 377 = mbk_sig487 
* net 378 = mbk_sig445 
* net 379 = mbk_sig444 
* net 380 = mbk_sig255 
* net 381 = mbk_sig254 
* net 382 = mbk_sig295 
* net 383 = mbk_sig296 
* net 384 = mbk_sig335 
* net 385 = mbk_sig336 
* net 386 = mbk_sig391 
* net 387 = mbk_sig390 
* net 388 = mbk_sig333 
* net 389 = mbk_sig291 
* net 390 = mbk_sig293 
* net 391 = mbk_sig118 
* net 392 = mbk_sig120 
* net 393 = mbk_sig141 
* net 394 = mbk_sig140 
* net 395 = mbk_sig71 
* net 396 = mbk_sig75 
* net 397 = mbk_sig65 
* net 398 = mbk_sig62 
* net 399 = mbk_sig28 
* net 400 = mbk_sig207 
* net 401 = mbk_sig215 
* net 402 = mbk_sig228 
* net 403 = mbk_sig227 
* net 404 = mbk_sig146 
* net 405 = mbk_sig170 
* net 406 = mbk_sig197 
* net 407 = mbk_sig42 
* net 408 = mbk_sig41 
* net 409 = mbk_sig208 
* net 410 = mbk_sig216 
* net 411 = mbk_sig229 
* net 412 = mbk_sig230 
* net 413 = mbk_sig148 
* net 414 = mbk_sig171 
* net 415 = mbk_sig198 
* net 416 = mbk_sig46 
* net 417 = mbk_sig48 
* net 418 = mbk_sig209 
* net 419 = mbk_sig217 
* net 420 = mbk_sig232 
* net 421 = mbk_sig231 
* net 422 = mbk_sig151 
* net 423 = mbk_sig174 
* net 424 = mbk_sig199 
* net 425 = mbk_sig54 
* net 426 = mbk_sig51 
* net 427 = mbk_sig210 
* net 428 = mbk_sig218 
* net 429 = mbk_sig233 
* net 430 = mbk_sig234 
* net 431 = mbk_sig152 
* net 432 = mbk_sig175 
* net 433 = mbk_sig200 
* net 434 = mbk_sig56 
* net 435 = mbk_sig58 
* net 436 = rbit_0_0.ram_127_1.m0_s 
* net 437 = rbit_0_0.ram_127_1.m1_s 
* net 438 = rbit_0_0.ram_127_0.m0_s 
* net 439 = rbit_0_0.ram_127_0.m1_s 
* net 440 = rbit_0_0.ram_126_1.m0_s 
* net 441 = rbit_0_0.ram_126_1.m1_s 
* net 442 = rbit_0_0.ram_126_0.m0_s 
* net 443 = rbit_0_0.ram_126_0.m1_s 
* net 444 = rbit_0_0.ram_125_1.m0_s 
* net 445 = rbit_0_0.ram_125_1.m1_s 
* net 446 = rbit_0_0.ram_125_0.m0_s 
* net 447 = rbit_0_0.ram_125_0.m1_s 
* net 448 = rbit_0_0.ram_124_1.m0_s 
* net 449 = rbit_0_0.ram_124_1.m1_s 
* net 450 = rbit_0_0.ram_124_0.m0_s 
* net 451 = rbit_0_0.ram_124_0.m1_s 
* net 452 = rbit_0_0.ram_123_1.m0_s 
* net 453 = rbit_0_0.ram_123_1.m1_s 
* net 454 = rbit_0_0.ram_123_0.m0_s 
* net 455 = rbit_0_0.ram_123_0.m1_s 
* net 456 = rbit_0_0.ram_122_1.m0_s 
* net 457 = rbit_0_0.ram_122_1.m1_s 
* net 458 = rbit_0_0.ram_122_0.m0_s 
* net 459 = rbit_0_0.ram_122_0.m1_s 
* net 460 = rbit_0_0.ram_121_1.m0_s 
* net 461 = rbit_0_0.ram_121_1.m1_s 
* net 462 = rbit_0_0.ram_121_0.m0_s 
* net 463 = rbit_0_0.ram_121_0.m1_s 
* net 464 = rbit_0_0.ram_120_1.m0_s 
* net 465 = rbit_0_0.ram_120_1.m1_s 
* net 466 = rbit_0_0.ram_120_0.m0_s 
* net 467 = rbit_0_0.ram_120_0.m1_s 
* net 468 = rbit_0_0.ram_119_1.m0_s 
* net 469 = rbit_0_0.ram_119_1.m1_s 
* net 470 = rbit_0_0.ram_119_0.m0_s 
* net 471 = rbit_0_0.ram_119_0.m1_s 
* net 472 = rbit_0_0.ram_118_1.m0_s 
* net 473 = rbit_0_0.ram_118_1.m1_s 
* net 474 = rbit_0_0.ram_118_0.m0_s 
* net 475 = rbit_0_0.ram_118_0.m1_s 
* net 476 = rbit_0_0.ram_117_1.m0_s 
* net 477 = rbit_0_0.ram_117_1.m1_s 
* net 478 = rbit_0_0.ram_117_0.m0_s 
* net 479 = rbit_0_0.ram_117_0.m1_s 
* net 480 = rbit_0_0.ram_116_1.m0_s 
* net 481 = rbit_0_0.ram_116_1.m1_s 
* net 482 = rbit_0_0.ram_116_0.m0_s 
* net 483 = rbit_0_0.ram_116_0.m1_s 
* net 484 = rbit_0_0.ram_115_1.m0_s 
* net 485 = rbit_0_0.ram_115_1.m1_s 
* net 486 = rbit_0_0.ram_115_0.m0_s 
* net 487 = rbit_0_0.ram_115_0.m1_s 
* net 488 = rbit_0_0.ram_114_1.m0_s 
* net 489 = rbit_0_0.ram_114_1.m1_s 
* net 490 = rbit_0_0.ram_114_0.m0_s 
* net 491 = rbit_0_0.ram_114_0.m1_s 
* net 492 = rbit_0_0.ram_113_1.m0_s 
* net 493 = rbit_0_0.ram_113_1.m1_s 
* net 494 = rbit_0_0.ram_113_0.m0_s 
* net 495 = rbit_0_0.ram_113_0.m1_s 
* net 496 = rbit_0_0.ram_112_1.m0_s 
* net 497 = rbit_0_0.ram_112_1.m1_s 
* net 498 = rbit_0_0.ram_112_0.m0_s 
* net 499 = rbit_0_0.ram_112_0.m1_s 
* net 500 = rbit_0_0.ram_111_1.m0_s 
* net 501 = rbit_0_0.ram_111_1.m1_s 
* net 502 = rbit_0_0.ram_111_0.m0_s 
* net 503 = rbit_0_0.ram_111_0.m1_s 
* net 504 = rbit_0_0.ram_110_1.m0_s 
* net 505 = rbit_0_0.ram_110_1.m1_s 
* net 506 = rbit_0_0.ram_110_0.m0_s 
* net 507 = rbit_0_0.ram_110_0.m1_s 
* net 508 = rbit_0_0.ram_109_1.m0_s 
* net 509 = rbit_0_0.ram_109_1.m1_s 
* net 510 = rbit_0_0.ram_109_0.m0_s 
* net 511 = rbit_0_0.ram_109_0.m1_s 
* net 512 = rbit_0_0.ram_108_1.m0_s 
* net 513 = rbit_0_0.ram_108_1.m1_s 
* net 514 = rbit_0_0.ram_108_0.m0_s 
* net 515 = rbit_0_0.ram_108_0.m1_s 
* net 516 = rbit_0_0.ram_107_1.m0_s 
* net 517 = rbit_0_0.ram_107_1.m1_s 
* net 518 = rbit_0_0.ram_107_0.m0_s 
* net 519 = rbit_0_0.ram_107_0.m1_s 
* net 520 = rbit_0_0.ram_106_1.m0_s 
* net 521 = rbit_0_0.ram_106_1.m1_s 
* net 522 = rbit_0_0.ram_106_0.m0_s 
* net 523 = rbit_0_0.ram_106_0.m1_s 
* net 524 = rbit_0_0.ram_105_1.m0_s 
* net 525 = rbit_0_0.ram_105_1.m1_s 
* net 526 = rbit_0_0.ram_105_0.m0_s 
* net 527 = rbit_0_0.ram_105_0.m1_s 
* net 528 = rbit_0_0.ram_104_1.m0_s 
* net 529 = rbit_0_0.ram_104_1.m1_s 
* net 530 = rbit_0_0.ram_104_0.m0_s 
* net 531 = rbit_0_0.ram_104_0.m1_s 
* net 532 = rbit_0_0.ram_103_1.m0_s 
* net 533 = rbit_0_0.ram_103_1.m1_s 
* net 534 = rbit_0_0.ram_103_0.m0_s 
* net 535 = rbit_0_0.ram_103_0.m1_s 
* net 536 = rbit_0_0.ram_102_1.m0_s 
* net 537 = rbit_0_0.ram_102_1.m1_s 
* net 538 = rbit_0_0.ram_102_0.m0_s 
* net 539 = rbit_0_0.ram_102_0.m1_s 
* net 540 = rbit_0_0.ram_101_1.m0_s 
* net 541 = rbit_0_0.ram_101_1.m1_s 
* net 542 = rbit_0_0.ram_101_0.m0_s 
* net 543 = rbit_0_0.ram_101_0.m1_s 
* net 544 = rbit_0_0.ram_100_1.m0_s 
* net 545 = rbit_0_0.ram_100_1.m1_s 
* net 546 = rbit_0_0.ram_100_0.m0_s 
* net 547 = rbit_0_0.ram_100_0.m1_s 
* net 548 = rbit_0_0.ram_99_1.m0_s 
* net 549 = rbit_0_0.ram_99_1.m1_s 
* net 550 = rbit_0_0.ram_99_0.m0_s 
* net 551 = rbit_0_0.ram_99_0.m1_s 
* net 552 = rbit_0_0.ram_98_1.m0_s 
* net 553 = rbit_0_0.ram_98_1.m1_s 
* net 554 = rbit_0_0.ram_98_0.m0_s 
* net 555 = rbit_0_0.ram_98_0.m1_s 
* net 556 = rbit_0_0.ram_97_1.m0_s 
* net 557 = rbit_0_0.ram_97_1.m1_s 
* net 558 = rbit_0_0.ram_97_0.m0_s 
* net 559 = rbit_0_0.ram_97_0.m1_s 
* net 560 = rbit_0_0.ram_96_1.m0_s 
* net 561 = rbit_0_0.ram_96_1.m1_s 
* net 562 = rbit_0_0.ram_96_0.m0_s 
* net 563 = rbit_0_0.ram_96_0.m1_s 
* net 564 = rbit_0_0.ram_95_1.m0_s 
* net 565 = rbit_0_0.ram_95_1.m1_s 
* net 566 = rbit_0_0.ram_95_0.m0_s 
* net 567 = rbit_0_0.ram_95_0.m1_s 
* net 568 = rbit_0_0.ram_94_1.m0_s 
* net 569 = rbit_0_0.ram_94_1.m1_s 
* net 570 = rbit_0_0.ram_94_0.m0_s 
* net 571 = rbit_0_0.ram_94_0.m1_s 
* net 572 = rbit_0_0.ram_93_1.m0_s 
* net 573 = rbit_0_0.ram_93_1.m1_s 
* net 574 = rbit_0_0.ram_93_0.m0_s 
* net 575 = rbit_0_0.ram_93_0.m1_s 
* net 576 = rbit_0_0.ram_92_1.m0_s 
* net 577 = rbit_0_0.ram_92_1.m1_s 
* net 578 = rbit_0_0.ram_92_0.m0_s 
* net 579 = rbit_0_0.ram_92_0.m1_s 
* net 580 = rbit_0_0.ram_91_1.m0_s 
* net 581 = rbit_0_0.ram_91_1.m1_s 
* net 582 = rbit_0_0.ram_91_0.m0_s 
* net 583 = rbit_0_0.ram_91_0.m1_s 
* net 584 = rbit_0_0.ram_90_1.m0_s 
* net 585 = rbit_0_0.ram_90_1.m1_s 
* net 586 = rbit_0_0.ram_90_0.m0_s 
* net 587 = rbit_0_0.ram_90_0.m1_s 
* net 588 = rbit_0_0.ram_89_1.m0_s 
* net 589 = rbit_0_0.ram_89_1.m1_s 
* net 590 = rbit_0_0.ram_89_0.m0_s 
* net 591 = rbit_0_0.ram_89_0.m1_s 
* net 592 = rbit_0_0.ram_88_1.m0_s 
* net 593 = rbit_0_0.ram_88_1.m1_s 
* net 594 = rbit_0_0.ram_88_0.m0_s 
* net 595 = rbit_0_0.ram_88_0.m1_s 
* net 596 = rbit_0_0.ram_87_1.m0_s 
* net 597 = rbit_0_0.ram_87_1.m1_s 
* net 598 = rbit_0_0.ram_87_0.m0_s 
* net 599 = rbit_0_0.ram_87_0.m1_s 
* net 600 = rbit_0_0.ram_86_1.m0_s 
* net 601 = rbit_0_0.ram_86_1.m1_s 
* net 602 = rbit_0_0.ram_86_0.m0_s 
* net 603 = rbit_0_0.ram_86_0.m1_s 
* net 604 = rbit_0_0.ram_85_1.m0_s 
* net 605 = rbit_0_0.ram_85_1.m1_s 
* net 606 = rbit_0_0.ram_85_0.m0_s 
* net 607 = rbit_0_0.ram_85_0.m1_s 
* net 608 = rbit_0_0.ram_84_1.m0_s 
* net 609 = rbit_0_0.ram_84_1.m1_s 
* net 610 = rbit_0_0.ram_84_0.m0_s 
* net 611 = rbit_0_0.ram_84_0.m1_s 
* net 612 = rbit_0_0.ram_83_1.m0_s 
* net 613 = rbit_0_0.ram_83_1.m1_s 
* net 614 = rbit_0_0.ram_83_0.m0_s 
* net 615 = rbit_0_0.ram_83_0.m1_s 
* net 616 = rbit_0_0.ram_82_1.m0_s 
* net 617 = rbit_0_0.ram_82_1.m1_s 
* net 618 = rbit_0_0.ram_82_0.m0_s 
* net 619 = rbit_0_0.ram_82_0.m1_s 
* net 620 = rbit_0_0.ram_81_1.m0_s 
* net 621 = rbit_0_0.ram_81_1.m1_s 
* net 622 = rbit_0_0.ram_81_0.m0_s 
* net 623 = rbit_0_0.ram_81_0.m1_s 
* net 624 = rbit_0_0.ram_80_1.m0_s 
* net 625 = rbit_0_0.ram_80_1.m1_s 
* net 626 = rbit_0_0.ram_80_0.m0_s 
* net 627 = rbit_0_0.ram_80_0.m1_s 
* net 628 = rbit_0_0.ram_79_1.m0_s 
* net 629 = rbit_0_0.ram_79_1.m1_s 
* net 630 = rbit_0_0.ram_79_0.m0_s 
* net 631 = rbit_0_0.ram_79_0.m1_s 
* net 632 = rbit_0_0.ram_78_1.m0_s 
* net 633 = rbit_0_0.ram_78_1.m1_s 
* net 634 = rbit_0_0.ram_78_0.m0_s 
* net 635 = rbit_0_0.ram_78_0.m1_s 
* net 636 = rbit_0_0.ram_77_1.m0_s 
* net 637 = rbit_0_0.ram_77_1.m1_s 
* net 638 = rbit_0_0.ram_77_0.m0_s 
* net 639 = rbit_0_0.ram_77_0.m1_s 
* net 640 = rbit_0_0.ram_76_1.m0_s 
* net 641 = rbit_0_0.ram_76_1.m1_s 
* net 642 = rbit_0_0.ram_76_0.m0_s 
* net 643 = rbit_0_0.ram_76_0.m1_s 
* net 644 = rbit_0_0.ram_75_1.m0_s 
* net 645 = rbit_0_0.ram_75_1.m1_s 
* net 646 = rbit_0_0.ram_75_0.m0_s 
* net 647 = rbit_0_0.ram_75_0.m1_s 
* net 648 = rbit_0_0.ram_74_1.m0_s 
* net 649 = rbit_0_0.ram_74_1.m1_s 
* net 650 = rbit_0_0.ram_74_0.m0_s 
* net 651 = rbit_0_0.ram_74_0.m1_s 
* net 652 = rbit_0_0.ram_73_1.m0_s 
* net 653 = rbit_0_0.ram_73_1.m1_s 
* net 654 = rbit_0_0.ram_73_0.m0_s 
* net 655 = rbit_0_0.ram_73_0.m1_s 
* net 656 = rbit_0_0.ram_72_1.m0_s 
* net 657 = rbit_0_0.ram_72_1.m1_s 
* net 658 = rbit_0_0.ram_72_0.m0_s 
* net 659 = rbit_0_0.ram_72_0.m1_s 
* net 660 = rbit_0_0.ram_71_1.m0_s 
* net 661 = rbit_0_0.ram_71_1.m1_s 
* net 662 = rbit_0_0.ram_71_0.m0_s 
* net 663 = rbit_0_0.ram_71_0.m1_s 
* net 664 = rbit_0_0.ram_70_1.m0_s 
* net 665 = rbit_0_0.ram_70_1.m1_s 
* net 666 = rbit_0_0.ram_70_0.m0_s 
* net 667 = rbit_0_0.ram_70_0.m1_s 
* net 668 = rbit_0_0.ram_69_1.m0_s 
* net 669 = rbit_0_0.ram_69_1.m1_s 
* net 670 = rbit_0_0.ram_69_0.m0_s 
* net 671 = rbit_0_0.ram_69_0.m1_s 
* net 672 = rbit_0_0.ram_68_1.m0_s 
* net 673 = rbit_0_0.ram_68_1.m1_s 
* net 674 = rbit_0_0.ram_68_0.m0_s 
* net 675 = rbit_0_0.ram_68_0.m1_s 
* net 676 = rbit_0_0.ram_67_1.m0_s 
* net 677 = rbit_0_0.ram_67_1.m1_s 
* net 678 = rbit_0_0.ram_67_0.m0_s 
* net 679 = rbit_0_0.ram_67_0.m1_s 
* net 680 = rbit_0_0.ram_66_1.m0_s 
* net 681 = rbit_0_0.ram_66_1.m1_s 
* net 682 = rbit_0_0.ram_66_0.m0_s 
* net 683 = rbit_0_0.ram_66_0.m1_s 
* net 684 = rbit_0_0.ram_65_1.m0_s 
* net 685 = rbit_0_0.ram_65_1.m1_s 
* net 686 = rbit_0_0.ram_65_0.m0_s 
* net 687 = rbit_0_0.ram_65_0.m1_s 
* net 688 = rbit_0_0.ram_64_1.m0_s 
* net 689 = rbit_0_0.ram_64_1.m1_s 
* net 690 = rbit_0_0.ram_64_0.m0_s 
* net 691 = rbit_0_0.ram_64_0.m1_s 
* net 692 = rbit_0_0.ram_63_1.m0_s 
* net 693 = rbit_0_0.ram_63_1.m1_s 
* net 694 = rbit_0_0.ram_63_0.m0_s 
* net 695 = rbit_0_0.ram_63_0.m1_s 
* net 696 = rbit_0_0.ram_62_1.m0_s 
* net 697 = rbit_0_0.ram_62_1.m1_s 
* net 698 = rbit_0_0.ram_62_0.m0_s 
* net 699 = rbit_0_0.ram_62_0.m1_s 
* net 700 = rbit_0_0.ram_61_1.m0_s 
* net 701 = rbit_0_0.ram_61_1.m1_s 
* net 702 = rbit_0_0.ram_61_0.m0_s 
* net 703 = rbit_0_0.ram_61_0.m1_s 
* net 704 = rbit_0_0.ram_60_1.m0_s 
* net 705 = rbit_0_0.ram_60_1.m1_s 
* net 706 = rbit_0_0.ram_60_0.m0_s 
* net 707 = rbit_0_0.ram_60_0.m1_s 
* net 708 = rbit_0_0.ram_59_1.m0_s 
* net 709 = rbit_0_0.ram_59_1.m1_s 
* net 710 = rbit_0_0.ram_59_0.m0_s 
* net 711 = rbit_0_0.ram_59_0.m1_s 
* net 712 = rbit_0_0.ram_58_1.m0_s 
* net 713 = rbit_0_0.ram_58_1.m1_s 
* net 714 = rbit_0_0.ram_58_0.m0_s 
* net 715 = rbit_0_0.ram_58_0.m1_s 
* net 716 = rbit_0_0.ram_57_1.m0_s 
* net 717 = rbit_0_0.ram_57_1.m1_s 
* net 718 = rbit_0_0.ram_57_0.m0_s 
* net 719 = rbit_0_0.ram_57_0.m1_s 
* net 720 = rbit_0_0.ram_56_1.m0_s 
* net 721 = rbit_0_0.ram_56_1.m1_s 
* net 722 = rbit_0_0.ram_56_0.m0_s 
* net 723 = rbit_0_0.ram_56_0.m1_s 
* net 724 = rbit_0_0.ram_55_1.m0_s 
* net 725 = rbit_0_0.ram_55_1.m1_s 
* net 726 = rbit_0_0.ram_55_0.m0_s 
* net 727 = rbit_0_0.ram_55_0.m1_s 
* net 728 = rbit_0_0.ram_54_1.m0_s 
* net 729 = rbit_0_0.ram_54_1.m1_s 
* net 730 = rbit_0_0.ram_54_0.m0_s 
* net 731 = rbit_0_0.ram_54_0.m1_s 
* net 732 = rbit_0_0.ram_53_1.m0_s 
* net 733 = rbit_0_0.ram_53_1.m1_s 
* net 734 = rbit_0_0.ram_53_0.m0_s 
* net 735 = rbit_0_0.ram_53_0.m1_s 
* net 736 = rbit_0_0.ram_52_1.m0_s 
* net 737 = rbit_0_0.ram_52_1.m1_s 
* net 738 = rbit_0_0.ram_52_0.m0_s 
* net 739 = rbit_0_0.ram_52_0.m1_s 
* net 740 = rbit_0_0.ram_51_1.m0_s 
* net 741 = rbit_0_0.ram_51_1.m1_s 
* net 742 = rbit_0_0.ram_51_0.m0_s 
* net 743 = rbit_0_0.ram_51_0.m1_s 
* net 744 = rbit_0_0.ram_50_1.m0_s 
* net 745 = rbit_0_0.ram_50_1.m1_s 
* net 746 = rbit_0_0.ram_50_0.m0_s 
* net 747 = rbit_0_0.ram_50_0.m1_s 
* net 748 = rbit_0_0.ram_49_1.m0_s 
* net 749 = rbit_0_0.ram_49_1.m1_s 
* net 750 = rbit_0_0.ram_49_0.m0_s 
* net 751 = rbit_0_0.ram_49_0.m1_s 
* net 752 = rbit_0_0.ram_48_1.m0_s 
* net 753 = rbit_0_0.ram_48_1.m1_s 
* net 754 = rbit_0_0.ram_48_0.m0_s 
* net 755 = rbit_0_0.ram_48_0.m1_s 
* net 756 = rbit_0_0.ram_47_1.m0_s 
* net 757 = rbit_0_0.ram_47_1.m1_s 
* net 758 = rbit_0_0.ram_47_0.m0_s 
* net 759 = rbit_0_0.ram_47_0.m1_s 
* net 760 = rbit_0_0.ram_46_1.m0_s 
* net 761 = rbit_0_0.ram_46_1.m1_s 
* net 762 = rbit_0_0.ram_46_0.m0_s 
* net 763 = rbit_0_0.ram_46_0.m1_s 
* net 764 = rbit_0_0.ram_45_1.m0_s 
* net 765 = rbit_0_0.ram_45_1.m1_s 
* net 766 = rbit_0_0.ram_45_0.m0_s 
* net 767 = rbit_0_0.ram_45_0.m1_s 
* net 768 = rbit_0_0.ram_44_1.m0_s 
* net 769 = rbit_0_0.ram_44_1.m1_s 
* net 770 = rbit_0_0.ram_44_0.m0_s 
* net 771 = rbit_0_0.ram_44_0.m1_s 
* net 772 = rbit_0_0.ram_43_1.m0_s 
* net 773 = rbit_0_0.ram_43_1.m1_s 
* net 774 = rbit_0_0.ram_43_0.m0_s 
* net 775 = rbit_0_0.ram_43_0.m1_s 
* net 776 = rbit_0_0.ram_42_1.m0_s 
* net 777 = rbit_0_0.ram_42_1.m1_s 
* net 778 = rbit_0_0.ram_42_0.m0_s 
* net 779 = rbit_0_0.ram_42_0.m1_s 
* net 780 = rbit_0_0.ram_41_1.m0_s 
* net 781 = rbit_0_0.ram_41_1.m1_s 
* net 782 = rbit_0_0.ram_41_0.m0_s 
* net 783 = rbit_0_0.ram_41_0.m1_s 
* net 784 = rbit_0_0.ram_40_1.m0_s 
* net 785 = rbit_0_0.ram_40_1.m1_s 
* net 786 = rbit_0_0.ram_40_0.m0_s 
* net 787 = rbit_0_0.ram_40_0.m1_s 
* net 788 = rbit_0_0.ram_39_1.m0_s 
* net 789 = rbit_0_0.ram_39_1.m1_s 
* net 790 = rbit_0_0.ram_39_0.m0_s 
* net 791 = rbit_0_0.ram_39_0.m1_s 
* net 792 = rbit_0_0.ram_38_1.m0_s 
* net 793 = rbit_0_0.ram_38_1.m1_s 
* net 794 = rbit_0_0.ram_38_0.m0_s 
* net 795 = rbit_0_0.ram_38_0.m1_s 
* net 796 = rbit_0_0.ram_37_1.m0_s 
* net 797 = rbit_0_0.ram_37_1.m1_s 
* net 798 = rbit_0_0.ram_37_0.m0_s 
* net 799 = rbit_0_0.ram_37_0.m1_s 
* net 800 = rbit_0_0.ram_36_1.m0_s 
* net 801 = rbit_0_0.ram_36_1.m1_s 
* net 802 = rbit_0_0.ram_36_0.m0_s 
* net 803 = rbit_0_0.ram_36_0.m1_s 
* net 804 = rbit_0_0.ram_35_1.m0_s 
* net 805 = rbit_0_0.ram_35_1.m1_s 
* net 806 = rbit_0_0.ram_35_0.m0_s 
* net 807 = rbit_0_0.ram_35_0.m1_s 
* net 808 = rbit_0_0.ram_34_1.m0_s 
* net 809 = rbit_0_0.ram_34_1.m1_s 
* net 810 = rbit_0_0.ram_34_0.m0_s 
* net 811 = rbit_0_0.ram_34_0.m1_s 
* net 812 = rbit_0_0.ram_33_1.m0_s 
* net 813 = rbit_0_0.ram_33_1.m1_s 
* net 814 = rbit_0_0.ram_33_0.m0_s 
* net 815 = rbit_0_0.ram_33_0.m1_s 
* net 816 = rbit_0_0.ram_32_1.m0_s 
* net 817 = rbit_0_0.ram_32_1.m1_s 
* net 818 = rbit_0_0.ram_32_0.m0_s 
* net 819 = rbit_0_0.ram_32_0.m1_s 
* net 820 = rbit_0_0.ram_31_1.m0_s 
* net 821 = rbit_0_0.ram_31_1.m1_s 
* net 822 = rbit_0_0.ram_31_0.m0_s 
* net 823 = rbit_0_0.ram_31_0.m1_s 
* net 824 = rbit_0_0.ram_30_1.m0_s 
* net 825 = rbit_0_0.ram_30_1.m1_s 
* net 826 = rbit_0_0.ram_30_0.m0_s 
* net 827 = rbit_0_0.ram_30_0.m1_s 
* net 828 = rbit_0_0.ram_29_1.m0_s 
* net 829 = rbit_0_0.ram_29_1.m1_s 
* net 830 = rbit_0_0.ram_29_0.m0_s 
* net 831 = rbit_0_0.ram_29_0.m1_s 
* net 832 = rbit_0_0.ram_28_1.m0_s 
* net 833 = rbit_0_0.ram_28_1.m1_s 
* net 834 = rbit_0_0.ram_28_0.m0_s 
* net 835 = rbit_0_0.ram_28_0.m1_s 
* net 836 = rbit_0_0.ram_27_1.m0_s 
* net 837 = rbit_0_0.ram_27_1.m1_s 
* net 838 = rbit_0_0.ram_27_0.m0_s 
* net 839 = rbit_0_0.ram_27_0.m1_s 
* net 840 = rbit_0_0.ram_26_1.m0_s 
* net 841 = rbit_0_0.ram_26_1.m1_s 
* net 842 = rbit_0_0.ram_26_0.m0_s 
* net 843 = rbit_0_0.ram_26_0.m1_s 
* net 844 = rbit_0_0.ram_25_1.m0_s 
* net 845 = rbit_0_0.ram_25_1.m1_s 
* net 846 = rbit_0_0.ram_25_0.m0_s 
* net 847 = rbit_0_0.ram_25_0.m1_s 
* net 848 = rbit_0_0.ram_24_1.m0_s 
* net 849 = rbit_0_0.ram_24_1.m1_s 
* net 850 = rbit_0_0.ram_24_0.m0_s 
* net 851 = rbit_0_0.ram_24_0.m1_s 
* net 852 = rbit_0_0.ram_23_1.m0_s 
* net 853 = rbit_0_0.ram_23_1.m1_s 
* net 854 = rbit_0_0.ram_23_0.m0_s 
* net 855 = rbit_0_0.ram_23_0.m1_s 
* net 856 = rbit_0_0.ram_22_1.m0_s 
* net 857 = rbit_0_0.ram_22_1.m1_s 
* net 858 = rbit_0_0.ram_22_0.m0_s 
* net 859 = rbit_0_0.ram_22_0.m1_s 
* net 860 = rbit_0_0.ram_21_1.m0_s 
* net 861 = rbit_0_0.ram_21_1.m1_s 
* net 862 = rbit_0_0.ram_21_0.m0_s 
* net 863 = rbit_0_0.ram_21_0.m1_s 
* net 864 = rbit_0_0.ram_20_1.m0_s 
* net 865 = rbit_0_0.ram_20_1.m1_s 
* net 866 = rbit_0_0.ram_20_0.m0_s 
* net 867 = rbit_0_0.ram_20_0.m1_s 
* net 868 = rbit_0_0.ram_19_1.m0_s 
* net 869 = rbit_0_0.ram_19_1.m1_s 
* net 870 = rbit_0_0.ram_19_0.m0_s 
* net 871 = rbit_0_0.ram_19_0.m1_s 
* net 872 = rbit_0_0.ram_18_1.m0_s 
* net 873 = rbit_0_0.ram_18_1.m1_s 
* net 874 = rbit_0_0.ram_18_0.m0_s 
* net 875 = rbit_0_0.ram_18_0.m1_s 
* net 876 = rbit_0_0.ram_17_1.m0_s 
* net 877 = rbit_0_0.ram_17_1.m1_s 
* net 878 = rbit_0_0.ram_17_0.m0_s 
* net 879 = rbit_0_0.ram_17_0.m1_s 
* net 880 = rbit_0_0.ram_16_1.m0_s 
* net 881 = rbit_0_0.ram_16_1.m1_s 
* net 882 = rbit_0_0.ram_16_0.m0_s 
* net 883 = rbit_0_0.ram_16_0.m1_s 
* net 884 = rbit_0_0.ram_15_1.m0_s 
* net 885 = rbit_0_0.ram_15_1.m1_s 
* net 886 = rbit_0_0.ram_15_0.m0_s 
* net 887 = rbit_0_0.ram_15_0.m1_s 
* net 888 = rbit_0_0.ram_14_1.m0_s 
* net 889 = rbit_0_0.ram_14_1.m1_s 
* net 890 = rbit_0_0.ram_14_0.m0_s 
* net 891 = rbit_0_0.ram_14_0.m1_s 
* net 892 = rbit_0_0.ram_13_1.m0_s 
* net 893 = rbit_0_0.ram_13_1.m1_s 
* net 894 = rbit_0_0.ram_13_0.m0_s 
* net 895 = rbit_0_0.ram_13_0.m1_s 
* net 896 = rbit_0_0.ram_12_1.m0_s 
* net 897 = rbit_0_0.ram_12_1.m1_s 
* net 898 = rbit_0_0.ram_12_0.m0_s 
* net 899 = rbit_0_0.ram_12_0.m1_s 
* net 900 = rbit_0_0.ram_11_1.m0_s 
* net 901 = rbit_0_0.ram_11_1.m1_s 
* net 902 = rbit_0_0.ram_11_0.m0_s 
* net 903 = rbit_0_0.ram_11_0.m1_s 
* net 904 = rbit_0_0.ram_10_1.m0_s 
* net 905 = rbit_0_0.ram_10_1.m1_s 
* net 906 = rbit_0_0.ram_10_0.m0_s 
* net 907 = rbit_0_0.ram_10_0.m1_s 
* net 908 = rbit_0_0.ram_9_1.m0_s 
* net 909 = rbit_0_0.ram_9_1.m1_s 
* net 910 = rbit_0_0.ram_9_0.m0_s 
* net 911 = rbit_0_0.ram_9_0.m1_s 
* net 912 = rbit_0_0.ram_8_1.m0_s 
* net 913 = rbit_0_0.ram_8_1.m1_s 
* net 914 = rbit_0_0.ram_8_0.m0_s 
* net 915 = rbit_0_0.ram_8_0.m1_s 
* net 916 = rbit_0_0.ram_7_1.m0_s 
* net 917 = rbit_0_0.ram_7_1.m1_s 
* net 918 = rbit_0_0.ram_7_0.m0_s 
* net 919 = rbit_0_0.ram_7_0.m1_s 
* net 920 = rbit_0_0.ram_6_1.m0_s 
* net 921 = rbit_0_0.ram_6_1.m1_s 
* net 922 = rbit_0_0.ram_6_0.m0_s 
* net 923 = rbit_0_0.ram_6_0.m1_s 
* net 924 = rbit_0_0.ram_5_1.m0_s 
* net 925 = rbit_0_0.ram_5_1.m1_s 
* net 926 = rbit_0_0.ram_5_0.m0_s 
* net 927 = rbit_0_0.ram_5_0.m1_s 
* net 928 = rbit_0_0.ram_4_1.m0_s 
* net 929 = rbit_0_0.ram_4_1.m1_s 
* net 930 = rbit_0_0.ram_4_0.m0_s 
* net 931 = rbit_0_0.ram_4_0.m1_s 
* net 932 = rbit_0_0.ram_3_1.m0_s 
* net 933 = rbit_0_0.ram_3_1.m1_s 
* net 934 = rbit_0_0.ram_3_0.m0_s 
* net 935 = rbit_0_0.ram_3_0.m1_s 
* net 936 = rbit_0_0.ram_2_1.m0_s 
* net 937 = rbit_0_0.ram_2_1.m1_s 
* net 938 = rbit_0_0.ram_2_0.m0_s 
* net 939 = rbit_0_0.ram_2_0.m1_s 
* net 940 = rbit_0_0.ram_1_1.m0_s 
* net 941 = rbit_0_0.ram_1_1.m1_s 
* net 942 = rbit_0_0.ram_1_0.m0_s 
* net 943 = rbit_0_0.ram_1_0.m1_s 
* net 944 = rbit_0_0.ram_0_1.m0_s 
* net 945 = rbit_0_0.ram_0_1.m1_s 
* net 946 = rbit_0_0.ram_0_0.m0_s 
* net 947 = rbit_0_0.ram_0_0.m1_s 
* net 948 = mbk_sig133 
* net 949 = mbk_sig109 
* net 950 = mbk_sig158 
* net 951 = mbk_sig108 
* net 952 = mbk_sig180 
* net 953 = mbk_sig4 
* net 954 = mbk_sig2 
* net 955 = mbk_sig66 
* net 956 = mbk_sig98 
* net 957 = mbk_sig90 
* net 958 = mbk_sig82 
* net 959 = rbit_1_0.ram_127_1.m0_s 
* net 960 = rbit_1_0.ram_127_1.m1_s 
* net 961 = rbit_1_0.ram_127_0.m0_s 
* net 962 = rbit_1_0.ram_127_0.m1_s 
* net 963 = rbit_1_0.ram_126_1.m0_s 
* net 964 = rbit_1_0.ram_126_1.m1_s 
* net 965 = rbit_1_0.ram_126_0.m0_s 
* net 966 = rbit_1_0.ram_126_0.m1_s 
* net 967 = rbit_1_0.ram_125_1.m0_s 
* net 968 = rbit_1_0.ram_125_1.m1_s 
* net 969 = rbit_1_0.ram_125_0.m0_s 
* net 970 = rbit_1_0.ram_125_0.m1_s 
* net 971 = rbit_1_0.ram_124_1.m0_s 
* net 972 = rbit_1_0.ram_124_1.m1_s 
* net 973 = rbit_1_0.ram_124_0.m0_s 
* net 974 = rbit_1_0.ram_124_0.m1_s 
* net 975 = rbit_1_0.ram_123_1.m0_s 
* net 976 = rbit_1_0.ram_123_1.m1_s 
* net 977 = rbit_1_0.ram_123_0.m0_s 
* net 978 = rbit_1_0.ram_123_0.m1_s 
* net 979 = rbit_1_0.ram_122_1.m0_s 
* net 980 = rbit_1_0.ram_122_1.m1_s 
* net 981 = rbit_1_0.ram_122_0.m0_s 
* net 982 = rbit_1_0.ram_122_0.m1_s 
* net 983 = rbit_1_0.ram_121_1.m0_s 
* net 984 = rbit_1_0.ram_121_1.m1_s 
* net 985 = rbit_1_0.ram_121_0.m0_s 
* net 986 = rbit_1_0.ram_121_0.m1_s 
* net 987 = rbit_1_0.ram_120_1.m0_s 
* net 988 = rbit_1_0.ram_120_1.m1_s 
* net 989 = rbit_1_0.ram_120_0.m0_s 
* net 990 = rbit_1_0.ram_120_0.m1_s 
* net 991 = rbit_1_0.ram_119_1.m0_s 
* net 992 = rbit_1_0.ram_119_1.m1_s 
* net 993 = rbit_1_0.ram_119_0.m0_s 
* net 994 = rbit_1_0.ram_119_0.m1_s 
* net 995 = rbit_1_0.ram_118_1.m0_s 
* net 996 = rbit_1_0.ram_118_1.m1_s 
* net 997 = rbit_1_0.ram_118_0.m0_s 
* net 998 = rbit_1_0.ram_118_0.m1_s 
* net 999 = rbit_1_0.ram_117_1.m0_s 
* net 1000 = rbit_1_0.ram_117_1.m1_s 
* net 1001 = rbit_1_0.ram_117_0.m0_s 
* net 1002 = rbit_1_0.ram_117_0.m1_s 
* net 1003 = rbit_1_0.ram_116_1.m0_s 
* net 1004 = rbit_1_0.ram_116_1.m1_s 
* net 1005 = rbit_1_0.ram_116_0.m0_s 
* net 1006 = rbit_1_0.ram_116_0.m1_s 
* net 1007 = rbit_1_0.ram_115_1.m0_s 
* net 1008 = rbit_1_0.ram_115_1.m1_s 
* net 1009 = rbit_1_0.ram_115_0.m0_s 
* net 1010 = rbit_1_0.ram_115_0.m1_s 
* net 1011 = rbit_1_0.ram_114_1.m0_s 
* net 1012 = rbit_1_0.ram_114_1.m1_s 
* net 1013 = rbit_1_0.ram_114_0.m0_s 
* net 1014 = rbit_1_0.ram_114_0.m1_s 
* net 1015 = rbit_1_0.ram_113_1.m0_s 
* net 1016 = rbit_1_0.ram_113_1.m1_s 
* net 1017 = rbit_1_0.ram_113_0.m0_s 
* net 1018 = rbit_1_0.ram_113_0.m1_s 
* net 1019 = rbit_1_0.ram_112_1.m0_s 
* net 1020 = rbit_1_0.ram_112_1.m1_s 
* net 1021 = rbit_1_0.ram_112_0.m0_s 
* net 1022 = rbit_1_0.ram_112_0.m1_s 
* net 1023 = rbit_1_0.ram_111_1.m0_s 
* net 1024 = rbit_1_0.ram_111_1.m1_s 
* net 1025 = rbit_1_0.ram_111_0.m0_s 
* net 1026 = rbit_1_0.ram_111_0.m1_s 
* net 1027 = rbit_1_0.ram_110_1.m0_s 
* net 1028 = rbit_1_0.ram_110_1.m1_s 
* net 1029 = rbit_1_0.ram_110_0.m0_s 
* net 1030 = rbit_1_0.ram_110_0.m1_s 
* net 1031 = rbit_1_0.ram_109_1.m0_s 
* net 1032 = rbit_1_0.ram_109_1.m1_s 
* net 1033 = rbit_1_0.ram_109_0.m0_s 
* net 1034 = rbit_1_0.ram_109_0.m1_s 
* net 1035 = rbit_1_0.ram_108_1.m0_s 
* net 1036 = rbit_1_0.ram_108_1.m1_s 
* net 1037 = rbit_1_0.ram_108_0.m0_s 
* net 1038 = rbit_1_0.ram_108_0.m1_s 
* net 1039 = rbit_1_0.ram_107_1.m0_s 
* net 1040 = rbit_1_0.ram_107_1.m1_s 
* net 1041 = rbit_1_0.ram_107_0.m0_s 
* net 1042 = rbit_1_0.ram_107_0.m1_s 
* net 1043 = rbit_1_0.ram_106_1.m0_s 
* net 1044 = rbit_1_0.ram_106_1.m1_s 
* net 1045 = rbit_1_0.ram_106_0.m0_s 
* net 1046 = rbit_1_0.ram_106_0.m1_s 
* net 1047 = rbit_1_0.ram_105_1.m0_s 
* net 1048 = rbit_1_0.ram_105_1.m1_s 
* net 1049 = rbit_1_0.ram_105_0.m0_s 
* net 1050 = rbit_1_0.ram_105_0.m1_s 
* net 1051 = rbit_1_0.ram_104_1.m0_s 
* net 1052 = rbit_1_0.ram_104_1.m1_s 
* net 1053 = rbit_1_0.ram_104_0.m0_s 
* net 1054 = rbit_1_0.ram_104_0.m1_s 
* net 1055 = rbit_1_0.ram_103_1.m0_s 
* net 1056 = rbit_1_0.ram_103_1.m1_s 
* net 1057 = rbit_1_0.ram_103_0.m0_s 
* net 1058 = rbit_1_0.ram_103_0.m1_s 
* net 1059 = rbit_1_0.ram_102_1.m0_s 
* net 1060 = rbit_1_0.ram_102_1.m1_s 
* net 1061 = rbit_1_0.ram_102_0.m0_s 
* net 1062 = rbit_1_0.ram_102_0.m1_s 
* net 1063 = rbit_1_0.ram_101_1.m0_s 
* net 1064 = rbit_1_0.ram_101_1.m1_s 
* net 1065 = rbit_1_0.ram_101_0.m0_s 
* net 1066 = rbit_1_0.ram_101_0.m1_s 
* net 1067 = rbit_1_0.ram_100_1.m0_s 
* net 1068 = rbit_1_0.ram_100_1.m1_s 
* net 1069 = rbit_1_0.ram_100_0.m0_s 
* net 1070 = rbit_1_0.ram_100_0.m1_s 
* net 1071 = rbit_1_0.ram_99_1.m0_s 
* net 1072 = rbit_1_0.ram_99_1.m1_s 
* net 1073 = rbit_1_0.ram_99_0.m0_s 
* net 1074 = rbit_1_0.ram_99_0.m1_s 
* net 1075 = rbit_1_0.ram_98_1.m0_s 
* net 1076 = rbit_1_0.ram_98_1.m1_s 
* net 1077 = rbit_1_0.ram_98_0.m0_s 
* net 1078 = rbit_1_0.ram_98_0.m1_s 
* net 1079 = rbit_1_0.ram_97_1.m0_s 
* net 1080 = rbit_1_0.ram_97_1.m1_s 
* net 1081 = rbit_1_0.ram_97_0.m0_s 
* net 1082 = rbit_1_0.ram_97_0.m1_s 
* net 1083 = rbit_1_0.ram_96_1.m0_s 
* net 1084 = rbit_1_0.ram_96_1.m1_s 
* net 1085 = rbit_1_0.ram_96_0.m0_s 
* net 1086 = rbit_1_0.ram_96_0.m1_s 
* net 1087 = rbit_1_0.ram_95_1.m0_s 
* net 1088 = rbit_1_0.ram_95_1.m1_s 
* net 1089 = rbit_1_0.ram_95_0.m0_s 
* net 1090 = rbit_1_0.ram_95_0.m1_s 
* net 1091 = rbit_1_0.ram_94_1.m0_s 
* net 1092 = rbit_1_0.ram_94_1.m1_s 
* net 1093 = rbit_1_0.ram_94_0.m0_s 
* net 1094 = rbit_1_0.ram_94_0.m1_s 
* net 1095 = rbit_1_0.ram_93_1.m0_s 
* net 1096 = rbit_1_0.ram_93_1.m1_s 
* net 1097 = rbit_1_0.ram_93_0.m0_s 
* net 1098 = rbit_1_0.ram_93_0.m1_s 
* net 1099 = rbit_1_0.ram_92_1.m0_s 
* net 1100 = rbit_1_0.ram_92_1.m1_s 
* net 1101 = rbit_1_0.ram_92_0.m0_s 
* net 1102 = rbit_1_0.ram_92_0.m1_s 
* net 1103 = rbit_1_0.ram_91_1.m0_s 
* net 1104 = rbit_1_0.ram_91_1.m1_s 
* net 1105 = rbit_1_0.ram_91_0.m0_s 
* net 1106 = rbit_1_0.ram_91_0.m1_s 
* net 1107 = rbit_1_0.ram_90_1.m0_s 
* net 1108 = rbit_1_0.ram_90_1.m1_s 
* net 1109 = rbit_1_0.ram_90_0.m0_s 
* net 1110 = rbit_1_0.ram_90_0.m1_s 
* net 1111 = rbit_1_0.ram_89_1.m0_s 
* net 1112 = rbit_1_0.ram_89_1.m1_s 
* net 1113 = rbit_1_0.ram_89_0.m0_s 
* net 1114 = rbit_1_0.ram_89_0.m1_s 
* net 1115 = rbit_1_0.ram_88_1.m0_s 
* net 1116 = rbit_1_0.ram_88_1.m1_s 
* net 1117 = rbit_1_0.ram_88_0.m0_s 
* net 1118 = rbit_1_0.ram_88_0.m1_s 
* net 1119 = rbit_1_0.ram_87_1.m0_s 
* net 1120 = rbit_1_0.ram_87_1.m1_s 
* net 1121 = rbit_1_0.ram_87_0.m0_s 
* net 1122 = rbit_1_0.ram_87_0.m1_s 
* net 1123 = rbit_1_0.ram_86_1.m0_s 
* net 1124 = rbit_1_0.ram_86_1.m1_s 
* net 1125 = rbit_1_0.ram_86_0.m0_s 
* net 1126 = rbit_1_0.ram_86_0.m1_s 
* net 1127 = rbit_1_0.ram_85_1.m0_s 
* net 1128 = rbit_1_0.ram_85_1.m1_s 
* net 1129 = rbit_1_0.ram_85_0.m0_s 
* net 1130 = rbit_1_0.ram_85_0.m1_s 
* net 1131 = rbit_1_0.ram_84_1.m0_s 
* net 1132 = rbit_1_0.ram_84_1.m1_s 
* net 1133 = rbit_1_0.ram_84_0.m0_s 
* net 1134 = rbit_1_0.ram_84_0.m1_s 
* net 1135 = rbit_1_0.ram_83_1.m0_s 
* net 1136 = rbit_1_0.ram_83_1.m1_s 
* net 1137 = rbit_1_0.ram_83_0.m0_s 
* net 1138 = rbit_1_0.ram_83_0.m1_s 
* net 1139 = rbit_1_0.ram_82_1.m0_s 
* net 1140 = rbit_1_0.ram_82_1.m1_s 
* net 1141 = rbit_1_0.ram_82_0.m0_s 
* net 1142 = rbit_1_0.ram_82_0.m1_s 
* net 1143 = rbit_1_0.ram_81_1.m0_s 
* net 1144 = rbit_1_0.ram_81_1.m1_s 
* net 1145 = rbit_1_0.ram_81_0.m0_s 
* net 1146 = rbit_1_0.ram_81_0.m1_s 
* net 1147 = rbit_1_0.ram_80_1.m0_s 
* net 1148 = rbit_1_0.ram_80_1.m1_s 
* net 1149 = rbit_1_0.ram_80_0.m0_s 
* net 1150 = rbit_1_0.ram_80_0.m1_s 
* net 1151 = rbit_1_0.ram_79_1.m0_s 
* net 1152 = rbit_1_0.ram_79_1.m1_s 
* net 1153 = rbit_1_0.ram_79_0.m0_s 
* net 1154 = rbit_1_0.ram_79_0.m1_s 
* net 1155 = rbit_1_0.ram_78_1.m0_s 
* net 1156 = rbit_1_0.ram_78_1.m1_s 
* net 1157 = rbit_1_0.ram_78_0.m0_s 
* net 1158 = rbit_1_0.ram_78_0.m1_s 
* net 1159 = rbit_1_0.ram_77_1.m0_s 
* net 1160 = rbit_1_0.ram_77_1.m1_s 
* net 1161 = rbit_1_0.ram_77_0.m0_s 
* net 1162 = rbit_1_0.ram_77_0.m1_s 
* net 1163 = rbit_1_0.ram_76_1.m0_s 
* net 1164 = rbit_1_0.ram_76_1.m1_s 
* net 1165 = rbit_1_0.ram_76_0.m0_s 
* net 1166 = rbit_1_0.ram_76_0.m1_s 
* net 1167 = rbit_1_0.ram_75_1.m0_s 
* net 1168 = rbit_1_0.ram_75_1.m1_s 
* net 1169 = rbit_1_0.ram_75_0.m0_s 
* net 1170 = rbit_1_0.ram_75_0.m1_s 
* net 1171 = rbit_1_0.ram_74_1.m0_s 
* net 1172 = rbit_1_0.ram_74_1.m1_s 
* net 1173 = rbit_1_0.ram_74_0.m0_s 
* net 1174 = rbit_1_0.ram_74_0.m1_s 
* net 1175 = rbit_1_0.ram_73_1.m0_s 
* net 1176 = rbit_1_0.ram_73_1.m1_s 
* net 1177 = rbit_1_0.ram_73_0.m0_s 
* net 1178 = rbit_1_0.ram_73_0.m1_s 
* net 1179 = rbit_1_0.ram_72_1.m0_s 
* net 1180 = rbit_1_0.ram_72_1.m1_s 
* net 1181 = rbit_1_0.ram_72_0.m0_s 
* net 1182 = rbit_1_0.ram_72_0.m1_s 
* net 1183 = rbit_1_0.ram_71_1.m0_s 
* net 1184 = rbit_1_0.ram_71_1.m1_s 
* net 1185 = rbit_1_0.ram_71_0.m0_s 
* net 1186 = rbit_1_0.ram_71_0.m1_s 
* net 1187 = rbit_1_0.ram_70_1.m0_s 
* net 1188 = rbit_1_0.ram_70_1.m1_s 
* net 1189 = rbit_1_0.ram_70_0.m0_s 
* net 1190 = rbit_1_0.ram_70_0.m1_s 
* net 1191 = rbit_1_0.ram_69_1.m0_s 
* net 1192 = rbit_1_0.ram_69_1.m1_s 
* net 1193 = rbit_1_0.ram_69_0.m0_s 
* net 1194 = rbit_1_0.ram_69_0.m1_s 
* net 1195 = rbit_1_0.ram_68_1.m0_s 
* net 1196 = rbit_1_0.ram_68_1.m1_s 
* net 1197 = rbit_1_0.ram_68_0.m0_s 
* net 1198 = rbit_1_0.ram_68_0.m1_s 
* net 1199 = rbit_1_0.ram_67_1.m0_s 
* net 1200 = rbit_1_0.ram_67_1.m1_s 
* net 1201 = rbit_1_0.ram_67_0.m0_s 
* net 1202 = rbit_1_0.ram_67_0.m1_s 
* net 1203 = rbit_1_0.ram_66_1.m0_s 
* net 1204 = rbit_1_0.ram_66_1.m1_s 
* net 1205 = rbit_1_0.ram_66_0.m0_s 
* net 1206 = rbit_1_0.ram_66_0.m1_s 
* net 1207 = rbit_1_0.ram_65_1.m0_s 
* net 1208 = rbit_1_0.ram_65_1.m1_s 
* net 1209 = rbit_1_0.ram_65_0.m0_s 
* net 1210 = rbit_1_0.ram_65_0.m1_s 
* net 1211 = rbit_1_0.ram_64_1.m0_s 
* net 1212 = rbit_1_0.ram_64_1.m1_s 
* net 1213 = rbit_1_0.ram_64_0.m0_s 
* net 1214 = rbit_1_0.ram_64_0.m1_s 
* net 1215 = rbit_1_0.ram_63_1.m0_s 
* net 1216 = rbit_1_0.ram_63_1.m1_s 
* net 1217 = rbit_1_0.ram_63_0.m0_s 
* net 1218 = rbit_1_0.ram_63_0.m1_s 
* net 1219 = rbit_1_0.ram_62_1.m0_s 
* net 1220 = rbit_1_0.ram_62_1.m1_s 
* net 1221 = rbit_1_0.ram_62_0.m0_s 
* net 1222 = rbit_1_0.ram_62_0.m1_s 
* net 1223 = rbit_1_0.ram_61_1.m0_s 
* net 1224 = rbit_1_0.ram_61_1.m1_s 
* net 1225 = rbit_1_0.ram_61_0.m0_s 
* net 1226 = rbit_1_0.ram_61_0.m1_s 
* net 1227 = rbit_1_0.ram_60_1.m0_s 
* net 1228 = rbit_1_0.ram_60_1.m1_s 
* net 1229 = rbit_1_0.ram_60_0.m0_s 
* net 1230 = rbit_1_0.ram_60_0.m1_s 
* net 1231 = rbit_1_0.ram_59_1.m0_s 
* net 1232 = rbit_1_0.ram_59_1.m1_s 
* net 1233 = rbit_1_0.ram_59_0.m0_s 
* net 1234 = rbit_1_0.ram_59_0.m1_s 
* net 1235 = rbit_1_0.ram_58_1.m0_s 
* net 1236 = rbit_1_0.ram_58_1.m1_s 
* net 1237 = rbit_1_0.ram_58_0.m0_s 
* net 1238 = rbit_1_0.ram_58_0.m1_s 
* net 1239 = rbit_1_0.ram_57_1.m0_s 
* net 1240 = rbit_1_0.ram_57_1.m1_s 
* net 1241 = rbit_1_0.ram_57_0.m0_s 
* net 1242 = rbit_1_0.ram_57_0.m1_s 
* net 1243 = rbit_1_0.ram_56_1.m0_s 
* net 1244 = rbit_1_0.ram_56_1.m1_s 
* net 1245 = rbit_1_0.ram_56_0.m0_s 
* net 1246 = rbit_1_0.ram_56_0.m1_s 
* net 1247 = rbit_1_0.ram_55_1.m0_s 
* net 1248 = rbit_1_0.ram_55_1.m1_s 
* net 1249 = rbit_1_0.ram_55_0.m0_s 
* net 1250 = rbit_1_0.ram_55_0.m1_s 
* net 1251 = rbit_1_0.ram_54_1.m0_s 
* net 1252 = rbit_1_0.ram_54_1.m1_s 
* net 1253 = rbit_1_0.ram_54_0.m0_s 
* net 1254 = rbit_1_0.ram_54_0.m1_s 
* net 1255 = rbit_1_0.ram_53_1.m0_s 
* net 1256 = rbit_1_0.ram_53_1.m1_s 
* net 1257 = rbit_1_0.ram_53_0.m0_s 
* net 1258 = rbit_1_0.ram_53_0.m1_s 
* net 1259 = rbit_1_0.ram_52_1.m0_s 
* net 1260 = rbit_1_0.ram_52_1.m1_s 
* net 1261 = rbit_1_0.ram_52_0.m0_s 
* net 1262 = rbit_1_0.ram_52_0.m1_s 
* net 1263 = rbit_1_0.ram_51_1.m0_s 
* net 1264 = rbit_1_0.ram_51_1.m1_s 
* net 1265 = rbit_1_0.ram_51_0.m0_s 
* net 1266 = rbit_1_0.ram_51_0.m1_s 
* net 1267 = rbit_1_0.ram_50_1.m0_s 
* net 1268 = rbit_1_0.ram_50_1.m1_s 
* net 1269 = rbit_1_0.ram_50_0.m0_s 
* net 1270 = rbit_1_0.ram_50_0.m1_s 
* net 1271 = rbit_1_0.ram_49_1.m0_s 
* net 1272 = rbit_1_0.ram_49_1.m1_s 
* net 1273 = rbit_1_0.ram_49_0.m0_s 
* net 1274 = rbit_1_0.ram_49_0.m1_s 
* net 1275 = rbit_1_0.ram_48_1.m0_s 
* net 1276 = rbit_1_0.ram_48_1.m1_s 
* net 1277 = rbit_1_0.ram_48_0.m0_s 
* net 1278 = rbit_1_0.ram_48_0.m1_s 
* net 1279 = rbit_1_0.ram_47_1.m0_s 
* net 1280 = rbit_1_0.ram_47_1.m1_s 
* net 1281 = rbit_1_0.ram_47_0.m0_s 
* net 1282 = rbit_1_0.ram_47_0.m1_s 
* net 1283 = rbit_1_0.ram_46_1.m0_s 
* net 1284 = rbit_1_0.ram_46_1.m1_s 
* net 1285 = rbit_1_0.ram_46_0.m0_s 
* net 1286 = rbit_1_0.ram_46_0.m1_s 
* net 1287 = rbit_1_0.ram_45_1.m0_s 
* net 1288 = rbit_1_0.ram_45_1.m1_s 
* net 1289 = rbit_1_0.ram_45_0.m0_s 
* net 1290 = rbit_1_0.ram_45_0.m1_s 
* net 1291 = rbit_1_0.ram_44_1.m0_s 
* net 1292 = rbit_1_0.ram_44_1.m1_s 
* net 1293 = rbit_1_0.ram_44_0.m0_s 
* net 1294 = rbit_1_0.ram_44_0.m1_s 
* net 1295 = rbit_1_0.ram_43_1.m0_s 
* net 1296 = rbit_1_0.ram_43_1.m1_s 
* net 1297 = rbit_1_0.ram_43_0.m0_s 
* net 1298 = rbit_1_0.ram_43_0.m1_s 
* net 1299 = rbit_1_0.ram_42_1.m0_s 
* net 1300 = rbit_1_0.ram_42_1.m1_s 
* net 1301 = rbit_1_0.ram_42_0.m0_s 
* net 1302 = rbit_1_0.ram_42_0.m1_s 
* net 1303 = rbit_1_0.ram_41_1.m0_s 
* net 1304 = rbit_1_0.ram_41_1.m1_s 
* net 1305 = rbit_1_0.ram_41_0.m0_s 
* net 1306 = rbit_1_0.ram_41_0.m1_s 
* net 1307 = rbit_1_0.ram_40_1.m0_s 
* net 1308 = rbit_1_0.ram_40_1.m1_s 
* net 1309 = rbit_1_0.ram_40_0.m0_s 
* net 1310 = rbit_1_0.ram_40_0.m1_s 
* net 1311 = rbit_1_0.ram_39_1.m0_s 
* net 1312 = rbit_1_0.ram_39_1.m1_s 
* net 1313 = rbit_1_0.ram_39_0.m0_s 
* net 1314 = rbit_1_0.ram_39_0.m1_s 
* net 1315 = rbit_1_0.ram_38_1.m0_s 
* net 1316 = rbit_1_0.ram_38_1.m1_s 
* net 1317 = rbit_1_0.ram_38_0.m0_s 
* net 1318 = rbit_1_0.ram_38_0.m1_s 
* net 1319 = rbit_1_0.ram_37_1.m0_s 
* net 1320 = rbit_1_0.ram_37_1.m1_s 
* net 1321 = rbit_1_0.ram_37_0.m0_s 
* net 1322 = rbit_1_0.ram_37_0.m1_s 
* net 1323 = rbit_1_0.ram_36_1.m0_s 
* net 1324 = rbit_1_0.ram_36_1.m1_s 
* net 1325 = rbit_1_0.ram_36_0.m0_s 
* net 1326 = rbit_1_0.ram_36_0.m1_s 
* net 1327 = rbit_1_0.ram_35_1.m0_s 
* net 1328 = rbit_1_0.ram_35_1.m1_s 
* net 1329 = rbit_1_0.ram_35_0.m0_s 
* net 1330 = rbit_1_0.ram_35_0.m1_s 
* net 1331 = rbit_1_0.ram_34_1.m0_s 
* net 1332 = rbit_1_0.ram_34_1.m1_s 
* net 1333 = rbit_1_0.ram_34_0.m0_s 
* net 1334 = rbit_1_0.ram_34_0.m1_s 
* net 1335 = rbit_1_0.ram_33_1.m0_s 
* net 1336 = rbit_1_0.ram_33_1.m1_s 
* net 1337 = rbit_1_0.ram_33_0.m0_s 
* net 1338 = rbit_1_0.ram_33_0.m1_s 
* net 1339 = rbit_1_0.ram_32_1.m0_s 
* net 1340 = rbit_1_0.ram_32_1.m1_s 
* net 1341 = rbit_1_0.ram_32_0.m0_s 
* net 1342 = rbit_1_0.ram_32_0.m1_s 
* net 1343 = rbit_1_0.ram_31_1.m0_s 
* net 1344 = rbit_1_0.ram_31_1.m1_s 
* net 1345 = rbit_1_0.ram_31_0.m0_s 
* net 1346 = rbit_1_0.ram_31_0.m1_s 
* net 1347 = rbit_1_0.ram_30_1.m0_s 
* net 1348 = rbit_1_0.ram_30_1.m1_s 
* net 1349 = rbit_1_0.ram_30_0.m0_s 
* net 1350 = rbit_1_0.ram_30_0.m1_s 
* net 1351 = rbit_1_0.ram_29_1.m0_s 
* net 1352 = rbit_1_0.ram_29_1.m1_s 
* net 1353 = rbit_1_0.ram_29_0.m0_s 
* net 1354 = rbit_1_0.ram_29_0.m1_s 
* net 1355 = rbit_1_0.ram_28_1.m0_s 
* net 1356 = rbit_1_0.ram_28_1.m1_s 
* net 1357 = rbit_1_0.ram_28_0.m0_s 
* net 1358 = rbit_1_0.ram_28_0.m1_s 
* net 1359 = rbit_1_0.ram_27_1.m0_s 
* net 1360 = rbit_1_0.ram_27_1.m1_s 
* net 1361 = rbit_1_0.ram_27_0.m0_s 
* net 1362 = rbit_1_0.ram_27_0.m1_s 
* net 1363 = rbit_1_0.ram_26_1.m0_s 
* net 1364 = rbit_1_0.ram_26_1.m1_s 
* net 1365 = rbit_1_0.ram_26_0.m0_s 
* net 1366 = rbit_1_0.ram_26_0.m1_s 
* net 1367 = rbit_1_0.ram_25_1.m0_s 
* net 1368 = rbit_1_0.ram_25_1.m1_s 
* net 1369 = rbit_1_0.ram_25_0.m0_s 
* net 1370 = rbit_1_0.ram_25_0.m1_s 
* net 1371 = rbit_1_0.ram_24_1.m0_s 
* net 1372 = rbit_1_0.ram_24_1.m1_s 
* net 1373 = rbit_1_0.ram_24_0.m0_s 
* net 1374 = rbit_1_0.ram_24_0.m1_s 
* net 1375 = rbit_1_0.ram_23_1.m0_s 
* net 1376 = rbit_1_0.ram_23_1.m1_s 
* net 1377 = rbit_1_0.ram_23_0.m0_s 
* net 1378 = rbit_1_0.ram_23_0.m1_s 
* net 1379 = rbit_1_0.ram_22_1.m0_s 
* net 1380 = rbit_1_0.ram_22_1.m1_s 
* net 1381 = rbit_1_0.ram_22_0.m0_s 
* net 1382 = rbit_1_0.ram_22_0.m1_s 
* net 1383 = rbit_1_0.ram_21_1.m0_s 
* net 1384 = rbit_1_0.ram_21_1.m1_s 
* net 1385 = rbit_1_0.ram_21_0.m0_s 
* net 1386 = rbit_1_0.ram_21_0.m1_s 
* net 1387 = rbit_1_0.ram_20_1.m0_s 
* net 1388 = rbit_1_0.ram_20_1.m1_s 
* net 1389 = rbit_1_0.ram_20_0.m0_s 
* net 1390 = rbit_1_0.ram_20_0.m1_s 
* net 1391 = rbit_1_0.ram_19_1.m0_s 
* net 1392 = rbit_1_0.ram_19_1.m1_s 
* net 1393 = rbit_1_0.ram_19_0.m0_s 
* net 1394 = rbit_1_0.ram_19_0.m1_s 
* net 1395 = rbit_1_0.ram_18_1.m0_s 
* net 1396 = rbit_1_0.ram_18_1.m1_s 
* net 1397 = rbit_1_0.ram_18_0.m0_s 
* net 1398 = rbit_1_0.ram_18_0.m1_s 
* net 1399 = rbit_1_0.ram_17_1.m0_s 
* net 1400 = rbit_1_0.ram_17_1.m1_s 
* net 1401 = rbit_1_0.ram_17_0.m0_s 
* net 1402 = rbit_1_0.ram_17_0.m1_s 
* net 1403 = rbit_1_0.ram_16_1.m0_s 
* net 1404 = rbit_1_0.ram_16_1.m1_s 
* net 1405 = rbit_1_0.ram_16_0.m0_s 
* net 1406 = rbit_1_0.ram_16_0.m1_s 
* net 1407 = rbit_1_0.ram_15_1.m0_s 
* net 1408 = rbit_1_0.ram_15_1.m1_s 
* net 1409 = rbit_1_0.ram_15_0.m0_s 
* net 1410 = rbit_1_0.ram_15_0.m1_s 
* net 1411 = rbit_1_0.ram_14_1.m0_s 
* net 1412 = rbit_1_0.ram_14_1.m1_s 
* net 1413 = rbit_1_0.ram_14_0.m0_s 
* net 1414 = rbit_1_0.ram_14_0.m1_s 
* net 1415 = rbit_1_0.ram_13_1.m0_s 
* net 1416 = rbit_1_0.ram_13_1.m1_s 
* net 1417 = rbit_1_0.ram_13_0.m0_s 
* net 1418 = rbit_1_0.ram_13_0.m1_s 
* net 1419 = rbit_1_0.ram_12_1.m0_s 
* net 1420 = rbit_1_0.ram_12_1.m1_s 
* net 1421 = rbit_1_0.ram_12_0.m0_s 
* net 1422 = rbit_1_0.ram_12_0.m1_s 
* net 1423 = rbit_1_0.ram_11_1.m0_s 
* net 1424 = rbit_1_0.ram_11_1.m1_s 
* net 1425 = rbit_1_0.ram_11_0.m0_s 
* net 1426 = rbit_1_0.ram_11_0.m1_s 
* net 1427 = rbit_1_0.ram_10_1.m0_s 
* net 1428 = rbit_1_0.ram_10_1.m1_s 
* net 1429 = rbit_1_0.ram_10_0.m0_s 
* net 1430 = rbit_1_0.ram_10_0.m1_s 
* net 1431 = rbit_1_0.ram_9_1.m0_s 
* net 1432 = rbit_1_0.ram_9_1.m1_s 
* net 1433 = rbit_1_0.ram_9_0.m0_s 
* net 1434 = rbit_1_0.ram_9_0.m1_s 
* net 1435 = rbit_1_0.ram_8_1.m0_s 
* net 1436 = rbit_1_0.ram_8_1.m1_s 
* net 1437 = rbit_1_0.ram_8_0.m0_s 
* net 1438 = rbit_1_0.ram_8_0.m1_s 
* net 1439 = rbit_1_0.ram_7_1.m0_s 
* net 1440 = rbit_1_0.ram_7_1.m1_s 
* net 1441 = rbit_1_0.ram_7_0.m0_s 
* net 1442 = rbit_1_0.ram_7_0.m1_s 
* net 1443 = rbit_1_0.ram_6_1.m0_s 
* net 1444 = rbit_1_0.ram_6_1.m1_s 
* net 1445 = rbit_1_0.ram_6_0.m0_s 
* net 1446 = rbit_1_0.ram_6_0.m1_s 
* net 1447 = rbit_1_0.ram_5_1.m0_s 
* net 1448 = rbit_1_0.ram_5_1.m1_s 
* net 1449 = rbit_1_0.ram_5_0.m0_s 
* net 1450 = rbit_1_0.ram_5_0.m1_s 
* net 1451 = rbit_1_0.ram_4_1.m0_s 
* net 1452 = rbit_1_0.ram_4_1.m1_s 
* net 1453 = rbit_1_0.ram_4_0.m0_s 
* net 1454 = rbit_1_0.ram_4_0.m1_s 
* net 1455 = rbit_1_0.ram_3_1.m0_s 
* net 1456 = rbit_1_0.ram_3_1.m1_s 
* net 1457 = rbit_1_0.ram_3_0.m0_s 
* net 1458 = rbit_1_0.ram_3_0.m1_s 
* net 1459 = rbit_1_0.ram_2_1.m0_s 
* net 1460 = rbit_1_0.ram_2_1.m1_s 
* net 1461 = rbit_1_0.ram_2_0.m0_s 
* net 1462 = rbit_1_0.ram_2_0.m1_s 
* net 1463 = rbit_1_0.ram_1_1.m0_s 
* net 1464 = rbit_1_0.ram_1_1.m1_s 
* net 1465 = rbit_1_0.ram_1_0.m0_s 
* net 1466 = rbit_1_0.ram_1_0.m1_s 
* net 1467 = rbit_1_0.ram_0_1.m0_s 
* net 1468 = rbit_1_0.ram_0_1.m1_s 
* net 1469 = rbit_1_0.ram_0_0.m0_s 
* net 1470 = rbit_1_0.ram_0_0.m1_s 
* net 1471 = mbk_sig134 
* net 1472 = mbk_sig110 
* net 1473 = mbk_sig160 
* net 1474 = mbk_sig111 
* net 1475 = mbk_sig181 
* net 1476 = mbk_sig11 
* net 1477 = mbk_sig8 
* net 1478 = mbk_sig67 
* net 1479 = mbk_sig99 
* net 1480 = mbk_sig91 
* net 1481 = mbk_sig83 
* net 1482 = rbit_2_0.ram_127_1.m0_s 
* net 1483 = rbit_2_0.ram_127_1.m1_s 
* net 1484 = rbit_2_0.ram_127_0.m0_s 
* net 1485 = rbit_2_0.ram_127_0.m1_s 
* net 1486 = rbit_2_0.ram_126_1.m0_s 
* net 1487 = rbit_2_0.ram_126_1.m1_s 
* net 1488 = rbit_2_0.ram_126_0.m0_s 
* net 1489 = rbit_2_0.ram_126_0.m1_s 
* net 1490 = rbit_2_0.ram_125_1.m0_s 
* net 1491 = rbit_2_0.ram_125_1.m1_s 
* net 1492 = rbit_2_0.ram_125_0.m0_s 
* net 1493 = rbit_2_0.ram_125_0.m1_s 
* net 1494 = rbit_2_0.ram_124_1.m0_s 
* net 1495 = rbit_2_0.ram_124_1.m1_s 
* net 1496 = rbit_2_0.ram_124_0.m0_s 
* net 1497 = rbit_2_0.ram_124_0.m1_s 
* net 1498 = rbit_2_0.ram_123_1.m0_s 
* net 1499 = rbit_2_0.ram_123_1.m1_s 
* net 1500 = rbit_2_0.ram_123_0.m0_s 
* net 1501 = rbit_2_0.ram_123_0.m1_s 
* net 1502 = rbit_2_0.ram_122_1.m0_s 
* net 1503 = rbit_2_0.ram_122_1.m1_s 
* net 1504 = rbit_2_0.ram_122_0.m0_s 
* net 1505 = rbit_2_0.ram_122_0.m1_s 
* net 1506 = rbit_2_0.ram_121_1.m0_s 
* net 1507 = rbit_2_0.ram_121_1.m1_s 
* net 1508 = rbit_2_0.ram_121_0.m0_s 
* net 1509 = rbit_2_0.ram_121_0.m1_s 
* net 1510 = rbit_2_0.ram_120_1.m0_s 
* net 1511 = rbit_2_0.ram_120_1.m1_s 
* net 1512 = rbit_2_0.ram_120_0.m0_s 
* net 1513 = rbit_2_0.ram_120_0.m1_s 
* net 1514 = rbit_2_0.ram_119_1.m0_s 
* net 1515 = rbit_2_0.ram_119_1.m1_s 
* net 1516 = rbit_2_0.ram_119_0.m0_s 
* net 1517 = rbit_2_0.ram_119_0.m1_s 
* net 1518 = rbit_2_0.ram_118_1.m0_s 
* net 1519 = rbit_2_0.ram_118_1.m1_s 
* net 1520 = rbit_2_0.ram_118_0.m0_s 
* net 1521 = rbit_2_0.ram_118_0.m1_s 
* net 1522 = rbit_2_0.ram_117_1.m0_s 
* net 1523 = rbit_2_0.ram_117_1.m1_s 
* net 1524 = rbit_2_0.ram_117_0.m0_s 
* net 1525 = rbit_2_0.ram_117_0.m1_s 
* net 1526 = rbit_2_0.ram_116_1.m0_s 
* net 1527 = rbit_2_0.ram_116_1.m1_s 
* net 1528 = rbit_2_0.ram_116_0.m0_s 
* net 1529 = rbit_2_0.ram_116_0.m1_s 
* net 1530 = rbit_2_0.ram_115_1.m0_s 
* net 1531 = rbit_2_0.ram_115_1.m1_s 
* net 1532 = rbit_2_0.ram_115_0.m0_s 
* net 1533 = rbit_2_0.ram_115_0.m1_s 
* net 1534 = rbit_2_0.ram_114_1.m0_s 
* net 1535 = rbit_2_0.ram_114_1.m1_s 
* net 1536 = rbit_2_0.ram_114_0.m0_s 
* net 1537 = rbit_2_0.ram_114_0.m1_s 
* net 1538 = rbit_2_0.ram_113_1.m0_s 
* net 1539 = rbit_2_0.ram_113_1.m1_s 
* net 1540 = rbit_2_0.ram_113_0.m0_s 
* net 1541 = rbit_2_0.ram_113_0.m1_s 
* net 1542 = rbit_2_0.ram_112_1.m0_s 
* net 1543 = rbit_2_0.ram_112_1.m1_s 
* net 1544 = rbit_2_0.ram_112_0.m0_s 
* net 1545 = rbit_2_0.ram_112_0.m1_s 
* net 1546 = rbit_2_0.ram_111_1.m0_s 
* net 1547 = rbit_2_0.ram_111_1.m1_s 
* net 1548 = rbit_2_0.ram_111_0.m0_s 
* net 1549 = rbit_2_0.ram_111_0.m1_s 
* net 1550 = rbit_2_0.ram_110_1.m0_s 
* net 1551 = rbit_2_0.ram_110_1.m1_s 
* net 1552 = rbit_2_0.ram_110_0.m0_s 
* net 1553 = rbit_2_0.ram_110_0.m1_s 
* net 1554 = rbit_2_0.ram_109_1.m0_s 
* net 1555 = rbit_2_0.ram_109_1.m1_s 
* net 1556 = rbit_2_0.ram_109_0.m0_s 
* net 1557 = rbit_2_0.ram_109_0.m1_s 
* net 1558 = rbit_2_0.ram_108_1.m0_s 
* net 1559 = rbit_2_0.ram_108_1.m1_s 
* net 1560 = rbit_2_0.ram_108_0.m0_s 
* net 1561 = rbit_2_0.ram_108_0.m1_s 
* net 1562 = rbit_2_0.ram_107_1.m0_s 
* net 1563 = rbit_2_0.ram_107_1.m1_s 
* net 1564 = rbit_2_0.ram_107_0.m0_s 
* net 1565 = rbit_2_0.ram_107_0.m1_s 
* net 1566 = rbit_2_0.ram_106_1.m0_s 
* net 1567 = rbit_2_0.ram_106_1.m1_s 
* net 1568 = rbit_2_0.ram_106_0.m0_s 
* net 1569 = rbit_2_0.ram_106_0.m1_s 
* net 1570 = rbit_2_0.ram_105_1.m0_s 
* net 1571 = rbit_2_0.ram_105_1.m1_s 
* net 1572 = rbit_2_0.ram_105_0.m0_s 
* net 1573 = rbit_2_0.ram_105_0.m1_s 
* net 1574 = rbit_2_0.ram_104_1.m0_s 
* net 1575 = rbit_2_0.ram_104_1.m1_s 
* net 1576 = rbit_2_0.ram_104_0.m0_s 
* net 1577 = rbit_2_0.ram_104_0.m1_s 
* net 1578 = rbit_2_0.ram_103_1.m0_s 
* net 1579 = rbit_2_0.ram_103_1.m1_s 
* net 1580 = rbit_2_0.ram_103_0.m0_s 
* net 1581 = rbit_2_0.ram_103_0.m1_s 
* net 1582 = rbit_2_0.ram_102_1.m0_s 
* net 1583 = rbit_2_0.ram_102_1.m1_s 
* net 1584 = rbit_2_0.ram_102_0.m0_s 
* net 1585 = rbit_2_0.ram_102_0.m1_s 
* net 1586 = rbit_2_0.ram_101_1.m0_s 
* net 1587 = rbit_2_0.ram_101_1.m1_s 
* net 1588 = rbit_2_0.ram_101_0.m0_s 
* net 1589 = rbit_2_0.ram_101_0.m1_s 
* net 1590 = rbit_2_0.ram_100_1.m0_s 
* net 1591 = rbit_2_0.ram_100_1.m1_s 
* net 1592 = rbit_2_0.ram_100_0.m0_s 
* net 1593 = rbit_2_0.ram_100_0.m1_s 
* net 1594 = rbit_2_0.ram_99_1.m0_s 
* net 1595 = rbit_2_0.ram_99_1.m1_s 
* net 1596 = rbit_2_0.ram_99_0.m0_s 
* net 1597 = rbit_2_0.ram_99_0.m1_s 
* net 1598 = rbit_2_0.ram_98_1.m0_s 
* net 1599 = rbit_2_0.ram_98_1.m1_s 
* net 1600 = rbit_2_0.ram_98_0.m0_s 
* net 1601 = rbit_2_0.ram_98_0.m1_s 
* net 1602 = rbit_2_0.ram_97_1.m0_s 
* net 1603 = rbit_2_0.ram_97_1.m1_s 
* net 1604 = rbit_2_0.ram_97_0.m0_s 
* net 1605 = rbit_2_0.ram_97_0.m1_s 
* net 1606 = rbit_2_0.ram_96_1.m0_s 
* net 1607 = rbit_2_0.ram_96_1.m1_s 
* net 1608 = rbit_2_0.ram_96_0.m0_s 
* net 1609 = rbit_2_0.ram_96_0.m1_s 
* net 1610 = rbit_2_0.ram_95_1.m0_s 
* net 1611 = rbit_2_0.ram_95_1.m1_s 
* net 1612 = rbit_2_0.ram_95_0.m0_s 
* net 1613 = rbit_2_0.ram_95_0.m1_s 
* net 1614 = rbit_2_0.ram_94_1.m0_s 
* net 1615 = rbit_2_0.ram_94_1.m1_s 
* net 1616 = rbit_2_0.ram_94_0.m0_s 
* net 1617 = rbit_2_0.ram_94_0.m1_s 
* net 1618 = rbit_2_0.ram_93_1.m0_s 
* net 1619 = rbit_2_0.ram_93_1.m1_s 
* net 1620 = rbit_2_0.ram_93_0.m0_s 
* net 1621 = rbit_2_0.ram_93_0.m1_s 
* net 1622 = rbit_2_0.ram_92_1.m0_s 
* net 1623 = rbit_2_0.ram_92_1.m1_s 
* net 1624 = rbit_2_0.ram_92_0.m0_s 
* net 1625 = rbit_2_0.ram_92_0.m1_s 
* net 1626 = rbit_2_0.ram_91_1.m0_s 
* net 1627 = rbit_2_0.ram_91_1.m1_s 
* net 1628 = rbit_2_0.ram_91_0.m0_s 
* net 1629 = rbit_2_0.ram_91_0.m1_s 
* net 1630 = rbit_2_0.ram_90_1.m0_s 
* net 1631 = rbit_2_0.ram_90_1.m1_s 
* net 1632 = rbit_2_0.ram_90_0.m0_s 
* net 1633 = rbit_2_0.ram_90_0.m1_s 
* net 1634 = rbit_2_0.ram_89_1.m0_s 
* net 1635 = rbit_2_0.ram_89_1.m1_s 
* net 1636 = rbit_2_0.ram_89_0.m0_s 
* net 1637 = rbit_2_0.ram_89_0.m1_s 
* net 1638 = rbit_2_0.ram_88_1.m0_s 
* net 1639 = rbit_2_0.ram_88_1.m1_s 
* net 1640 = rbit_2_0.ram_88_0.m0_s 
* net 1641 = rbit_2_0.ram_88_0.m1_s 
* net 1642 = rbit_2_0.ram_87_1.m0_s 
* net 1643 = rbit_2_0.ram_87_1.m1_s 
* net 1644 = rbit_2_0.ram_87_0.m0_s 
* net 1645 = rbit_2_0.ram_87_0.m1_s 
* net 1646 = rbit_2_0.ram_86_1.m0_s 
* net 1647 = rbit_2_0.ram_86_1.m1_s 
* net 1648 = rbit_2_0.ram_86_0.m0_s 
* net 1649 = rbit_2_0.ram_86_0.m1_s 
* net 1650 = rbit_2_0.ram_85_1.m0_s 
* net 1651 = rbit_2_0.ram_85_1.m1_s 
* net 1652 = rbit_2_0.ram_85_0.m0_s 
* net 1653 = rbit_2_0.ram_85_0.m1_s 
* net 1654 = rbit_2_0.ram_84_1.m0_s 
* net 1655 = rbit_2_0.ram_84_1.m1_s 
* net 1656 = rbit_2_0.ram_84_0.m0_s 
* net 1657 = rbit_2_0.ram_84_0.m1_s 
* net 1658 = rbit_2_0.ram_83_1.m0_s 
* net 1659 = rbit_2_0.ram_83_1.m1_s 
* net 1660 = rbit_2_0.ram_83_0.m0_s 
* net 1661 = rbit_2_0.ram_83_0.m1_s 
* net 1662 = rbit_2_0.ram_82_1.m0_s 
* net 1663 = rbit_2_0.ram_82_1.m1_s 
* net 1664 = rbit_2_0.ram_82_0.m0_s 
* net 1665 = rbit_2_0.ram_82_0.m1_s 
* net 1666 = rbit_2_0.ram_81_1.m0_s 
* net 1667 = rbit_2_0.ram_81_1.m1_s 
* net 1668 = rbit_2_0.ram_81_0.m0_s 
* net 1669 = rbit_2_0.ram_81_0.m1_s 
* net 1670 = rbit_2_0.ram_80_1.m0_s 
* net 1671 = rbit_2_0.ram_80_1.m1_s 
* net 1672 = rbit_2_0.ram_80_0.m0_s 
* net 1673 = rbit_2_0.ram_80_0.m1_s 
* net 1674 = rbit_2_0.ram_79_1.m0_s 
* net 1675 = rbit_2_0.ram_79_1.m1_s 
* net 1676 = rbit_2_0.ram_79_0.m0_s 
* net 1677 = rbit_2_0.ram_79_0.m1_s 
* net 1678 = rbit_2_0.ram_78_1.m0_s 
* net 1679 = rbit_2_0.ram_78_1.m1_s 
* net 1680 = rbit_2_0.ram_78_0.m0_s 
* net 1681 = rbit_2_0.ram_78_0.m1_s 
* net 1682 = rbit_2_0.ram_77_1.m0_s 
* net 1683 = rbit_2_0.ram_77_1.m1_s 
* net 1684 = rbit_2_0.ram_77_0.m0_s 
* net 1685 = rbit_2_0.ram_77_0.m1_s 
* net 1686 = rbit_2_0.ram_76_1.m0_s 
* net 1687 = rbit_2_0.ram_76_1.m1_s 
* net 1688 = rbit_2_0.ram_76_0.m0_s 
* net 1689 = rbit_2_0.ram_76_0.m1_s 
* net 1690 = rbit_2_0.ram_75_1.m0_s 
* net 1691 = rbit_2_0.ram_75_1.m1_s 
* net 1692 = rbit_2_0.ram_75_0.m0_s 
* net 1693 = rbit_2_0.ram_75_0.m1_s 
* net 1694 = rbit_2_0.ram_74_1.m0_s 
* net 1695 = rbit_2_0.ram_74_1.m1_s 
* net 1696 = rbit_2_0.ram_74_0.m0_s 
* net 1697 = rbit_2_0.ram_74_0.m1_s 
* net 1698 = rbit_2_0.ram_73_1.m0_s 
* net 1699 = rbit_2_0.ram_73_1.m1_s 
* net 1700 = rbit_2_0.ram_73_0.m0_s 
* net 1701 = rbit_2_0.ram_73_0.m1_s 
* net 1702 = rbit_2_0.ram_72_1.m0_s 
* net 1703 = rbit_2_0.ram_72_1.m1_s 
* net 1704 = rbit_2_0.ram_72_0.m0_s 
* net 1705 = rbit_2_0.ram_72_0.m1_s 
* net 1706 = rbit_2_0.ram_71_1.m0_s 
* net 1707 = rbit_2_0.ram_71_1.m1_s 
* net 1708 = rbit_2_0.ram_71_0.m0_s 
* net 1709 = rbit_2_0.ram_71_0.m1_s 
* net 1710 = rbit_2_0.ram_70_1.m0_s 
* net 1711 = rbit_2_0.ram_70_1.m1_s 
* net 1712 = rbit_2_0.ram_70_0.m0_s 
* net 1713 = rbit_2_0.ram_70_0.m1_s 
* net 1714 = rbit_2_0.ram_69_1.m0_s 
* net 1715 = rbit_2_0.ram_69_1.m1_s 
* net 1716 = rbit_2_0.ram_69_0.m0_s 
* net 1717 = rbit_2_0.ram_69_0.m1_s 
* net 1718 = rbit_2_0.ram_68_1.m0_s 
* net 1719 = rbit_2_0.ram_68_1.m1_s 
* net 1720 = rbit_2_0.ram_68_0.m0_s 
* net 1721 = rbit_2_0.ram_68_0.m1_s 
* net 1722 = rbit_2_0.ram_67_1.m0_s 
* net 1723 = rbit_2_0.ram_67_1.m1_s 
* net 1724 = rbit_2_0.ram_67_0.m0_s 
* net 1725 = rbit_2_0.ram_67_0.m1_s 
* net 1726 = rbit_2_0.ram_66_1.m0_s 
* net 1727 = rbit_2_0.ram_66_1.m1_s 
* net 1728 = rbit_2_0.ram_66_0.m0_s 
* net 1729 = rbit_2_0.ram_66_0.m1_s 
* net 1730 = rbit_2_0.ram_65_1.m0_s 
* net 1731 = rbit_2_0.ram_65_1.m1_s 
* net 1732 = rbit_2_0.ram_65_0.m0_s 
* net 1733 = rbit_2_0.ram_65_0.m1_s 
* net 1734 = rbit_2_0.ram_64_1.m0_s 
* net 1735 = rbit_2_0.ram_64_1.m1_s 
* net 1736 = rbit_2_0.ram_64_0.m0_s 
* net 1737 = rbit_2_0.ram_64_0.m1_s 
* net 1738 = rbit_2_0.ram_63_1.m0_s 
* net 1739 = rbit_2_0.ram_63_1.m1_s 
* net 1740 = rbit_2_0.ram_63_0.m0_s 
* net 1741 = rbit_2_0.ram_63_0.m1_s 
* net 1742 = rbit_2_0.ram_62_1.m0_s 
* net 1743 = rbit_2_0.ram_62_1.m1_s 
* net 1744 = rbit_2_0.ram_62_0.m0_s 
* net 1745 = rbit_2_0.ram_62_0.m1_s 
* net 1746 = rbit_2_0.ram_61_1.m0_s 
* net 1747 = rbit_2_0.ram_61_1.m1_s 
* net 1748 = rbit_2_0.ram_61_0.m0_s 
* net 1749 = rbit_2_0.ram_61_0.m1_s 
* net 1750 = rbit_2_0.ram_60_1.m0_s 
* net 1751 = rbit_2_0.ram_60_1.m1_s 
* net 1752 = rbit_2_0.ram_60_0.m0_s 
* net 1753 = rbit_2_0.ram_60_0.m1_s 
* net 1754 = rbit_2_0.ram_59_1.m0_s 
* net 1755 = rbit_2_0.ram_59_1.m1_s 
* net 1756 = rbit_2_0.ram_59_0.m0_s 
* net 1757 = rbit_2_0.ram_59_0.m1_s 
* net 1758 = rbit_2_0.ram_58_1.m0_s 
* net 1759 = rbit_2_0.ram_58_1.m1_s 
* net 1760 = rbit_2_0.ram_58_0.m0_s 
* net 1761 = rbit_2_0.ram_58_0.m1_s 
* net 1762 = rbit_2_0.ram_57_1.m0_s 
* net 1763 = rbit_2_0.ram_57_1.m1_s 
* net 1764 = rbit_2_0.ram_57_0.m0_s 
* net 1765 = rbit_2_0.ram_57_0.m1_s 
* net 1766 = rbit_2_0.ram_56_1.m0_s 
* net 1767 = rbit_2_0.ram_56_1.m1_s 
* net 1768 = rbit_2_0.ram_56_0.m0_s 
* net 1769 = rbit_2_0.ram_56_0.m1_s 
* net 1770 = rbit_2_0.ram_55_1.m0_s 
* net 1771 = rbit_2_0.ram_55_1.m1_s 
* net 1772 = rbit_2_0.ram_55_0.m0_s 
* net 1773 = rbit_2_0.ram_55_0.m1_s 
* net 1774 = rbit_2_0.ram_54_1.m0_s 
* net 1775 = rbit_2_0.ram_54_1.m1_s 
* net 1776 = rbit_2_0.ram_54_0.m0_s 
* net 1777 = rbit_2_0.ram_54_0.m1_s 
* net 1778 = rbit_2_0.ram_53_1.m0_s 
* net 1779 = rbit_2_0.ram_53_1.m1_s 
* net 1780 = rbit_2_0.ram_53_0.m0_s 
* net 1781 = rbit_2_0.ram_53_0.m1_s 
* net 1782 = rbit_2_0.ram_52_1.m0_s 
* net 1783 = rbit_2_0.ram_52_1.m1_s 
* net 1784 = rbit_2_0.ram_52_0.m0_s 
* net 1785 = rbit_2_0.ram_52_0.m1_s 
* net 1786 = rbit_2_0.ram_51_1.m0_s 
* net 1787 = rbit_2_0.ram_51_1.m1_s 
* net 1788 = rbit_2_0.ram_51_0.m0_s 
* net 1789 = rbit_2_0.ram_51_0.m1_s 
* net 1790 = rbit_2_0.ram_50_1.m0_s 
* net 1791 = rbit_2_0.ram_50_1.m1_s 
* net 1792 = rbit_2_0.ram_50_0.m0_s 
* net 1793 = rbit_2_0.ram_50_0.m1_s 
* net 1794 = rbit_2_0.ram_49_1.m0_s 
* net 1795 = rbit_2_0.ram_49_1.m1_s 
* net 1796 = rbit_2_0.ram_49_0.m0_s 
* net 1797 = rbit_2_0.ram_49_0.m1_s 
* net 1798 = rbit_2_0.ram_48_1.m0_s 
* net 1799 = rbit_2_0.ram_48_1.m1_s 
* net 1800 = rbit_2_0.ram_48_0.m0_s 
* net 1801 = rbit_2_0.ram_48_0.m1_s 
* net 1802 = rbit_2_0.ram_47_1.m0_s 
* net 1803 = rbit_2_0.ram_47_1.m1_s 
* net 1804 = rbit_2_0.ram_47_0.m0_s 
* net 1805 = rbit_2_0.ram_47_0.m1_s 
* net 1806 = rbit_2_0.ram_46_1.m0_s 
* net 1807 = rbit_2_0.ram_46_1.m1_s 
* net 1808 = rbit_2_0.ram_46_0.m0_s 
* net 1809 = rbit_2_0.ram_46_0.m1_s 
* net 1810 = rbit_2_0.ram_45_1.m0_s 
* net 1811 = rbit_2_0.ram_45_1.m1_s 
* net 1812 = rbit_2_0.ram_45_0.m0_s 
* net 1813 = rbit_2_0.ram_45_0.m1_s 
* net 1814 = rbit_2_0.ram_44_1.m0_s 
* net 1815 = rbit_2_0.ram_44_1.m1_s 
* net 1816 = rbit_2_0.ram_44_0.m0_s 
* net 1817 = rbit_2_0.ram_44_0.m1_s 
* net 1818 = rbit_2_0.ram_43_1.m0_s 
* net 1819 = rbit_2_0.ram_43_1.m1_s 
* net 1820 = rbit_2_0.ram_43_0.m0_s 
* net 1821 = rbit_2_0.ram_43_0.m1_s 
* net 1822 = rbit_2_0.ram_42_1.m0_s 
* net 1823 = rbit_2_0.ram_42_1.m1_s 
* net 1824 = rbit_2_0.ram_42_0.m0_s 
* net 1825 = rbit_2_0.ram_42_0.m1_s 
* net 1826 = rbit_2_0.ram_41_1.m0_s 
* net 1827 = rbit_2_0.ram_41_1.m1_s 
* net 1828 = rbit_2_0.ram_41_0.m0_s 
* net 1829 = rbit_2_0.ram_41_0.m1_s 
* net 1830 = rbit_2_0.ram_40_1.m0_s 
* net 1831 = rbit_2_0.ram_40_1.m1_s 
* net 1832 = rbit_2_0.ram_40_0.m0_s 
* net 1833 = rbit_2_0.ram_40_0.m1_s 
* net 1834 = rbit_2_0.ram_39_1.m0_s 
* net 1835 = rbit_2_0.ram_39_1.m1_s 
* net 1836 = rbit_2_0.ram_39_0.m0_s 
* net 1837 = rbit_2_0.ram_39_0.m1_s 
* net 1838 = rbit_2_0.ram_38_1.m0_s 
* net 1839 = rbit_2_0.ram_38_1.m1_s 
* net 1840 = rbit_2_0.ram_38_0.m0_s 
* net 1841 = rbit_2_0.ram_38_0.m1_s 
* net 1842 = rbit_2_0.ram_37_1.m0_s 
* net 1843 = rbit_2_0.ram_37_1.m1_s 
* net 1844 = rbit_2_0.ram_37_0.m0_s 
* net 1845 = rbit_2_0.ram_37_0.m1_s 
* net 1846 = rbit_2_0.ram_36_1.m0_s 
* net 1847 = rbit_2_0.ram_36_1.m1_s 
* net 1848 = rbit_2_0.ram_36_0.m0_s 
* net 1849 = rbit_2_0.ram_36_0.m1_s 
* net 1850 = rbit_2_0.ram_35_1.m0_s 
* net 1851 = rbit_2_0.ram_35_1.m1_s 
* net 1852 = rbit_2_0.ram_35_0.m0_s 
* net 1853 = rbit_2_0.ram_35_0.m1_s 
* net 1854 = rbit_2_0.ram_34_1.m0_s 
* net 1855 = rbit_2_0.ram_34_1.m1_s 
* net 1856 = rbit_2_0.ram_34_0.m0_s 
* net 1857 = rbit_2_0.ram_34_0.m1_s 
* net 1858 = rbit_2_0.ram_33_1.m0_s 
* net 1859 = rbit_2_0.ram_33_1.m1_s 
* net 1860 = rbit_2_0.ram_33_0.m0_s 
* net 1861 = rbit_2_0.ram_33_0.m1_s 
* net 1862 = rbit_2_0.ram_32_1.m0_s 
* net 1863 = rbit_2_0.ram_32_1.m1_s 
* net 1864 = rbit_2_0.ram_32_0.m0_s 
* net 1865 = rbit_2_0.ram_32_0.m1_s 
* net 1866 = rbit_2_0.ram_31_1.m0_s 
* net 1867 = rbit_2_0.ram_31_1.m1_s 
* net 1868 = rbit_2_0.ram_31_0.m0_s 
* net 1869 = rbit_2_0.ram_31_0.m1_s 
* net 1870 = rbit_2_0.ram_30_1.m0_s 
* net 1871 = rbit_2_0.ram_30_1.m1_s 
* net 1872 = rbit_2_0.ram_30_0.m0_s 
* net 1873 = rbit_2_0.ram_30_0.m1_s 
* net 1874 = rbit_2_0.ram_29_1.m0_s 
* net 1875 = rbit_2_0.ram_29_1.m1_s 
* net 1876 = rbit_2_0.ram_29_0.m0_s 
* net 1877 = rbit_2_0.ram_29_0.m1_s 
* net 1878 = rbit_2_0.ram_28_1.m0_s 
* net 1879 = rbit_2_0.ram_28_1.m1_s 
* net 1880 = rbit_2_0.ram_28_0.m0_s 
* net 1881 = rbit_2_0.ram_28_0.m1_s 
* net 1882 = rbit_2_0.ram_27_1.m0_s 
* net 1883 = rbit_2_0.ram_27_1.m1_s 
* net 1884 = rbit_2_0.ram_27_0.m0_s 
* net 1885 = rbit_2_0.ram_27_0.m1_s 
* net 1886 = rbit_2_0.ram_26_1.m0_s 
* net 1887 = rbit_2_0.ram_26_1.m1_s 
* net 1888 = rbit_2_0.ram_26_0.m0_s 
* net 1889 = rbit_2_0.ram_26_0.m1_s 
* net 1890 = rbit_2_0.ram_25_1.m0_s 
* net 1891 = rbit_2_0.ram_25_1.m1_s 
* net 1892 = rbit_2_0.ram_25_0.m0_s 
* net 1893 = rbit_2_0.ram_25_0.m1_s 
* net 1894 = rbit_2_0.ram_24_1.m0_s 
* net 1895 = rbit_2_0.ram_24_1.m1_s 
* net 1896 = rbit_2_0.ram_24_0.m0_s 
* net 1897 = rbit_2_0.ram_24_0.m1_s 
* net 1898 = rbit_2_0.ram_23_1.m0_s 
* net 1899 = rbit_2_0.ram_23_1.m1_s 
* net 1900 = rbit_2_0.ram_23_0.m0_s 
* net 1901 = rbit_2_0.ram_23_0.m1_s 
* net 1902 = rbit_2_0.ram_22_1.m0_s 
* net 1903 = rbit_2_0.ram_22_1.m1_s 
* net 1904 = rbit_2_0.ram_22_0.m0_s 
* net 1905 = rbit_2_0.ram_22_0.m1_s 
* net 1906 = rbit_2_0.ram_21_1.m0_s 
* net 1907 = rbit_2_0.ram_21_1.m1_s 
* net 1908 = rbit_2_0.ram_21_0.m0_s 
* net 1909 = rbit_2_0.ram_21_0.m1_s 
* net 1910 = rbit_2_0.ram_20_1.m0_s 
* net 1911 = rbit_2_0.ram_20_1.m1_s 
* net 1912 = rbit_2_0.ram_20_0.m0_s 
* net 1913 = rbit_2_0.ram_20_0.m1_s 
* net 1914 = rbit_2_0.ram_19_1.m0_s 
* net 1915 = rbit_2_0.ram_19_1.m1_s 
* net 1916 = rbit_2_0.ram_19_0.m0_s 
* net 1917 = rbit_2_0.ram_19_0.m1_s 
* net 1918 = rbit_2_0.ram_18_1.m0_s 
* net 1919 = rbit_2_0.ram_18_1.m1_s 
* net 1920 = rbit_2_0.ram_18_0.m0_s 
* net 1921 = rbit_2_0.ram_18_0.m1_s 
* net 1922 = rbit_2_0.ram_17_1.m0_s 
* net 1923 = rbit_2_0.ram_17_1.m1_s 
* net 1924 = rbit_2_0.ram_17_0.m0_s 
* net 1925 = rbit_2_0.ram_17_0.m1_s 
* net 1926 = rbit_2_0.ram_16_1.m0_s 
* net 1927 = rbit_2_0.ram_16_1.m1_s 
* net 1928 = rbit_2_0.ram_16_0.m0_s 
* net 1929 = rbit_2_0.ram_16_0.m1_s 
* net 1930 = rbit_2_0.ram_15_1.m0_s 
* net 1931 = rbit_2_0.ram_15_1.m1_s 
* net 1932 = rbit_2_0.ram_15_0.m0_s 
* net 1933 = rbit_2_0.ram_15_0.m1_s 
* net 1934 = rbit_2_0.ram_14_1.m0_s 
* net 1935 = rbit_2_0.ram_14_1.m1_s 
* net 1936 = rbit_2_0.ram_14_0.m0_s 
* net 1937 = rbit_2_0.ram_14_0.m1_s 
* net 1938 = rbit_2_0.ram_13_1.m0_s 
* net 1939 = rbit_2_0.ram_13_1.m1_s 
* net 1940 = rbit_2_0.ram_13_0.m0_s 
* net 1941 = rbit_2_0.ram_13_0.m1_s 
* net 1942 = rbit_2_0.ram_12_1.m0_s 
* net 1943 = rbit_2_0.ram_12_1.m1_s 
* net 1944 = rbit_2_0.ram_12_0.m0_s 
* net 1945 = rbit_2_0.ram_12_0.m1_s 
* net 1946 = rbit_2_0.ram_11_1.m0_s 
* net 1947 = rbit_2_0.ram_11_1.m1_s 
* net 1948 = rbit_2_0.ram_11_0.m0_s 
* net 1949 = rbit_2_0.ram_11_0.m1_s 
* net 1950 = rbit_2_0.ram_10_1.m0_s 
* net 1951 = rbit_2_0.ram_10_1.m1_s 
* net 1952 = rbit_2_0.ram_10_0.m0_s 
* net 1953 = rbit_2_0.ram_10_0.m1_s 
* net 1954 = rbit_2_0.ram_9_1.m0_s 
* net 1955 = rbit_2_0.ram_9_1.m1_s 
* net 1956 = rbit_2_0.ram_9_0.m0_s 
* net 1957 = rbit_2_0.ram_9_0.m1_s 
* net 1958 = rbit_2_0.ram_8_1.m0_s 
* net 1959 = rbit_2_0.ram_8_1.m1_s 
* net 1960 = rbit_2_0.ram_8_0.m0_s 
* net 1961 = rbit_2_0.ram_8_0.m1_s 
* net 1962 = rbit_2_0.ram_7_1.m0_s 
* net 1963 = rbit_2_0.ram_7_1.m1_s 
* net 1964 = rbit_2_0.ram_7_0.m0_s 
* net 1965 = rbit_2_0.ram_7_0.m1_s 
* net 1966 = rbit_2_0.ram_6_1.m0_s 
* net 1967 = rbit_2_0.ram_6_1.m1_s 
* net 1968 = rbit_2_0.ram_6_0.m0_s 
* net 1969 = rbit_2_0.ram_6_0.m1_s 
* net 1970 = rbit_2_0.ram_5_1.m0_s 
* net 1971 = rbit_2_0.ram_5_1.m1_s 
* net 1972 = rbit_2_0.ram_5_0.m0_s 
* net 1973 = rbit_2_0.ram_5_0.m1_s 
* net 1974 = rbit_2_0.ram_4_1.m0_s 
* net 1975 = rbit_2_0.ram_4_1.m1_s 
* net 1976 = rbit_2_0.ram_4_0.m0_s 
* net 1977 = rbit_2_0.ram_4_0.m1_s 
* net 1978 = rbit_2_0.ram_3_1.m0_s 
* net 1979 = rbit_2_0.ram_3_1.m1_s 
* net 1980 = rbit_2_0.ram_3_0.m0_s 
* net 1981 = rbit_2_0.ram_3_0.m1_s 
* net 1982 = rbit_2_0.ram_2_1.m0_s 
* net 1983 = rbit_2_0.ram_2_1.m1_s 
* net 1984 = rbit_2_0.ram_2_0.m0_s 
* net 1985 = rbit_2_0.ram_2_0.m1_s 
* net 1986 = rbit_2_0.ram_1_1.m0_s 
* net 1987 = rbit_2_0.ram_1_1.m1_s 
* net 1988 = rbit_2_0.ram_1_0.m0_s 
* net 1989 = rbit_2_0.ram_1_0.m1_s 
* net 1990 = rbit_2_0.ram_0_1.m0_s 
* net 1991 = rbit_2_0.ram_0_1.m1_s 
* net 1992 = rbit_2_0.ram_0_0.m0_s 
* net 1993 = rbit_2_0.ram_0_0.m1_s 
* net 1994 = mbk_sig137 
* net 1995 = mbk_sig113 
* net 1996 = mbk_sig162 
* net 1997 = mbk_sig112 
* net 1998 = mbk_sig182 
* net 1999 = mbk_sig16 
* net 2000 = mbk_sig14 
* net 2001 = mbk_sig68 
* net 2002 = mbk_sig100 
* net 2003 = mbk_sig92 
* net 2004 = mbk_sig84 
* net 2005 = rbit_3_0.ram_127_1.m0_s 
* net 2006 = rbit_3_0.ram_127_1.m1_s 
* net 2007 = rbit_3_0.ram_127_0.m0_s 
* net 2008 = rbit_3_0.ram_127_0.m1_s 
* net 2009 = rbit_3_0.ram_126_1.m0_s 
* net 2010 = rbit_3_0.ram_126_1.m1_s 
* net 2011 = rbit_3_0.ram_126_0.m0_s 
* net 2012 = rbit_3_0.ram_126_0.m1_s 
* net 2013 = rbit_3_0.ram_125_1.m0_s 
* net 2014 = rbit_3_0.ram_125_1.m1_s 
* net 2015 = rbit_3_0.ram_125_0.m0_s 
* net 2016 = rbit_3_0.ram_125_0.m1_s 
* net 2017 = rbit_3_0.ram_124_1.m0_s 
* net 2018 = rbit_3_0.ram_124_1.m1_s 
* net 2019 = rbit_3_0.ram_124_0.m0_s 
* net 2020 = rbit_3_0.ram_124_0.m1_s 
* net 2021 = rbit_3_0.ram_123_1.m0_s 
* net 2022 = rbit_3_0.ram_123_1.m1_s 
* net 2023 = rbit_3_0.ram_123_0.m0_s 
* net 2024 = rbit_3_0.ram_123_0.m1_s 
* net 2025 = rbit_3_0.ram_122_1.m0_s 
* net 2026 = rbit_3_0.ram_122_1.m1_s 
* net 2027 = rbit_3_0.ram_122_0.m0_s 
* net 2028 = rbit_3_0.ram_122_0.m1_s 
* net 2029 = rbit_3_0.ram_121_1.m0_s 
* net 2030 = rbit_3_0.ram_121_1.m1_s 
* net 2031 = rbit_3_0.ram_121_0.m0_s 
* net 2032 = rbit_3_0.ram_121_0.m1_s 
* net 2033 = rbit_3_0.ram_120_1.m0_s 
* net 2034 = rbit_3_0.ram_120_1.m1_s 
* net 2035 = rbit_3_0.ram_120_0.m0_s 
* net 2036 = rbit_3_0.ram_120_0.m1_s 
* net 2037 = rbit_3_0.ram_119_1.m0_s 
* net 2038 = rbit_3_0.ram_119_1.m1_s 
* net 2039 = rbit_3_0.ram_119_0.m0_s 
* net 2040 = rbit_3_0.ram_119_0.m1_s 
* net 2041 = rbit_3_0.ram_118_1.m0_s 
* net 2042 = rbit_3_0.ram_118_1.m1_s 
* net 2043 = rbit_3_0.ram_118_0.m0_s 
* net 2044 = rbit_3_0.ram_118_0.m1_s 
* net 2045 = rbit_3_0.ram_117_1.m0_s 
* net 2046 = rbit_3_0.ram_117_1.m1_s 
* net 2047 = rbit_3_0.ram_117_0.m0_s 
* net 2048 = rbit_3_0.ram_117_0.m1_s 
* net 2049 = rbit_3_0.ram_116_1.m0_s 
* net 2050 = rbit_3_0.ram_116_1.m1_s 
* net 2051 = rbit_3_0.ram_116_0.m0_s 
* net 2052 = rbit_3_0.ram_116_0.m1_s 
* net 2053 = rbit_3_0.ram_115_1.m0_s 
* net 2054 = rbit_3_0.ram_115_1.m1_s 
* net 2055 = rbit_3_0.ram_115_0.m0_s 
* net 2056 = rbit_3_0.ram_115_0.m1_s 
* net 2057 = rbit_3_0.ram_114_1.m0_s 
* net 2058 = rbit_3_0.ram_114_1.m1_s 
* net 2059 = rbit_3_0.ram_114_0.m0_s 
* net 2060 = rbit_3_0.ram_114_0.m1_s 
* net 2061 = rbit_3_0.ram_113_1.m0_s 
* net 2062 = rbit_3_0.ram_113_1.m1_s 
* net 2063 = rbit_3_0.ram_113_0.m0_s 
* net 2064 = rbit_3_0.ram_113_0.m1_s 
* net 2065 = rbit_3_0.ram_112_1.m0_s 
* net 2066 = rbit_3_0.ram_112_1.m1_s 
* net 2067 = rbit_3_0.ram_112_0.m0_s 
* net 2068 = rbit_3_0.ram_112_0.m1_s 
* net 2069 = rbit_3_0.ram_111_1.m0_s 
* net 2070 = rbit_3_0.ram_111_1.m1_s 
* net 2071 = rbit_3_0.ram_111_0.m0_s 
* net 2072 = rbit_3_0.ram_111_0.m1_s 
* net 2073 = rbit_3_0.ram_110_1.m0_s 
* net 2074 = rbit_3_0.ram_110_1.m1_s 
* net 2075 = rbit_3_0.ram_110_0.m0_s 
* net 2076 = rbit_3_0.ram_110_0.m1_s 
* net 2077 = rbit_3_0.ram_109_1.m0_s 
* net 2078 = rbit_3_0.ram_109_1.m1_s 
* net 2079 = rbit_3_0.ram_109_0.m0_s 
* net 2080 = rbit_3_0.ram_109_0.m1_s 
* net 2081 = rbit_3_0.ram_108_1.m0_s 
* net 2082 = rbit_3_0.ram_108_1.m1_s 
* net 2083 = rbit_3_0.ram_108_0.m0_s 
* net 2084 = rbit_3_0.ram_108_0.m1_s 
* net 2085 = rbit_3_0.ram_107_1.m0_s 
* net 2086 = rbit_3_0.ram_107_1.m1_s 
* net 2087 = rbit_3_0.ram_107_0.m0_s 
* net 2088 = rbit_3_0.ram_107_0.m1_s 
* net 2089 = rbit_3_0.ram_106_1.m0_s 
* net 2090 = rbit_3_0.ram_106_1.m1_s 
* net 2091 = rbit_3_0.ram_106_0.m0_s 
* net 2092 = rbit_3_0.ram_106_0.m1_s 
* net 2093 = rbit_3_0.ram_105_1.m0_s 
* net 2094 = rbit_3_0.ram_105_1.m1_s 
* net 2095 = rbit_3_0.ram_105_0.m0_s 
* net 2096 = rbit_3_0.ram_105_0.m1_s 
* net 2097 = rbit_3_0.ram_104_1.m0_s 
* net 2098 = rbit_3_0.ram_104_1.m1_s 
* net 2099 = rbit_3_0.ram_104_0.m0_s 
* net 2100 = rbit_3_0.ram_104_0.m1_s 
* net 2101 = rbit_3_0.ram_103_1.m0_s 
* net 2102 = rbit_3_0.ram_103_1.m1_s 
* net 2103 = rbit_3_0.ram_103_0.m0_s 
* net 2104 = rbit_3_0.ram_103_0.m1_s 
* net 2105 = rbit_3_0.ram_102_1.m0_s 
* net 2106 = rbit_3_0.ram_102_1.m1_s 
* net 2107 = rbit_3_0.ram_102_0.m0_s 
* net 2108 = rbit_3_0.ram_102_0.m1_s 
* net 2109 = rbit_3_0.ram_101_1.m0_s 
* net 2110 = rbit_3_0.ram_101_1.m1_s 
* net 2111 = rbit_3_0.ram_101_0.m0_s 
* net 2112 = rbit_3_0.ram_101_0.m1_s 
* net 2113 = rbit_3_0.ram_100_1.m0_s 
* net 2114 = rbit_3_0.ram_100_1.m1_s 
* net 2115 = rbit_3_0.ram_100_0.m0_s 
* net 2116 = rbit_3_0.ram_100_0.m1_s 
* net 2117 = rbit_3_0.ram_99_1.m0_s 
* net 2118 = rbit_3_0.ram_99_1.m1_s 
* net 2119 = rbit_3_0.ram_99_0.m0_s 
* net 2120 = rbit_3_0.ram_99_0.m1_s 
* net 2121 = rbit_3_0.ram_98_1.m0_s 
* net 2122 = rbit_3_0.ram_98_1.m1_s 
* net 2123 = rbit_3_0.ram_98_0.m0_s 
* net 2124 = rbit_3_0.ram_98_0.m1_s 
* net 2125 = rbit_3_0.ram_97_1.m0_s 
* net 2126 = rbit_3_0.ram_97_1.m1_s 
* net 2127 = rbit_3_0.ram_97_0.m0_s 
* net 2128 = rbit_3_0.ram_97_0.m1_s 
* net 2129 = rbit_3_0.ram_96_1.m0_s 
* net 2130 = rbit_3_0.ram_96_1.m1_s 
* net 2131 = rbit_3_0.ram_96_0.m0_s 
* net 2132 = rbit_3_0.ram_96_0.m1_s 
* net 2133 = rbit_3_0.ram_95_1.m0_s 
* net 2134 = rbit_3_0.ram_95_1.m1_s 
* net 2135 = rbit_3_0.ram_95_0.m0_s 
* net 2136 = rbit_3_0.ram_95_0.m1_s 
* net 2137 = rbit_3_0.ram_94_1.m0_s 
* net 2138 = rbit_3_0.ram_94_1.m1_s 
* net 2139 = rbit_3_0.ram_94_0.m0_s 
* net 2140 = rbit_3_0.ram_94_0.m1_s 
* net 2141 = rbit_3_0.ram_93_1.m0_s 
* net 2142 = rbit_3_0.ram_93_1.m1_s 
* net 2143 = rbit_3_0.ram_93_0.m0_s 
* net 2144 = rbit_3_0.ram_93_0.m1_s 
* net 2145 = rbit_3_0.ram_92_1.m0_s 
* net 2146 = rbit_3_0.ram_92_1.m1_s 
* net 2147 = rbit_3_0.ram_92_0.m0_s 
* net 2148 = rbit_3_0.ram_92_0.m1_s 
* net 2149 = rbit_3_0.ram_91_1.m0_s 
* net 2150 = rbit_3_0.ram_91_1.m1_s 
* net 2151 = rbit_3_0.ram_91_0.m0_s 
* net 2152 = rbit_3_0.ram_91_0.m1_s 
* net 2153 = rbit_3_0.ram_90_1.m0_s 
* net 2154 = rbit_3_0.ram_90_1.m1_s 
* net 2155 = rbit_3_0.ram_90_0.m0_s 
* net 2156 = rbit_3_0.ram_90_0.m1_s 
* net 2157 = rbit_3_0.ram_89_1.m0_s 
* net 2158 = rbit_3_0.ram_89_1.m1_s 
* net 2159 = rbit_3_0.ram_89_0.m0_s 
* net 2160 = rbit_3_0.ram_89_0.m1_s 
* net 2161 = rbit_3_0.ram_88_1.m0_s 
* net 2162 = rbit_3_0.ram_88_1.m1_s 
* net 2163 = rbit_3_0.ram_88_0.m0_s 
* net 2164 = rbit_3_0.ram_88_0.m1_s 
* net 2165 = rbit_3_0.ram_87_1.m0_s 
* net 2166 = rbit_3_0.ram_87_1.m1_s 
* net 2167 = rbit_3_0.ram_87_0.m0_s 
* net 2168 = rbit_3_0.ram_87_0.m1_s 
* net 2169 = rbit_3_0.ram_86_1.m0_s 
* net 2170 = rbit_3_0.ram_86_1.m1_s 
* net 2171 = rbit_3_0.ram_86_0.m0_s 
* net 2172 = rbit_3_0.ram_86_0.m1_s 
* net 2173 = rbit_3_0.ram_85_1.m0_s 
* net 2174 = rbit_3_0.ram_85_1.m1_s 
* net 2175 = rbit_3_0.ram_85_0.m0_s 
* net 2176 = rbit_3_0.ram_85_0.m1_s 
* net 2177 = rbit_3_0.ram_84_1.m0_s 
* net 2178 = rbit_3_0.ram_84_1.m1_s 
* net 2179 = rbit_3_0.ram_84_0.m0_s 
* net 2180 = rbit_3_0.ram_84_0.m1_s 
* net 2181 = rbit_3_0.ram_83_1.m0_s 
* net 2182 = rbit_3_0.ram_83_1.m1_s 
* net 2183 = rbit_3_0.ram_83_0.m0_s 
* net 2184 = rbit_3_0.ram_83_0.m1_s 
* net 2185 = rbit_3_0.ram_82_1.m0_s 
* net 2186 = rbit_3_0.ram_82_1.m1_s 
* net 2187 = rbit_3_0.ram_82_0.m0_s 
* net 2188 = rbit_3_0.ram_82_0.m1_s 
* net 2189 = rbit_3_0.ram_81_1.m0_s 
* net 2190 = rbit_3_0.ram_81_1.m1_s 
* net 2191 = rbit_3_0.ram_81_0.m0_s 
* net 2192 = rbit_3_0.ram_81_0.m1_s 
* net 2193 = rbit_3_0.ram_80_1.m0_s 
* net 2194 = rbit_3_0.ram_80_1.m1_s 
* net 2195 = rbit_3_0.ram_80_0.m0_s 
* net 2196 = rbit_3_0.ram_80_0.m1_s 
* net 2197 = rbit_3_0.ram_79_1.m0_s 
* net 2198 = rbit_3_0.ram_79_1.m1_s 
* net 2199 = rbit_3_0.ram_79_0.m0_s 
* net 2200 = rbit_3_0.ram_79_0.m1_s 
* net 2201 = rbit_3_0.ram_78_1.m0_s 
* net 2202 = rbit_3_0.ram_78_1.m1_s 
* net 2203 = rbit_3_0.ram_78_0.m0_s 
* net 2204 = rbit_3_0.ram_78_0.m1_s 
* net 2205 = rbit_3_0.ram_77_1.m0_s 
* net 2206 = rbit_3_0.ram_77_1.m1_s 
* net 2207 = rbit_3_0.ram_77_0.m0_s 
* net 2208 = rbit_3_0.ram_77_0.m1_s 
* net 2209 = rbit_3_0.ram_76_1.m0_s 
* net 2210 = rbit_3_0.ram_76_1.m1_s 
* net 2211 = rbit_3_0.ram_76_0.m0_s 
* net 2212 = rbit_3_0.ram_76_0.m1_s 
* net 2213 = rbit_3_0.ram_75_1.m0_s 
* net 2214 = rbit_3_0.ram_75_1.m1_s 
* net 2215 = rbit_3_0.ram_75_0.m0_s 
* net 2216 = rbit_3_0.ram_75_0.m1_s 
* net 2217 = rbit_3_0.ram_74_1.m0_s 
* net 2218 = rbit_3_0.ram_74_1.m1_s 
* net 2219 = rbit_3_0.ram_74_0.m0_s 
* net 2220 = rbit_3_0.ram_74_0.m1_s 
* net 2221 = rbit_3_0.ram_73_1.m0_s 
* net 2222 = rbit_3_0.ram_73_1.m1_s 
* net 2223 = rbit_3_0.ram_73_0.m0_s 
* net 2224 = rbit_3_0.ram_73_0.m1_s 
* net 2225 = rbit_3_0.ram_72_1.m0_s 
* net 2226 = rbit_3_0.ram_72_1.m1_s 
* net 2227 = rbit_3_0.ram_72_0.m0_s 
* net 2228 = rbit_3_0.ram_72_0.m1_s 
* net 2229 = rbit_3_0.ram_71_1.m0_s 
* net 2230 = rbit_3_0.ram_71_1.m1_s 
* net 2231 = rbit_3_0.ram_71_0.m0_s 
* net 2232 = rbit_3_0.ram_71_0.m1_s 
* net 2233 = rbit_3_0.ram_70_1.m0_s 
* net 2234 = rbit_3_0.ram_70_1.m1_s 
* net 2235 = rbit_3_0.ram_70_0.m0_s 
* net 2236 = rbit_3_0.ram_70_0.m1_s 
* net 2237 = rbit_3_0.ram_69_1.m0_s 
* net 2238 = rbit_3_0.ram_69_1.m1_s 
* net 2239 = rbit_3_0.ram_69_0.m0_s 
* net 2240 = rbit_3_0.ram_69_0.m1_s 
* net 2241 = rbit_3_0.ram_68_1.m0_s 
* net 2242 = rbit_3_0.ram_68_1.m1_s 
* net 2243 = rbit_3_0.ram_68_0.m0_s 
* net 2244 = rbit_3_0.ram_68_0.m1_s 
* net 2245 = rbit_3_0.ram_67_1.m0_s 
* net 2246 = rbit_3_0.ram_67_1.m1_s 
* net 2247 = rbit_3_0.ram_67_0.m0_s 
* net 2248 = rbit_3_0.ram_67_0.m1_s 
* net 2249 = rbit_3_0.ram_66_1.m0_s 
* net 2250 = rbit_3_0.ram_66_1.m1_s 
* net 2251 = rbit_3_0.ram_66_0.m0_s 
* net 2252 = rbit_3_0.ram_66_0.m1_s 
* net 2253 = rbit_3_0.ram_65_1.m0_s 
* net 2254 = rbit_3_0.ram_65_1.m1_s 
* net 2255 = rbit_3_0.ram_65_0.m0_s 
* net 2256 = rbit_3_0.ram_65_0.m1_s 
* net 2257 = rbit_3_0.ram_64_1.m0_s 
* net 2258 = rbit_3_0.ram_64_1.m1_s 
* net 2259 = rbit_3_0.ram_64_0.m0_s 
* net 2260 = rbit_3_0.ram_64_0.m1_s 
* net 2261 = rbit_3_0.ram_63_1.m0_s 
* net 2262 = rbit_3_0.ram_63_1.m1_s 
* net 2263 = rbit_3_0.ram_63_0.m0_s 
* net 2264 = rbit_3_0.ram_63_0.m1_s 
* net 2265 = rbit_3_0.ram_62_1.m0_s 
* net 2266 = rbit_3_0.ram_62_1.m1_s 
* net 2267 = rbit_3_0.ram_62_0.m0_s 
* net 2268 = rbit_3_0.ram_62_0.m1_s 
* net 2269 = rbit_3_0.ram_61_1.m0_s 
* net 2270 = rbit_3_0.ram_61_1.m1_s 
* net 2271 = rbit_3_0.ram_61_0.m0_s 
* net 2272 = rbit_3_0.ram_61_0.m1_s 
* net 2273 = rbit_3_0.ram_60_1.m0_s 
* net 2274 = rbit_3_0.ram_60_1.m1_s 
* net 2275 = rbit_3_0.ram_60_0.m0_s 
* net 2276 = rbit_3_0.ram_60_0.m1_s 
* net 2277 = rbit_3_0.ram_59_1.m0_s 
* net 2278 = rbit_3_0.ram_59_1.m1_s 
* net 2279 = rbit_3_0.ram_59_0.m0_s 
* net 2280 = rbit_3_0.ram_59_0.m1_s 
* net 2281 = rbit_3_0.ram_58_1.m0_s 
* net 2282 = rbit_3_0.ram_58_1.m1_s 
* net 2283 = rbit_3_0.ram_58_0.m0_s 
* net 2284 = rbit_3_0.ram_58_0.m1_s 
* net 2285 = rbit_3_0.ram_57_1.m0_s 
* net 2286 = rbit_3_0.ram_57_1.m1_s 
* net 2287 = rbit_3_0.ram_57_0.m0_s 
* net 2288 = rbit_3_0.ram_57_0.m1_s 
* net 2289 = rbit_3_0.ram_56_1.m0_s 
* net 2290 = rbit_3_0.ram_56_1.m1_s 
* net 2291 = rbit_3_0.ram_56_0.m0_s 
* net 2292 = rbit_3_0.ram_56_0.m1_s 
* net 2293 = rbit_3_0.ram_55_1.m0_s 
* net 2294 = rbit_3_0.ram_55_1.m1_s 
* net 2295 = rbit_3_0.ram_55_0.m0_s 
* net 2296 = rbit_3_0.ram_55_0.m1_s 
* net 2297 = rbit_3_0.ram_54_1.m0_s 
* net 2298 = rbit_3_0.ram_54_1.m1_s 
* net 2299 = rbit_3_0.ram_54_0.m0_s 
* net 2300 = rbit_3_0.ram_54_0.m1_s 
* net 2301 = rbit_3_0.ram_53_1.m0_s 
* net 2302 = rbit_3_0.ram_53_1.m1_s 
* net 2303 = rbit_3_0.ram_53_0.m0_s 
* net 2304 = rbit_3_0.ram_53_0.m1_s 
* net 2305 = rbit_3_0.ram_52_1.m0_s 
* net 2306 = rbit_3_0.ram_52_1.m1_s 
* net 2307 = rbit_3_0.ram_52_0.m0_s 
* net 2308 = rbit_3_0.ram_52_0.m1_s 
* net 2309 = rbit_3_0.ram_51_1.m0_s 
* net 2310 = rbit_3_0.ram_51_1.m1_s 
* net 2311 = rbit_3_0.ram_51_0.m0_s 
* net 2312 = rbit_3_0.ram_51_0.m1_s 
* net 2313 = rbit_3_0.ram_50_1.m0_s 
* net 2314 = rbit_3_0.ram_50_1.m1_s 
* net 2315 = rbit_3_0.ram_50_0.m0_s 
* net 2316 = rbit_3_0.ram_50_0.m1_s 
* net 2317 = rbit_3_0.ram_49_1.m0_s 
* net 2318 = rbit_3_0.ram_49_1.m1_s 
* net 2319 = rbit_3_0.ram_49_0.m0_s 
* net 2320 = rbit_3_0.ram_49_0.m1_s 
* net 2321 = rbit_3_0.ram_48_1.m0_s 
* net 2322 = rbit_3_0.ram_48_1.m1_s 
* net 2323 = rbit_3_0.ram_48_0.m0_s 
* net 2324 = rbit_3_0.ram_48_0.m1_s 
* net 2325 = rbit_3_0.ram_47_1.m0_s 
* net 2326 = rbit_3_0.ram_47_1.m1_s 
* net 2327 = rbit_3_0.ram_47_0.m0_s 
* net 2328 = rbit_3_0.ram_47_0.m1_s 
* net 2329 = rbit_3_0.ram_46_1.m0_s 
* net 2330 = rbit_3_0.ram_46_1.m1_s 
* net 2331 = rbit_3_0.ram_46_0.m0_s 
* net 2332 = rbit_3_0.ram_46_0.m1_s 
* net 2333 = rbit_3_0.ram_45_1.m0_s 
* net 2334 = rbit_3_0.ram_45_1.m1_s 
* net 2335 = rbit_3_0.ram_45_0.m0_s 
* net 2336 = rbit_3_0.ram_45_0.m1_s 
* net 2337 = rbit_3_0.ram_44_1.m0_s 
* net 2338 = rbit_3_0.ram_44_1.m1_s 
* net 2339 = rbit_3_0.ram_44_0.m0_s 
* net 2340 = rbit_3_0.ram_44_0.m1_s 
* net 2341 = rbit_3_0.ram_43_1.m0_s 
* net 2342 = rbit_3_0.ram_43_1.m1_s 
* net 2343 = rbit_3_0.ram_43_0.m0_s 
* net 2344 = rbit_3_0.ram_43_0.m1_s 
* net 2345 = rbit_3_0.ram_42_1.m0_s 
* net 2346 = rbit_3_0.ram_42_1.m1_s 
* net 2347 = rbit_3_0.ram_42_0.m0_s 
* net 2348 = rbit_3_0.ram_42_0.m1_s 
* net 2349 = rbit_3_0.ram_41_1.m0_s 
* net 2350 = rbit_3_0.ram_41_1.m1_s 
* net 2351 = rbit_3_0.ram_41_0.m0_s 
* net 2352 = rbit_3_0.ram_41_0.m1_s 
* net 2353 = rbit_3_0.ram_40_1.m0_s 
* net 2354 = rbit_3_0.ram_40_1.m1_s 
* net 2355 = rbit_3_0.ram_40_0.m0_s 
* net 2356 = rbit_3_0.ram_40_0.m1_s 
* net 2357 = rbit_3_0.ram_39_1.m0_s 
* net 2358 = rbit_3_0.ram_39_1.m1_s 
* net 2359 = rbit_3_0.ram_39_0.m0_s 
* net 2360 = rbit_3_0.ram_39_0.m1_s 
* net 2361 = rbit_3_0.ram_38_1.m0_s 
* net 2362 = rbit_3_0.ram_38_1.m1_s 
* net 2363 = rbit_3_0.ram_38_0.m0_s 
* net 2364 = rbit_3_0.ram_38_0.m1_s 
* net 2365 = rbit_3_0.ram_37_1.m0_s 
* net 2366 = rbit_3_0.ram_37_1.m1_s 
* net 2367 = rbit_3_0.ram_37_0.m0_s 
* net 2368 = rbit_3_0.ram_37_0.m1_s 
* net 2369 = rbit_3_0.ram_36_1.m0_s 
* net 2370 = rbit_3_0.ram_36_1.m1_s 
* net 2371 = rbit_3_0.ram_36_0.m0_s 
* net 2372 = rbit_3_0.ram_36_0.m1_s 
* net 2373 = rbit_3_0.ram_35_1.m0_s 
* net 2374 = rbit_3_0.ram_35_1.m1_s 
* net 2375 = rbit_3_0.ram_35_0.m0_s 
* net 2376 = rbit_3_0.ram_35_0.m1_s 
* net 2377 = rbit_3_0.ram_34_1.m0_s 
* net 2378 = rbit_3_0.ram_34_1.m1_s 
* net 2379 = rbit_3_0.ram_34_0.m0_s 
* net 2380 = rbit_3_0.ram_34_0.m1_s 
* net 2381 = rbit_3_0.ram_33_1.m0_s 
* net 2382 = rbit_3_0.ram_33_1.m1_s 
* net 2383 = rbit_3_0.ram_33_0.m0_s 
* net 2384 = rbit_3_0.ram_33_0.m1_s 
* net 2385 = rbit_3_0.ram_32_1.m0_s 
* net 2386 = rbit_3_0.ram_32_1.m1_s 
* net 2387 = rbit_3_0.ram_32_0.m0_s 
* net 2388 = rbit_3_0.ram_32_0.m1_s 
* net 2389 = rbit_3_0.ram_31_1.m0_s 
* net 2390 = rbit_3_0.ram_31_1.m1_s 
* net 2391 = rbit_3_0.ram_31_0.m0_s 
* net 2392 = rbit_3_0.ram_31_0.m1_s 
* net 2393 = rbit_3_0.ram_30_1.m0_s 
* net 2394 = rbit_3_0.ram_30_1.m1_s 
* net 2395 = rbit_3_0.ram_30_0.m0_s 
* net 2396 = rbit_3_0.ram_30_0.m1_s 
* net 2397 = rbit_3_0.ram_29_1.m0_s 
* net 2398 = rbit_3_0.ram_29_1.m1_s 
* net 2399 = rbit_3_0.ram_29_0.m0_s 
* net 2400 = rbit_3_0.ram_29_0.m1_s 
* net 2401 = rbit_3_0.ram_28_1.m0_s 
* net 2402 = rbit_3_0.ram_28_1.m1_s 
* net 2403 = rbit_3_0.ram_28_0.m0_s 
* net 2404 = rbit_3_0.ram_28_0.m1_s 
* net 2405 = rbit_3_0.ram_27_1.m0_s 
* net 2406 = rbit_3_0.ram_27_1.m1_s 
* net 2407 = rbit_3_0.ram_27_0.m0_s 
* net 2408 = rbit_3_0.ram_27_0.m1_s 
* net 2409 = rbit_3_0.ram_26_1.m0_s 
* net 2410 = rbit_3_0.ram_26_1.m1_s 
* net 2411 = rbit_3_0.ram_26_0.m0_s 
* net 2412 = rbit_3_0.ram_26_0.m1_s 
* net 2413 = rbit_3_0.ram_25_1.m0_s 
* net 2414 = rbit_3_0.ram_25_1.m1_s 
* net 2415 = rbit_3_0.ram_25_0.m0_s 
* net 2416 = rbit_3_0.ram_25_0.m1_s 
* net 2417 = rbit_3_0.ram_24_1.m0_s 
* net 2418 = rbit_3_0.ram_24_1.m1_s 
* net 2419 = rbit_3_0.ram_24_0.m0_s 
* net 2420 = rbit_3_0.ram_24_0.m1_s 
* net 2421 = rbit_3_0.ram_23_1.m0_s 
* net 2422 = rbit_3_0.ram_23_1.m1_s 
* net 2423 = rbit_3_0.ram_23_0.m0_s 
* net 2424 = rbit_3_0.ram_23_0.m1_s 
* net 2425 = rbit_3_0.ram_22_1.m0_s 
* net 2426 = rbit_3_0.ram_22_1.m1_s 
* net 2427 = rbit_3_0.ram_22_0.m0_s 
* net 2428 = rbit_3_0.ram_22_0.m1_s 
* net 2429 = rbit_3_0.ram_21_1.m0_s 
* net 2430 = rbit_3_0.ram_21_1.m1_s 
* net 2431 = rbit_3_0.ram_21_0.m0_s 
* net 2432 = rbit_3_0.ram_21_0.m1_s 
* net 2433 = rbit_3_0.ram_20_1.m0_s 
* net 2434 = rbit_3_0.ram_20_1.m1_s 
* net 2435 = rbit_3_0.ram_20_0.m0_s 
* net 2436 = rbit_3_0.ram_20_0.m1_s 
* net 2437 = rbit_3_0.ram_19_1.m0_s 
* net 2438 = rbit_3_0.ram_19_1.m1_s 
* net 2439 = rbit_3_0.ram_19_0.m0_s 
* net 2440 = rbit_3_0.ram_19_0.m1_s 
* net 2441 = rbit_3_0.ram_18_1.m0_s 
* net 2442 = rbit_3_0.ram_18_1.m1_s 
* net 2443 = rbit_3_0.ram_18_0.m0_s 
* net 2444 = rbit_3_0.ram_18_0.m1_s 
* net 2445 = rbit_3_0.ram_17_1.m0_s 
* net 2446 = rbit_3_0.ram_17_1.m1_s 
* net 2447 = rbit_3_0.ram_17_0.m0_s 
* net 2448 = rbit_3_0.ram_17_0.m1_s 
* net 2449 = rbit_3_0.ram_16_1.m0_s 
* net 2450 = rbit_3_0.ram_16_1.m1_s 
* net 2451 = rbit_3_0.ram_16_0.m0_s 
* net 2452 = rbit_3_0.ram_16_0.m1_s 
* net 2453 = rbit_3_0.ram_15_1.m0_s 
* net 2454 = rbit_3_0.ram_15_1.m1_s 
* net 2455 = rbit_3_0.ram_15_0.m0_s 
* net 2456 = rbit_3_0.ram_15_0.m1_s 
* net 2457 = rbit_3_0.ram_14_1.m0_s 
* net 2458 = rbit_3_0.ram_14_1.m1_s 
* net 2459 = rbit_3_0.ram_14_0.m0_s 
* net 2460 = rbit_3_0.ram_14_0.m1_s 
* net 2461 = rbit_3_0.ram_13_1.m0_s 
* net 2462 = rbit_3_0.ram_13_1.m1_s 
* net 2463 = rbit_3_0.ram_13_0.m0_s 
* net 2464 = rbit_3_0.ram_13_0.m1_s 
* net 2465 = rbit_3_0.ram_12_1.m0_s 
* net 2466 = rbit_3_0.ram_12_1.m1_s 
* net 2467 = rbit_3_0.ram_12_0.m0_s 
* net 2468 = rbit_3_0.ram_12_0.m1_s 
* net 2469 = rbit_3_0.ram_11_1.m0_s 
* net 2470 = rbit_3_0.ram_11_1.m1_s 
* net 2471 = rbit_3_0.ram_11_0.m0_s 
* net 2472 = rbit_3_0.ram_11_0.m1_s 
* net 2473 = rbit_3_0.ram_10_1.m0_s 
* net 2474 = rbit_3_0.ram_10_1.m1_s 
* net 2475 = rbit_3_0.ram_10_0.m0_s 
* net 2476 = rbit_3_0.ram_10_0.m1_s 
* net 2477 = rbit_3_0.ram_9_1.m0_s 
* net 2478 = rbit_3_0.ram_9_1.m1_s 
* net 2479 = rbit_3_0.ram_9_0.m0_s 
* net 2480 = rbit_3_0.ram_9_0.m1_s 
* net 2481 = rbit_3_0.ram_8_1.m0_s 
* net 2482 = rbit_3_0.ram_8_1.m1_s 
* net 2483 = rbit_3_0.ram_8_0.m0_s 
* net 2484 = rbit_3_0.ram_8_0.m1_s 
* net 2485 = rbit_3_0.ram_7_1.m0_s 
* net 2486 = rbit_3_0.ram_7_1.m1_s 
* net 2487 = rbit_3_0.ram_7_0.m0_s 
* net 2488 = rbit_3_0.ram_7_0.m1_s 
* net 2489 = rbit_3_0.ram_6_1.m0_s 
* net 2490 = rbit_3_0.ram_6_1.m1_s 
* net 2491 = rbit_3_0.ram_6_0.m0_s 
* net 2492 = rbit_3_0.ram_6_0.m1_s 
* net 2493 = rbit_3_0.ram_5_1.m0_s 
* net 2494 = rbit_3_0.ram_5_1.m1_s 
* net 2495 = rbit_3_0.ram_5_0.m0_s 
* net 2496 = rbit_3_0.ram_5_0.m1_s 
* net 2497 = rbit_3_0.ram_4_1.m0_s 
* net 2498 = rbit_3_0.ram_4_1.m1_s 
* net 2499 = rbit_3_0.ram_4_0.m0_s 
* net 2500 = rbit_3_0.ram_4_0.m1_s 
* net 2501 = rbit_3_0.ram_3_1.m0_s 
* net 2502 = rbit_3_0.ram_3_1.m1_s 
* net 2503 = rbit_3_0.ram_3_0.m0_s 
* net 2504 = rbit_3_0.ram_3_0.m1_s 
* net 2505 = rbit_3_0.ram_2_1.m0_s 
* net 2506 = rbit_3_0.ram_2_1.m1_s 
* net 2507 = rbit_3_0.ram_2_0.m0_s 
* net 2508 = rbit_3_0.ram_2_0.m1_s 
* net 2509 = rbit_3_0.ram_1_1.m0_s 
* net 2510 = rbit_3_0.ram_1_1.m1_s 
* net 2511 = rbit_3_0.ram_1_0.m0_s 
* net 2512 = rbit_3_0.ram_1_0.m1_s 
* net 2513 = rbit_3_0.ram_0_1.m0_s 
* net 2514 = rbit_3_0.ram_0_1.m1_s 
* net 2515 = rbit_3_0.ram_0_0.m0_s 
* net 2516 = rbit_3_0.ram_0_0.m1_s 
* net 2517 = mbk_sig138 
* net 2518 = mbk_sig114 
* net 2519 = mbk_sig164 
* net 2520 = mbk_sig115 
* net 2521 = mbk_sig183 
* net 2522 = mbk_sig22 
* net 2523 = mbk_sig18 
* net 2524 = mbk_sig69 
* net 2525 = mbk_sig101 
* net 2526 = mbk_sig93 
* net 2527 = mbk_sig85 
* net 2528 = mbk_sig5201 
* net 2529 = mbk_sig5195 
* net 2530 = mbk_sig5199 
* net 2531 = mbk_sig5198 
* net 2532 = mbk_sig5196 
* net 2533 = decod.decd_31.wld[0] 
* net 2534 = decod.decd_31.wld[2] 
* net 2535 = decod.decd_31.wld[1] 
* net 2536 = decod.decd_31.wld[3] 
* net 2537 = decod.decd_31.cd 
* net 2538 = mbk_sig5138 
* net 2539 = mbk_sig5080 
* net 2540 = mbk_sig5079 
* net 2541 = decod.decg_31.wlg[2] 
* net 2542 = mbk_sig5136 
* net 2543 = decod.decg_31.wlg[1] 
* net 2544 = mbk_sig5074 
* net 2545 = decod.decg_31.wlg[0] 
* net 2546 = mbk_sig5075 
* net 2547 = decod.decg_31.wlg[3] 
* net 2548 = mbk_sig5175 
* net 2549 = decod.decd_30.wld[0] 
* net 2550 = decod.decd_30.wld[2] 
* net 2551 = decod.decd_30.wld[1] 
* net 2552 = decod.decd_30.wld[3] 
* net 2553 = decod.decd_30.cd 
* net 2554 = mbk_sig4984 
* net 2555 = mbk_sig4944 
* net 2556 = mbk_sig4942 
* net 2557 = decod.decg_30.wlg[2] 
* net 2558 = mbk_sig4981 
* net 2559 = decod.decg_30.wlg[1] 
* net 2560 = mbk_sig4940 
* net 2561 = decod.decg_30.wlg[0] 
* net 2562 = mbk_sig4901 
* net 2563 = decod.decg_30.wlg[3] 
* net 2564 = mbk_sig4982 
* net 2565 = decod.decd_29.wld[0] 
* net 2566 = decod.decd_29.wld[2] 
* net 2567 = decod.decd_29.wld[1] 
* net 2568 = decod.decd_29.wld[3] 
* net 2569 = decod.decd_29.cd 
* net 2570 = mbk_sig4846 
* net 2571 = mbk_sig4790 
* net 2572 = mbk_sig4748 
* net 2573 = decod.decg_29.wlg[2] 
* net 2574 = mbk_sig4787 
* net 2575 = decod.decg_29.wlg[1] 
* net 2576 = mbk_sig4786 
* net 2577 = decod.decg_29.wlg[0] 
* net 2578 = mbk_sig4747 
* net 2579 = decod.decg_29.wlg[3] 
* net 2580 = mbk_sig4844 
* net 2581 = decod.decd_28.wld[0] 
* net 2582 = decod.decd_28.wld[2] 
* net 2583 = decod.decd_28.wld[1] 
* net 2584 = decod.decd_28.wld[3] 
* net 2585 = decod.decd_28.cd 
* net 2586 = mbk_sig4672 
* net 2587 = mbk_sig4614 
* net 2588 = mbk_sig4613 
* net 2589 = decod.decg_28.wlg[2] 
* net 2590 = mbk_sig4669 
* net 2591 = decod.decg_28.wlg[1] 
* net 2592 = mbk_sig4610 
* net 2593 = decod.decg_28.wlg[0] 
* net 2594 = mbk_sig4608 
* net 2595 = decod.decg_28.wlg[3] 
* net 2596 = mbk_sig4710 
* net 2597 = decod.decd_27.wld[0] 
* net 2598 = decod.decd_27.wld[2] 
* net 2599 = decod.decd_27.wld[1] 
* net 2600 = decod.decd_27.wld[3] 
* net 2601 = decod.decd_27.cd 
* net 2602 = mbk_sig4519 
* net 2603 = mbk_sig4478 
* net 2604 = mbk_sig4476 
* net 2605 = decod.decg_27.wlg[2] 
* net 2606 = mbk_sig4516 
* net 2607 = decod.decg_27.wlg[1] 
* net 2608 = mbk_sig4474 
* net 2609 = decod.decg_27.wlg[0] 
* net 2610 = mbk_sig4434 
* net 2611 = decod.decg_27.wlg[3] 
* net 2612 = mbk_sig4517 
* net 2613 = decod.decd_26.wld[0] 
* net 2614 = decod.decd_26.wld[2] 
* net 2615 = decod.decd_26.wld[1] 
* net 2616 = decod.decd_26.wld[3] 
* net 2617 = decod.decd_26.cd 
* net 2618 = mbk_sig4380 
* net 2619 = mbk_sig4325 
* net 2620 = mbk_sig4323 
* net 2621 = decod.decg_26.wlg[2] 
* net 2622 = mbk_sig4321 
* net 2623 = decod.decg_26.wlg[1] 
* net 2624 = mbk_sig4320 
* net 2625 = decod.decg_26.wlg[0] 
* net 2626 = mbk_sig4282 
* net 2627 = decod.decg_26.wlg[3] 
* net 2628 = mbk_sig4378 
* net 2629 = decod.decd_25.wld[0] 
* net 2630 = decod.decd_25.wld[2] 
* net 2631 = decod.decd_25.wld[1] 
* net 2632 = decod.decd_25.wld[3] 
* net 2633 = decod.decd_25.cd 
* net 2634 = mbk_sig4244 
* net 2635 = mbk_sig4130 
* net 2636 = mbk_sig4129 
* net 2637 = decod.decg_25.wlg[2] 
* net 2638 = mbk_sig4185 
* net 2639 = decod.decg_25.wlg[1] 
* net 2640 = mbk_sig4131 
* net 2641 = decod.decg_25.wlg[0] 
* net 2642 = mbk_sig4127 
* net 2643 = decod.decg_25.wlg[3] 
* net 2644 = mbk_sig4242 
* net 2645 = decod.decd_24.wld[0] 
* net 2646 = decod.decd_24.wld[2] 
* net 2647 = decod.decd_24.wld[1] 
* net 2648 = decod.decd_24.wld[3] 
* net 2649 = decod.decd_24.cd 
* net 2650 = mbk_sig4053 
* net 2651 = mbk_sig4012 
* net 2652 = mbk_sig4010 
* net 2653 = decod.decg_24.wlg[2] 
* net 2654 = mbk_sig4051 
* net 2655 = decod.decg_24.wlg[1] 
* net 2656 = mbk_sig4008 
* net 2657 = decod.decg_24.wlg[0] 
* net 2658 = mbk_sig3953 
* net 2659 = decod.decg_24.wlg[3] 
* net 2660 = mbk_sig4090 
* net 2661 = decod.decd_23.wld[0] 
* net 2662 = decod.decd_23.wld[2] 
* net 2663 = decod.decd_23.wld[1] 
* net 2664 = decod.decd_23.wld[3] 
* net 2665 = decod.decd_23.cd 
* net 2666 = mbk_sig3899 
* net 2667 = mbk_sig3859 
* net 2668 = mbk_sig3857 
* net 2669 = decod.decg_23.wlg[2] 
* net 2670 = mbk_sig3896 
* net 2671 = decod.decg_23.wlg[1] 
* net 2672 = mbk_sig3855 
* net 2673 = decod.decg_23.wlg[0] 
* net 2674 = mbk_sig3817 
* net 2675 = decod.decg_23.wlg[3] 
* net 2676 = mbk_sig3897 
* net 2677 = decod.decd_22.wld[0] 
* net 2678 = decod.decd_22.wld[2] 
* net 2679 = decod.decd_22.wld[1] 
* net 2680 = decod.decd_22.wld[3] 
* net 2681 = decod.decd_22.cd 
* net 2682 = mbk_sig3778 
* net 2683 = mbk_sig3664 
* net 2684 = mbk_sig3663 
* net 2685 = decod.decg_22.wlg[2] 
* net 2686 = mbk_sig3720 
* net 2687 = decod.decg_22.wlg[1] 
* net 2688 = mbk_sig3719 
* net 2689 = decod.decg_22.wlg[0] 
* net 2690 = mbk_sig3662 
* net 2691 = decod.decg_22.wlg[3] 
* net 2692 = mbk_sig3776 
* net 2693 = decod.decd_21.wld[0] 
* net 2694 = decod.decd_21.wld[2] 
* net 2695 = decod.decd_21.wld[1] 
* net 2696 = decod.decd_21.wld[3] 
* net 2697 = decod.decd_21.cd 
* net 2698 = mbk_sig3588 
* net 2699 = mbk_sig3531 
* net 2700 = mbk_sig3530 
* net 2701 = decod.decg_21.wlg[2] 
* net 2702 = mbk_sig3586 
* net 2703 = decod.decg_21.wlg[1] 
* net 2704 = mbk_sig3526 
* net 2705 = decod.decg_21.wlg[0] 
* net 2706 = mbk_sig3527 
* net 2707 = decod.decg_21.wlg[3] 
* net 2708 = mbk_sig3625 
* net 2709 = decod.decd_20.wld[0] 
* net 2710 = decod.decd_20.wld[2] 
* net 2711 = decod.decd_20.wld[1] 
* net 2712 = decod.decd_20.wld[3] 
* net 2713 = decod.decd_20.cd 
* net 2714 = mbk_sig3434 
* net 2715 = mbk_sig3394 
* net 2716 = mbk_sig3392 
* net 2717 = decod.decg_20.wlg[2] 
* net 2718 = mbk_sig3431 
* net 2719 = decod.decg_20.wlg[1] 
* net 2720 = mbk_sig3390 
* net 2721 = decod.decg_20.wlg[0] 
* net 2722 = mbk_sig3351 
* net 2723 = decod.decg_20.wlg[3] 
* net 2724 = mbk_sig3432 
* net 2725 = decod.decd_19.wld[0] 
* net 2726 = decod.decd_19.wld[2] 
* net 2727 = decod.decd_19.wld[1] 
* net 2728 = decod.decd_19.wld[3] 
* net 2729 = decod.decd_19.cd 
* net 2730 = mbk_sig3296 
* net 2731 = mbk_sig3240 
* net 2732 = mbk_sig3198 
* net 2733 = decod.decg_19.wlg[2] 
* net 2734 = mbk_sig3237 
* net 2735 = decod.decg_19.wlg[1] 
* net 2736 = mbk_sig3236 
* net 2737 = decod.decg_19.wlg[0] 
* net 2738 = mbk_sig3197 
* net 2739 = decod.decg_19.wlg[3] 
* net 2740 = mbk_sig3294 
* net 2741 = decod.decd_18.wld[0] 
* net 2742 = decod.decd_18.wld[2] 
* net 2743 = decod.decd_18.wld[1] 
* net 2744 = decod.decd_18.wld[3] 
* net 2745 = decod.decd_18.cd 
* net 2746 = mbk_sig3122 
* net 2747 = mbk_sig3064 
* net 2748 = mbk_sig3063 
* net 2749 = decod.decg_18.wlg[2] 
* net 2750 = mbk_sig3119 
* net 2751 = decod.decg_18.wlg[1] 
* net 2752 = mbk_sig3060 
* net 2753 = decod.decg_18.wlg[0] 
* net 2754 = mbk_sig3058 
* net 2755 = decod.decg_18.wlg[3] 
* net 2756 = mbk_sig3160 
* net 2757 = decod.decd_17.wld[0] 
* net 2758 = decod.decd_17.wld[2] 
* net 2759 = decod.decd_17.wld[1] 
* net 2760 = decod.decd_17.wld[3] 
* net 2761 = decod.decd_17.cd 
* net 2762 = mbk_sig2969 
* net 2763 = mbk_sig2928 
* net 2764 = mbk_sig2926 
* net 2765 = decod.decg_17.wlg[2] 
* net 2766 = mbk_sig2966 
* net 2767 = decod.decg_17.wlg[1] 
* net 2768 = mbk_sig2924 
* net 2769 = decod.decg_17.wlg[0] 
* net 2770 = mbk_sig2885 
* net 2771 = decod.decg_17.wlg[3] 
* net 2772 = mbk_sig2967 
* net 2773 = decod.decd_16.wld[0] 
* net 2774 = decod.decd_16.wld[2] 
* net 2775 = decod.decd_16.wld[1] 
* net 2776 = decod.decd_16.wld[3] 
* net 2777 = decod.decd_16.cd 
* net 2778 = mbk_sig2831 
* net 2779 = mbk_sig2775 
* net 2780 = mbk_sig2773 
* net 2781 = decod.decg_16.wlg[2] 
* net 2782 = mbk_sig2771 
* net 2783 = decod.decg_16.wlg[1] 
* net 2784 = mbk_sig2770 
* net 2785 = decod.decg_16.wlg[0] 
* net 2786 = mbk_sig2732 
* net 2787 = decod.decg_16.wlg[3] 
* net 2788 = mbk_sig2829 
* net 2789 = decod.decd_15.wld[0] 
* net 2790 = decod.decd_15.wld[2] 
* net 2791 = decod.decd_15.wld[1] 
* net 2792 = decod.decd_15.wld[3] 
* net 2793 = decod.decd_15.cd 
* net 2794 = mbk_sig2694 
* net 2795 = mbk_sig2580 
* net 2796 = mbk_sig2579 
* net 2797 = decod.decg_15.wlg[2] 
* net 2798 = mbk_sig2635 
* net 2799 = decod.decg_15.wlg[1] 
* net 2800 = mbk_sig2581 
* net 2801 = decod.decg_15.wlg[0] 
* net 2802 = mbk_sig2577 
* net 2803 = decod.decg_15.wlg[3] 
* net 2804 = mbk_sig2692 
* net 2805 = decod.decd_14.wld[0] 
* net 2806 = decod.decd_14.wld[2] 
* net 2807 = decod.decd_14.wld[1] 
* net 2808 = decod.decd_14.wld[3] 
* net 2809 = decod.decd_14.cd 
* net 2810 = mbk_sig2503 
* net 2811 = mbk_sig2462 
* net 2812 = mbk_sig2460 
* net 2813 = decod.decg_14.wlg[2] 
* net 2814 = mbk_sig2501 
* net 2815 = decod.decg_14.wlg[1] 
* net 2816 = mbk_sig2458 
* net 2817 = decod.decg_14.wlg[0] 
* net 2818 = mbk_sig2403 
* net 2819 = decod.decg_14.wlg[3] 
* net 2820 = mbk_sig2540 
* net 2821 = decod.decd_13.wld[0] 
* net 2822 = decod.decd_13.wld[2] 
* net 2823 = decod.decd_13.wld[1] 
* net 2824 = decod.decd_13.wld[3] 
* net 2825 = decod.decd_13.cd 
* net 2826 = mbk_sig2349 
* net 2827 = mbk_sig2309 
* net 2828 = mbk_sig2307 
* net 2829 = decod.decg_13.wlg[2] 
* net 2830 = mbk_sig2346 
* net 2831 = decod.decg_13.wlg[1] 
* net 2832 = mbk_sig2305 
* net 2833 = decod.decg_13.wlg[0] 
* net 2834 = mbk_sig2267 
* net 2835 = decod.decg_13.wlg[3] 
* net 2836 = mbk_sig2347 
* net 2837 = decod.decd_12.wld[0] 
* net 2838 = decod.decd_12.wld[2] 
* net 2839 = decod.decd_12.wld[1] 
* net 2840 = decod.decd_12.wld[3] 
* net 2841 = decod.decd_12.cd 
* net 2842 = mbk_sig2228 
* net 2843 = mbk_sig2114 
* net 2844 = mbk_sig2113 
* net 2845 = decod.decg_12.wlg[2] 
* net 2846 = mbk_sig2169 
* net 2847 = decod.decg_12.wlg[1] 
* net 2848 = mbk_sig2170 
* net 2849 = decod.decg_12.wlg[0] 
* net 2850 = mbk_sig2112 
* net 2851 = decod.decg_12.wlg[3] 
* net 2852 = mbk_sig2226 
* net 2853 = decod.decd_11.wld[0] 
* net 2854 = decod.decd_11.wld[2] 
* net 2855 = decod.decd_11.wld[1] 
* net 2856 = decod.decd_11.wld[3] 
* net 2857 = decod.decd_11.cd 
* net 2858 = mbk_sig2038 
* net 2859 = mbk_sig1981 
* net 2860 = mbk_sig1980 
* net 2861 = decod.decg_11.wlg[2] 
* net 2862 = mbk_sig2036 
* net 2863 = decod.decg_11.wlg[1] 
* net 2864 = mbk_sig1976 
* net 2865 = decod.decg_11.wlg[0] 
* net 2866 = mbk_sig1977 
* net 2867 = decod.decg_11.wlg[3] 
* net 2868 = mbk_sig2075 
* net 2869 = decod.decd_10.wld[0] 
* net 2870 = decod.decd_10.wld[2] 
* net 2871 = decod.decd_10.wld[1] 
* net 2872 = decod.decd_10.wld[3] 
* net 2873 = decod.decd_10.cd 
* net 2874 = mbk_sig1884 
* net 2875 = mbk_sig1844 
* net 2876 = mbk_sig1842 
* net 2877 = decod.decg_10.wlg[2] 
* net 2878 = mbk_sig1881 
* net 2879 = decod.decg_10.wlg[1] 
* net 2880 = mbk_sig1840 
* net 2881 = decod.decg_10.wlg[0] 
* net 2882 = mbk_sig1801 
* net 2883 = decod.decg_10.wlg[3] 
* net 2884 = mbk_sig1882 
* net 2885 = decod.decd_9.wld[0] 
* net 2886 = decod.decd_9.wld[2] 
* net 2887 = decod.decd_9.wld[1] 
* net 2888 = decod.decd_9.wld[3] 
* net 2889 = decod.decd_9.cd 
* net 2890 = mbk_sig1746 
* net 2891 = mbk_sig1690 
* net 2892 = mbk_sig1648 
* net 2893 = decod.decg_9.wlg[2] 
* net 2894 = mbk_sig1687 
* net 2895 = decod.decg_9.wlg[1] 
* net 2896 = mbk_sig1686 
* net 2897 = decod.decg_9.wlg[0] 
* net 2898 = mbk_sig1647 
* net 2899 = decod.decg_9.wlg[3] 
* net 2900 = mbk_sig1744 
* net 2901 = decod.decd_8.wld[0] 
* net 2902 = decod.decd_8.wld[2] 
* net 2903 = decod.decd_8.wld[1] 
* net 2904 = decod.decd_8.wld[3] 
* net 2905 = decod.decd_8.cd 
* net 2906 = mbk_sig1572 
* net 2907 = mbk_sig1514 
* net 2908 = mbk_sig1513 
* net 2909 = decod.decg_8.wlg[2] 
* net 2910 = mbk_sig1569 
* net 2911 = decod.decg_8.wlg[1] 
* net 2912 = mbk_sig1510 
* net 2913 = decod.decg_8.wlg[0] 
* net 2914 = mbk_sig1508 
* net 2915 = decod.decg_8.wlg[3] 
* net 2916 = mbk_sig1610 
* net 2917 = decod.decd_7.wld[0] 
* net 2918 = decod.decd_7.wld[2] 
* net 2919 = decod.decd_7.wld[1] 
* net 2920 = decod.decd_7.wld[3] 
* net 2921 = decod.decd_7.cd 
* net 2922 = mbk_sig1419 
* net 2923 = mbk_sig1379 
* net 2924 = mbk_sig1377 
* net 2925 = decod.decg_7.wlg[2] 
* net 2926 = mbk_sig1416 
* net 2927 = decod.decg_7.wlg[1] 
* net 2928 = mbk_sig1375 
* net 2929 = decod.decg_7.wlg[0] 
* net 2930 = mbk_sig1335 
* net 2931 = decod.decg_7.wlg[3] 
* net 2932 = mbk_sig1417 
* net 2933 = decod.decd_6.wld[0] 
* net 2934 = decod.decd_6.wld[2] 
* net 2935 = decod.decd_6.wld[1] 
* net 2936 = decod.decd_6.wld[3] 
* net 2937 = decod.decd_6.cd 
* net 2938 = mbk_sig1281 
* net 2939 = mbk_sig1225 
* net 2940 = mbk_sig1223 
* net 2941 = decod.decg_6.wlg[2] 
* net 2942 = mbk_sig1221 
* net 2943 = decod.decg_6.wlg[1] 
* net 2944 = mbk_sig1220 
* net 2945 = decod.decg_6.wlg[0] 
* net 2946 = mbk_sig1182 
* net 2947 = decod.decg_6.wlg[3] 
* net 2948 = mbk_sig1279 
* net 2949 = decod.decd_5.wld[0] 
* net 2950 = decod.decd_5.wld[2] 
* net 2951 = decod.decd_5.wld[1] 
* net 2952 = decod.decd_5.wld[3] 
* net 2953 = decod.decd_5.cd 
* net 2954 = mbk_sig1144 
* net 2955 = mbk_sig1030 
* net 2956 = mbk_sig1029 
* net 2957 = decod.decg_5.wlg[2] 
* net 2958 = mbk_sig1085 
* net 2959 = decod.decg_5.wlg[1] 
* net 2960 = mbk_sig1031 
* net 2961 = decod.decg_5.wlg[0] 
* net 2962 = mbk_sig1027 
* net 2963 = decod.decg_5.wlg[3] 
* net 2964 = mbk_sig1142 
* net 2965 = decod.decd_4.wld[0] 
* net 2966 = decod.decd_4.wld[2] 
* net 2967 = decod.decd_4.wld[1] 
* net 2968 = decod.decd_4.wld[3] 
* net 2969 = decod.decd_4.cd 
* net 2970 = mbk_sig953 
* net 2971 = mbk_sig913 
* net 2972 = mbk_sig911 
* net 2973 = decod.decg_4.wlg[2] 
* net 2974 = mbk_sig951 
* net 2975 = decod.decg_4.wlg[1] 
* net 2976 = mbk_sig909 
* net 2977 = decod.decg_4.wlg[0] 
* net 2978 = mbk_sig853 
* net 2979 = decod.decg_4.wlg[3] 
* net 2980 = mbk_sig990 
* net 2981 = decod.decd_3.wld[0] 
* net 2982 = decod.decd_3.wld[2] 
* net 2983 = decod.decd_3.wld[1] 
* net 2984 = decod.decd_3.wld[3] 
* net 2985 = decod.decd_3.cd 
* net 2986 = mbk_sig799 
* net 2987 = mbk_sig760 
* net 2988 = mbk_sig758 
* net 2989 = decod.decg_3.wlg[2] 
* net 2990 = mbk_sig756 
* net 2991 = decod.decg_3.wlg[1] 
* net 2992 = mbk_sig755 
* net 2993 = decod.decg_3.wlg[0] 
* net 2994 = mbk_sig717 
* net 2995 = decod.decg_3.wlg[3] 
* net 2996 = mbk_sig797 
* net 2997 = decod.decd_2.wld[0] 
* net 2998 = decod.decd_2.wld[2] 
* net 2999 = decod.decd_2.wld[1] 
* net 3000 = decod.decd_2.wld[3] 
* net 3001 = decod.decd_2.cd 
* net 3002 = mbk_sig678 
* net 3003 = mbk_sig565 
* net 3004 = mbk_sig564 
* net 3005 = decod.decg_2.wlg[2] 
* net 3006 = mbk_sig619 
* net 3007 = decod.decg_2.wlg[1] 
* net 3008 = mbk_sig620 
* net 3009 = decod.decg_2.wlg[0] 
* net 3010 = mbk_sig562 
* net 3011 = decod.decg_2.wlg[3] 
* net 3012 = mbk_sig676 
* net 3013 = decod.decd_1.wld[0] 
* net 3014 = decod.decd_1.wld[2] 
* net 3015 = decod.decd_1.wld[1] 
* net 3016 = decod.decd_1.wld[3] 
* net 3017 = decod.decd_1.cd 
* net 3018 = mbk_sig488 
* net 3019 = mbk_sig447 
* net 3020 = mbk_sig446 
* net 3021 = decod.decg_1.wlg[2] 
* net 3022 = mbk_sig486 
* net 3023 = decod.decg_1.wlg[1] 
* net 3024 = mbk_sig443 
* net 3025 = decod.decg_1.wlg[0] 
* net 3026 = mbk_sig388 
* net 3027 = decod.decg_1.wlg[3] 
* net 3028 = mbk_sig525 
* net 3029 = decod.decd_0.wld[0] 
* net 3030 = decod.decd_0.wld[2] 
* net 3031 = decod.decd_0.wld[1] 
* net 3032 = decod.decd_0.wld[3] 
* net 3033 = decod.decd_0.cd 
* net 3034 = mbk_sig334 
* net 3035 = mbk_sig294 
* net 3036 = mbk_sig292 
* net 3037 = decod.decg_0.wlg[2] 
* net 3038 = mbk_sig331 
* net 3039 = decod.decg_0.wlg[1] 
* net 3040 = mbk_sig290 
* net 3041 = decod.decg_0.wlg[0] 
* net 3042 = mbk_sig252 
* net 3043 = decod.decg_0.wlg[3] 
* net 3044 = mbk_sig332 
* net 3045 = mbk_sig202 
* net 3046 = mbk_sig203 
* net 3047 = mbk_sig185 
* net 3048 = mbk_sig196 
* net 3049 = mbk_sig187 
* net 3050 = mbk_sig178 
* net 3051 = decod.adr_1.adr_n[7] 
* net 3052 = mbk_sig186 
* net 3053 = mbk_sig166 
* net 3054 = mbk_sig177 
* net 3055 = mbk_sig179 
* net 3056 = mbk_sig167 
* net 3057 = mbk_sig165 
* net 3058 = mbk_sig168 
* net 3059 = mbk_sig155 
* net 3060 = mbk_sig154 
* net 3061 = mbk_sig156 
* net 3062 = mbk_sig116 
* net 3063 = mbk_sig121 
* net 3064 = decod.decd_0.cp[3] 
* net 3065 = mbk_sig142 
* net 3066 = mbk_sig143 
* net 3067 = decod.decd_0.cp[1] 
* net 3068 = decod.decd_0.cp[2] 
* net 3069 = mbk_sig117 
* net 3070 = mbk_sig119 
* net 3071 = decod.decd_0.cp[0] 
* net 3072 = mbk_sig107 
* net 3073 = mbk_sig106 
* net 3074 = mbk_sig80 
* net 3075 = mbk_sig72 
* net 3076 = mbk_sig74 
* net 3077 = mbk_sig5 
* net 3078 = mbk_sig70 
* net 3079 = mbk_sig73 
* net 3080 = mbk_sig64 
* net 3081 = mbk_sig44 
* net 3082 = mbk_sig61 
* net 3083 = mbk_sig6 
* net 3084 = mbk_sig63 
* net 3085 = decod.compg.cmk[0] 
* net 3086 = mbk_sig25 
* net 3087 = rbit_0_1.ram_127_1.m0_s 
* net 3088 = rbit_0_1.ram_127_1.m1_s 
* net 3089 = rbit_0_1.ram_127_0.m0_s 
* net 3090 = rbit_0_1.ram_127_0.m1_s 
* net 3091 = rbit_0_1.ram_126_1.m0_s 
* net 3092 = rbit_0_1.ram_126_1.m1_s 
* net 3093 = rbit_0_1.ram_126_0.m0_s 
* net 3094 = rbit_0_1.ram_126_0.m1_s 
* net 3095 = rbit_0_1.ram_125_1.m0_s 
* net 3096 = rbit_0_1.ram_125_1.m1_s 
* net 3097 = rbit_0_1.ram_125_0.m0_s 
* net 3098 = rbit_0_1.ram_125_0.m1_s 
* net 3099 = rbit_0_1.ram_124_1.m0_s 
* net 3100 = rbit_0_1.ram_124_1.m1_s 
* net 3101 = rbit_0_1.ram_124_0.m0_s 
* net 3102 = rbit_0_1.ram_124_0.m1_s 
* net 3103 = rbit_0_1.ram_123_1.m0_s 
* net 3104 = rbit_0_1.ram_123_1.m1_s 
* net 3105 = rbit_0_1.ram_123_0.m0_s 
* net 3106 = rbit_0_1.ram_123_0.m1_s 
* net 3107 = rbit_0_1.ram_122_1.m0_s 
* net 3108 = rbit_0_1.ram_122_1.m1_s 
* net 3109 = rbit_0_1.ram_122_0.m0_s 
* net 3110 = rbit_0_1.ram_122_0.m1_s 
* net 3111 = rbit_0_1.ram_121_1.m0_s 
* net 3112 = rbit_0_1.ram_121_1.m1_s 
* net 3113 = rbit_0_1.ram_121_0.m0_s 
* net 3114 = rbit_0_1.ram_121_0.m1_s 
* net 3115 = rbit_0_1.ram_120_1.m0_s 
* net 3116 = rbit_0_1.ram_120_1.m1_s 
* net 3117 = rbit_0_1.ram_120_0.m0_s 
* net 3118 = rbit_0_1.ram_120_0.m1_s 
* net 3119 = rbit_0_1.ram_119_1.m0_s 
* net 3120 = rbit_0_1.ram_119_1.m1_s 
* net 3121 = rbit_0_1.ram_119_0.m0_s 
* net 3122 = rbit_0_1.ram_119_0.m1_s 
* net 3123 = rbit_0_1.ram_118_1.m0_s 
* net 3124 = rbit_0_1.ram_118_1.m1_s 
* net 3125 = rbit_0_1.ram_118_0.m0_s 
* net 3126 = rbit_0_1.ram_118_0.m1_s 
* net 3127 = rbit_0_1.ram_117_1.m0_s 
* net 3128 = rbit_0_1.ram_117_1.m1_s 
* net 3129 = rbit_0_1.ram_117_0.m0_s 
* net 3130 = rbit_0_1.ram_117_0.m1_s 
* net 3131 = rbit_0_1.ram_116_1.m0_s 
* net 3132 = rbit_0_1.ram_116_1.m1_s 
* net 3133 = rbit_0_1.ram_116_0.m0_s 
* net 3134 = rbit_0_1.ram_116_0.m1_s 
* net 3135 = rbit_0_1.ram_115_1.m0_s 
* net 3136 = rbit_0_1.ram_115_1.m1_s 
* net 3137 = rbit_0_1.ram_115_0.m0_s 
* net 3138 = rbit_0_1.ram_115_0.m1_s 
* net 3139 = rbit_0_1.ram_114_1.m0_s 
* net 3140 = rbit_0_1.ram_114_1.m1_s 
* net 3141 = rbit_0_1.ram_114_0.m0_s 
* net 3142 = rbit_0_1.ram_114_0.m1_s 
* net 3143 = rbit_0_1.ram_113_1.m0_s 
* net 3144 = rbit_0_1.ram_113_1.m1_s 
* net 3145 = rbit_0_1.ram_113_0.m0_s 
* net 3146 = rbit_0_1.ram_113_0.m1_s 
* net 3147 = rbit_0_1.ram_112_1.m0_s 
* net 3148 = rbit_0_1.ram_112_1.m1_s 
* net 3149 = rbit_0_1.ram_112_0.m0_s 
* net 3150 = rbit_0_1.ram_112_0.m1_s 
* net 3151 = rbit_0_1.ram_111_1.m0_s 
* net 3152 = rbit_0_1.ram_111_1.m1_s 
* net 3153 = rbit_0_1.ram_111_0.m0_s 
* net 3154 = rbit_0_1.ram_111_0.m1_s 
* net 3155 = rbit_0_1.ram_110_1.m0_s 
* net 3156 = rbit_0_1.ram_110_1.m1_s 
* net 3157 = rbit_0_1.ram_110_0.m0_s 
* net 3158 = rbit_0_1.ram_110_0.m1_s 
* net 3159 = rbit_0_1.ram_109_1.m0_s 
* net 3160 = rbit_0_1.ram_109_1.m1_s 
* net 3161 = rbit_0_1.ram_109_0.m0_s 
* net 3162 = rbit_0_1.ram_109_0.m1_s 
* net 3163 = rbit_0_1.ram_108_1.m0_s 
* net 3164 = rbit_0_1.ram_108_1.m1_s 
* net 3165 = rbit_0_1.ram_108_0.m0_s 
* net 3166 = rbit_0_1.ram_108_0.m1_s 
* net 3167 = rbit_0_1.ram_107_1.m0_s 
* net 3168 = rbit_0_1.ram_107_1.m1_s 
* net 3169 = rbit_0_1.ram_107_0.m0_s 
* net 3170 = rbit_0_1.ram_107_0.m1_s 
* net 3171 = rbit_0_1.ram_106_1.m0_s 
* net 3172 = rbit_0_1.ram_106_1.m1_s 
* net 3173 = rbit_0_1.ram_106_0.m0_s 
* net 3174 = rbit_0_1.ram_106_0.m1_s 
* net 3175 = rbit_0_1.ram_105_1.m0_s 
* net 3176 = rbit_0_1.ram_105_1.m1_s 
* net 3177 = rbit_0_1.ram_105_0.m0_s 
* net 3178 = rbit_0_1.ram_105_0.m1_s 
* net 3179 = rbit_0_1.ram_104_1.m0_s 
* net 3180 = rbit_0_1.ram_104_1.m1_s 
* net 3181 = rbit_0_1.ram_104_0.m0_s 
* net 3182 = rbit_0_1.ram_104_0.m1_s 
* net 3183 = rbit_0_1.ram_103_1.m0_s 
* net 3184 = rbit_0_1.ram_103_1.m1_s 
* net 3185 = rbit_0_1.ram_103_0.m0_s 
* net 3186 = rbit_0_1.ram_103_0.m1_s 
* net 3187 = rbit_0_1.ram_102_1.m0_s 
* net 3188 = rbit_0_1.ram_102_1.m1_s 
* net 3189 = rbit_0_1.ram_102_0.m0_s 
* net 3190 = rbit_0_1.ram_102_0.m1_s 
* net 3191 = rbit_0_1.ram_101_1.m0_s 
* net 3192 = rbit_0_1.ram_101_1.m1_s 
* net 3193 = rbit_0_1.ram_101_0.m0_s 
* net 3194 = rbit_0_1.ram_101_0.m1_s 
* net 3195 = rbit_0_1.ram_100_1.m0_s 
* net 3196 = rbit_0_1.ram_100_1.m1_s 
* net 3197 = rbit_0_1.ram_100_0.m0_s 
* net 3198 = rbit_0_1.ram_100_0.m1_s 
* net 3199 = rbit_0_1.ram_99_1.m0_s 
* net 3200 = rbit_0_1.ram_99_1.m1_s 
* net 3201 = rbit_0_1.ram_99_0.m0_s 
* net 3202 = rbit_0_1.ram_99_0.m1_s 
* net 3203 = rbit_0_1.ram_98_1.m0_s 
* net 3204 = rbit_0_1.ram_98_1.m1_s 
* net 3205 = rbit_0_1.ram_98_0.m0_s 
* net 3206 = rbit_0_1.ram_98_0.m1_s 
* net 3207 = rbit_0_1.ram_97_1.m0_s 
* net 3208 = rbit_0_1.ram_97_1.m1_s 
* net 3209 = rbit_0_1.ram_97_0.m0_s 
* net 3210 = rbit_0_1.ram_97_0.m1_s 
* net 3211 = rbit_0_1.ram_96_1.m0_s 
* net 3212 = rbit_0_1.ram_96_1.m1_s 
* net 3213 = rbit_0_1.ram_96_0.m0_s 
* net 3214 = rbit_0_1.ram_96_0.m1_s 
* net 3215 = rbit_0_1.ram_95_1.m0_s 
* net 3216 = rbit_0_1.ram_95_1.m1_s 
* net 3217 = rbit_0_1.ram_95_0.m0_s 
* net 3218 = rbit_0_1.ram_95_0.m1_s 
* net 3219 = rbit_0_1.ram_94_1.m0_s 
* net 3220 = rbit_0_1.ram_94_1.m1_s 
* net 3221 = rbit_0_1.ram_94_0.m0_s 
* net 3222 = rbit_0_1.ram_94_0.m1_s 
* net 3223 = rbit_0_1.ram_93_1.m0_s 
* net 3224 = rbit_0_1.ram_93_1.m1_s 
* net 3225 = rbit_0_1.ram_93_0.m0_s 
* net 3226 = rbit_0_1.ram_93_0.m1_s 
* net 3227 = rbit_0_1.ram_92_1.m0_s 
* net 3228 = rbit_0_1.ram_92_1.m1_s 
* net 3229 = rbit_0_1.ram_92_0.m0_s 
* net 3230 = rbit_0_1.ram_92_0.m1_s 
* net 3231 = rbit_0_1.ram_91_1.m0_s 
* net 3232 = rbit_0_1.ram_91_1.m1_s 
* net 3233 = rbit_0_1.ram_91_0.m0_s 
* net 3234 = rbit_0_1.ram_91_0.m1_s 
* net 3235 = rbit_0_1.ram_90_1.m0_s 
* net 3236 = rbit_0_1.ram_90_1.m1_s 
* net 3237 = rbit_0_1.ram_90_0.m0_s 
* net 3238 = rbit_0_1.ram_90_0.m1_s 
* net 3239 = rbit_0_1.ram_89_1.m0_s 
* net 3240 = rbit_0_1.ram_89_1.m1_s 
* net 3241 = rbit_0_1.ram_89_0.m0_s 
* net 3242 = rbit_0_1.ram_89_0.m1_s 
* net 3243 = rbit_0_1.ram_88_1.m0_s 
* net 3244 = rbit_0_1.ram_88_1.m1_s 
* net 3245 = rbit_0_1.ram_88_0.m0_s 
* net 3246 = rbit_0_1.ram_88_0.m1_s 
* net 3247 = rbit_0_1.ram_87_1.m0_s 
* net 3248 = rbit_0_1.ram_87_1.m1_s 
* net 3249 = rbit_0_1.ram_87_0.m0_s 
* net 3250 = rbit_0_1.ram_87_0.m1_s 
* net 3251 = rbit_0_1.ram_86_1.m0_s 
* net 3252 = rbit_0_1.ram_86_1.m1_s 
* net 3253 = rbit_0_1.ram_86_0.m0_s 
* net 3254 = rbit_0_1.ram_86_0.m1_s 
* net 3255 = rbit_0_1.ram_85_1.m0_s 
* net 3256 = rbit_0_1.ram_85_1.m1_s 
* net 3257 = rbit_0_1.ram_85_0.m0_s 
* net 3258 = rbit_0_1.ram_85_0.m1_s 
* net 3259 = rbit_0_1.ram_84_1.m0_s 
* net 3260 = rbit_0_1.ram_84_1.m1_s 
* net 3261 = rbit_0_1.ram_84_0.m0_s 
* net 3262 = rbit_0_1.ram_84_0.m1_s 
* net 3263 = rbit_0_1.ram_83_1.m0_s 
* net 3264 = rbit_0_1.ram_83_1.m1_s 
* net 3265 = rbit_0_1.ram_83_0.m0_s 
* net 3266 = rbit_0_1.ram_83_0.m1_s 
* net 3267 = rbit_0_1.ram_82_1.m0_s 
* net 3268 = rbit_0_1.ram_82_1.m1_s 
* net 3269 = rbit_0_1.ram_82_0.m0_s 
* net 3270 = rbit_0_1.ram_82_0.m1_s 
* net 3271 = rbit_0_1.ram_81_1.m0_s 
* net 3272 = rbit_0_1.ram_81_1.m1_s 
* net 3273 = rbit_0_1.ram_81_0.m0_s 
* net 3274 = rbit_0_1.ram_81_0.m1_s 
* net 3275 = rbit_0_1.ram_80_1.m0_s 
* net 3276 = rbit_0_1.ram_80_1.m1_s 
* net 3277 = rbit_0_1.ram_80_0.m0_s 
* net 3278 = rbit_0_1.ram_80_0.m1_s 
* net 3279 = rbit_0_1.ram_79_1.m0_s 
* net 3280 = rbit_0_1.ram_79_1.m1_s 
* net 3281 = rbit_0_1.ram_79_0.m0_s 
* net 3282 = rbit_0_1.ram_79_0.m1_s 
* net 3283 = rbit_0_1.ram_78_1.m0_s 
* net 3284 = rbit_0_1.ram_78_1.m1_s 
* net 3285 = rbit_0_1.ram_78_0.m0_s 
* net 3286 = rbit_0_1.ram_78_0.m1_s 
* net 3287 = rbit_0_1.ram_77_1.m0_s 
* net 3288 = rbit_0_1.ram_77_1.m1_s 
* net 3289 = rbit_0_1.ram_77_0.m0_s 
* net 3290 = rbit_0_1.ram_77_0.m1_s 
* net 3291 = rbit_0_1.ram_76_1.m0_s 
* net 3292 = rbit_0_1.ram_76_1.m1_s 
* net 3293 = rbit_0_1.ram_76_0.m0_s 
* net 3294 = rbit_0_1.ram_76_0.m1_s 
* net 3295 = rbit_0_1.ram_75_1.m0_s 
* net 3296 = rbit_0_1.ram_75_1.m1_s 
* net 3297 = rbit_0_1.ram_75_0.m0_s 
* net 3298 = rbit_0_1.ram_75_0.m1_s 
* net 3299 = rbit_0_1.ram_74_1.m0_s 
* net 3300 = rbit_0_1.ram_74_1.m1_s 
* net 3301 = rbit_0_1.ram_74_0.m0_s 
* net 3302 = rbit_0_1.ram_74_0.m1_s 
* net 3303 = rbit_0_1.ram_73_1.m0_s 
* net 3304 = rbit_0_1.ram_73_1.m1_s 
* net 3305 = rbit_0_1.ram_73_0.m0_s 
* net 3306 = rbit_0_1.ram_73_0.m1_s 
* net 3307 = rbit_0_1.ram_72_1.m0_s 
* net 3308 = rbit_0_1.ram_72_1.m1_s 
* net 3309 = rbit_0_1.ram_72_0.m0_s 
* net 3310 = rbit_0_1.ram_72_0.m1_s 
* net 3311 = rbit_0_1.ram_71_1.m0_s 
* net 3312 = rbit_0_1.ram_71_1.m1_s 
* net 3313 = rbit_0_1.ram_71_0.m0_s 
* net 3314 = rbit_0_1.ram_71_0.m1_s 
* net 3315 = rbit_0_1.ram_70_1.m0_s 
* net 3316 = rbit_0_1.ram_70_1.m1_s 
* net 3317 = rbit_0_1.ram_70_0.m0_s 
* net 3318 = rbit_0_1.ram_70_0.m1_s 
* net 3319 = rbit_0_1.ram_69_1.m0_s 
* net 3320 = rbit_0_1.ram_69_1.m1_s 
* net 3321 = rbit_0_1.ram_69_0.m0_s 
* net 3322 = rbit_0_1.ram_69_0.m1_s 
* net 3323 = rbit_0_1.ram_68_1.m0_s 
* net 3324 = rbit_0_1.ram_68_1.m1_s 
* net 3325 = rbit_0_1.ram_68_0.m0_s 
* net 3326 = rbit_0_1.ram_68_0.m1_s 
* net 3327 = rbit_0_1.ram_67_1.m0_s 
* net 3328 = rbit_0_1.ram_67_1.m1_s 
* net 3329 = rbit_0_1.ram_67_0.m0_s 
* net 3330 = rbit_0_1.ram_67_0.m1_s 
* net 3331 = rbit_0_1.ram_66_1.m0_s 
* net 3332 = rbit_0_1.ram_66_1.m1_s 
* net 3333 = rbit_0_1.ram_66_0.m0_s 
* net 3334 = rbit_0_1.ram_66_0.m1_s 
* net 3335 = rbit_0_1.ram_65_1.m0_s 
* net 3336 = rbit_0_1.ram_65_1.m1_s 
* net 3337 = rbit_0_1.ram_65_0.m0_s 
* net 3338 = rbit_0_1.ram_65_0.m1_s 
* net 3339 = rbit_0_1.ram_64_1.m0_s 
* net 3340 = rbit_0_1.ram_64_1.m1_s 
* net 3341 = rbit_0_1.ram_64_0.m0_s 
* net 3342 = rbit_0_1.ram_64_0.m1_s 
* net 3343 = rbit_0_1.ram_63_1.m0_s 
* net 3344 = rbit_0_1.ram_63_1.m1_s 
* net 3345 = rbit_0_1.ram_63_0.m0_s 
* net 3346 = rbit_0_1.ram_63_0.m1_s 
* net 3347 = rbit_0_1.ram_62_1.m0_s 
* net 3348 = rbit_0_1.ram_62_1.m1_s 
* net 3349 = rbit_0_1.ram_62_0.m0_s 
* net 3350 = rbit_0_1.ram_62_0.m1_s 
* net 3351 = rbit_0_1.ram_61_1.m0_s 
* net 3352 = rbit_0_1.ram_61_1.m1_s 
* net 3353 = rbit_0_1.ram_61_0.m0_s 
* net 3354 = rbit_0_1.ram_61_0.m1_s 
* net 3355 = rbit_0_1.ram_60_1.m0_s 
* net 3356 = rbit_0_1.ram_60_1.m1_s 
* net 3357 = rbit_0_1.ram_60_0.m0_s 
* net 3358 = rbit_0_1.ram_60_0.m1_s 
* net 3359 = rbit_0_1.ram_59_1.m0_s 
* net 3360 = rbit_0_1.ram_59_1.m1_s 
* net 3361 = rbit_0_1.ram_59_0.m0_s 
* net 3362 = rbit_0_1.ram_59_0.m1_s 
* net 3363 = rbit_0_1.ram_58_1.m0_s 
* net 3364 = rbit_0_1.ram_58_1.m1_s 
* net 3365 = rbit_0_1.ram_58_0.m0_s 
* net 3366 = rbit_0_1.ram_58_0.m1_s 
* net 3367 = rbit_0_1.ram_57_1.m0_s 
* net 3368 = rbit_0_1.ram_57_1.m1_s 
* net 3369 = rbit_0_1.ram_57_0.m0_s 
* net 3370 = rbit_0_1.ram_57_0.m1_s 
* net 3371 = rbit_0_1.ram_56_1.m0_s 
* net 3372 = rbit_0_1.ram_56_1.m1_s 
* net 3373 = rbit_0_1.ram_56_0.m0_s 
* net 3374 = rbit_0_1.ram_56_0.m1_s 
* net 3375 = rbit_0_1.ram_55_1.m0_s 
* net 3376 = rbit_0_1.ram_55_1.m1_s 
* net 3377 = rbit_0_1.ram_55_0.m0_s 
* net 3378 = rbit_0_1.ram_55_0.m1_s 
* net 3379 = rbit_0_1.ram_54_1.m0_s 
* net 3380 = rbit_0_1.ram_54_1.m1_s 
* net 3381 = rbit_0_1.ram_54_0.m0_s 
* net 3382 = rbit_0_1.ram_54_0.m1_s 
* net 3383 = rbit_0_1.ram_53_1.m0_s 
* net 3384 = rbit_0_1.ram_53_1.m1_s 
* net 3385 = rbit_0_1.ram_53_0.m0_s 
* net 3386 = rbit_0_1.ram_53_0.m1_s 
* net 3387 = rbit_0_1.ram_52_1.m0_s 
* net 3388 = rbit_0_1.ram_52_1.m1_s 
* net 3389 = rbit_0_1.ram_52_0.m0_s 
* net 3390 = rbit_0_1.ram_52_0.m1_s 
* net 3391 = rbit_0_1.ram_51_1.m0_s 
* net 3392 = rbit_0_1.ram_51_1.m1_s 
* net 3393 = rbit_0_1.ram_51_0.m0_s 
* net 3394 = rbit_0_1.ram_51_0.m1_s 
* net 3395 = rbit_0_1.ram_50_1.m0_s 
* net 3396 = rbit_0_1.ram_50_1.m1_s 
* net 3397 = rbit_0_1.ram_50_0.m0_s 
* net 3398 = rbit_0_1.ram_50_0.m1_s 
* net 3399 = rbit_0_1.ram_49_1.m0_s 
* net 3400 = rbit_0_1.ram_49_1.m1_s 
* net 3401 = rbit_0_1.ram_49_0.m0_s 
* net 3402 = rbit_0_1.ram_49_0.m1_s 
* net 3403 = rbit_0_1.ram_48_1.m0_s 
* net 3404 = rbit_0_1.ram_48_1.m1_s 
* net 3405 = rbit_0_1.ram_48_0.m0_s 
* net 3406 = rbit_0_1.ram_48_0.m1_s 
* net 3407 = rbit_0_1.ram_47_1.m0_s 
* net 3408 = rbit_0_1.ram_47_1.m1_s 
* net 3409 = rbit_0_1.ram_47_0.m0_s 
* net 3410 = rbit_0_1.ram_47_0.m1_s 
* net 3411 = rbit_0_1.ram_46_1.m0_s 
* net 3412 = rbit_0_1.ram_46_1.m1_s 
* net 3413 = rbit_0_1.ram_46_0.m0_s 
* net 3414 = rbit_0_1.ram_46_0.m1_s 
* net 3415 = rbit_0_1.ram_45_1.m0_s 
* net 3416 = rbit_0_1.ram_45_1.m1_s 
* net 3417 = rbit_0_1.ram_45_0.m0_s 
* net 3418 = rbit_0_1.ram_45_0.m1_s 
* net 3419 = rbit_0_1.ram_44_1.m0_s 
* net 3420 = rbit_0_1.ram_44_1.m1_s 
* net 3421 = rbit_0_1.ram_44_0.m0_s 
* net 3422 = rbit_0_1.ram_44_0.m1_s 
* net 3423 = rbit_0_1.ram_43_1.m0_s 
* net 3424 = rbit_0_1.ram_43_1.m1_s 
* net 3425 = rbit_0_1.ram_43_0.m0_s 
* net 3426 = rbit_0_1.ram_43_0.m1_s 
* net 3427 = rbit_0_1.ram_42_1.m0_s 
* net 3428 = rbit_0_1.ram_42_1.m1_s 
* net 3429 = rbit_0_1.ram_42_0.m0_s 
* net 3430 = rbit_0_1.ram_42_0.m1_s 
* net 3431 = rbit_0_1.ram_41_1.m0_s 
* net 3432 = rbit_0_1.ram_41_1.m1_s 
* net 3433 = rbit_0_1.ram_41_0.m0_s 
* net 3434 = rbit_0_1.ram_41_0.m1_s 
* net 3435 = rbit_0_1.ram_40_1.m0_s 
* net 3436 = rbit_0_1.ram_40_1.m1_s 
* net 3437 = rbit_0_1.ram_40_0.m0_s 
* net 3438 = rbit_0_1.ram_40_0.m1_s 
* net 3439 = rbit_0_1.ram_39_1.m0_s 
* net 3440 = rbit_0_1.ram_39_1.m1_s 
* net 3441 = rbit_0_1.ram_39_0.m0_s 
* net 3442 = rbit_0_1.ram_39_0.m1_s 
* net 3443 = rbit_0_1.ram_38_1.m0_s 
* net 3444 = rbit_0_1.ram_38_1.m1_s 
* net 3445 = rbit_0_1.ram_38_0.m0_s 
* net 3446 = rbit_0_1.ram_38_0.m1_s 
* net 3447 = rbit_0_1.ram_37_1.m0_s 
* net 3448 = rbit_0_1.ram_37_1.m1_s 
* net 3449 = rbit_0_1.ram_37_0.m0_s 
* net 3450 = rbit_0_1.ram_37_0.m1_s 
* net 3451 = rbit_0_1.ram_36_1.m0_s 
* net 3452 = rbit_0_1.ram_36_1.m1_s 
* net 3453 = rbit_0_1.ram_36_0.m0_s 
* net 3454 = rbit_0_1.ram_36_0.m1_s 
* net 3455 = rbit_0_1.ram_35_1.m0_s 
* net 3456 = rbit_0_1.ram_35_1.m1_s 
* net 3457 = rbit_0_1.ram_35_0.m0_s 
* net 3458 = rbit_0_1.ram_35_0.m1_s 
* net 3459 = rbit_0_1.ram_34_1.m0_s 
* net 3460 = rbit_0_1.ram_34_1.m1_s 
* net 3461 = rbit_0_1.ram_34_0.m0_s 
* net 3462 = rbit_0_1.ram_34_0.m1_s 
* net 3463 = rbit_0_1.ram_33_1.m0_s 
* net 3464 = rbit_0_1.ram_33_1.m1_s 
* net 3465 = rbit_0_1.ram_33_0.m0_s 
* net 3466 = rbit_0_1.ram_33_0.m1_s 
* net 3467 = rbit_0_1.ram_32_1.m0_s 
* net 3468 = rbit_0_1.ram_32_1.m1_s 
* net 3469 = rbit_0_1.ram_32_0.m0_s 
* net 3470 = rbit_0_1.ram_32_0.m1_s 
* net 3471 = rbit_0_1.ram_31_1.m0_s 
* net 3472 = rbit_0_1.ram_31_1.m1_s 
* net 3473 = rbit_0_1.ram_31_0.m0_s 
* net 3474 = rbit_0_1.ram_31_0.m1_s 
* net 3475 = rbit_0_1.ram_30_1.m0_s 
* net 3476 = rbit_0_1.ram_30_1.m1_s 
* net 3477 = rbit_0_1.ram_30_0.m0_s 
* net 3478 = rbit_0_1.ram_30_0.m1_s 
* net 3479 = rbit_0_1.ram_29_1.m0_s 
* net 3480 = rbit_0_1.ram_29_1.m1_s 
* net 3481 = rbit_0_1.ram_29_0.m0_s 
* net 3482 = rbit_0_1.ram_29_0.m1_s 
* net 3483 = rbit_0_1.ram_28_1.m0_s 
* net 3484 = rbit_0_1.ram_28_1.m1_s 
* net 3485 = rbit_0_1.ram_28_0.m0_s 
* net 3486 = rbit_0_1.ram_28_0.m1_s 
* net 3487 = rbit_0_1.ram_27_1.m0_s 
* net 3488 = rbit_0_1.ram_27_1.m1_s 
* net 3489 = rbit_0_1.ram_27_0.m0_s 
* net 3490 = rbit_0_1.ram_27_0.m1_s 
* net 3491 = rbit_0_1.ram_26_1.m0_s 
* net 3492 = rbit_0_1.ram_26_1.m1_s 
* net 3493 = rbit_0_1.ram_26_0.m0_s 
* net 3494 = rbit_0_1.ram_26_0.m1_s 
* net 3495 = rbit_0_1.ram_25_1.m0_s 
* net 3496 = rbit_0_1.ram_25_1.m1_s 
* net 3497 = rbit_0_1.ram_25_0.m0_s 
* net 3498 = rbit_0_1.ram_25_0.m1_s 
* net 3499 = rbit_0_1.ram_24_1.m0_s 
* net 3500 = rbit_0_1.ram_24_1.m1_s 
* net 3501 = rbit_0_1.ram_24_0.m0_s 
* net 3502 = rbit_0_1.ram_24_0.m1_s 
* net 3503 = rbit_0_1.ram_23_1.m0_s 
* net 3504 = rbit_0_1.ram_23_1.m1_s 
* net 3505 = rbit_0_1.ram_23_0.m0_s 
* net 3506 = rbit_0_1.ram_23_0.m1_s 
* net 3507 = rbit_0_1.ram_22_1.m0_s 
* net 3508 = rbit_0_1.ram_22_1.m1_s 
* net 3509 = rbit_0_1.ram_22_0.m0_s 
* net 3510 = rbit_0_1.ram_22_0.m1_s 
* net 3511 = rbit_0_1.ram_21_1.m0_s 
* net 3512 = rbit_0_1.ram_21_1.m1_s 
* net 3513 = rbit_0_1.ram_21_0.m0_s 
* net 3514 = rbit_0_1.ram_21_0.m1_s 
* net 3515 = rbit_0_1.ram_20_1.m0_s 
* net 3516 = rbit_0_1.ram_20_1.m1_s 
* net 3517 = rbit_0_1.ram_20_0.m0_s 
* net 3518 = rbit_0_1.ram_20_0.m1_s 
* net 3519 = rbit_0_1.ram_19_1.m0_s 
* net 3520 = rbit_0_1.ram_19_1.m1_s 
* net 3521 = rbit_0_1.ram_19_0.m0_s 
* net 3522 = rbit_0_1.ram_19_0.m1_s 
* net 3523 = rbit_0_1.ram_18_1.m0_s 
* net 3524 = rbit_0_1.ram_18_1.m1_s 
* net 3525 = rbit_0_1.ram_18_0.m0_s 
* net 3526 = rbit_0_1.ram_18_0.m1_s 
* net 3527 = rbit_0_1.ram_17_1.m0_s 
* net 3528 = rbit_0_1.ram_17_1.m1_s 
* net 3529 = rbit_0_1.ram_17_0.m0_s 
* net 3530 = rbit_0_1.ram_17_0.m1_s 
* net 3531 = rbit_0_1.ram_16_1.m0_s 
* net 3532 = rbit_0_1.ram_16_1.m1_s 
* net 3533 = rbit_0_1.ram_16_0.m0_s 
* net 3534 = rbit_0_1.ram_16_0.m1_s 
* net 3535 = rbit_0_1.ram_15_1.m0_s 
* net 3536 = rbit_0_1.ram_15_1.m1_s 
* net 3537 = rbit_0_1.ram_15_0.m0_s 
* net 3538 = rbit_0_1.ram_15_0.m1_s 
* net 3539 = rbit_0_1.ram_14_1.m0_s 
* net 3540 = rbit_0_1.ram_14_1.m1_s 
* net 3541 = rbit_0_1.ram_14_0.m0_s 
* net 3542 = rbit_0_1.ram_14_0.m1_s 
* net 3543 = rbit_0_1.ram_13_1.m0_s 
* net 3544 = rbit_0_1.ram_13_1.m1_s 
* net 3545 = rbit_0_1.ram_13_0.m0_s 
* net 3546 = rbit_0_1.ram_13_0.m1_s 
* net 3547 = rbit_0_1.ram_12_1.m0_s 
* net 3548 = rbit_0_1.ram_12_1.m1_s 
* net 3549 = rbit_0_1.ram_12_0.m0_s 
* net 3550 = rbit_0_1.ram_12_0.m1_s 
* net 3551 = rbit_0_1.ram_11_1.m0_s 
* net 3552 = rbit_0_1.ram_11_1.m1_s 
* net 3553 = rbit_0_1.ram_11_0.m0_s 
* net 3554 = rbit_0_1.ram_11_0.m1_s 
* net 3555 = rbit_0_1.ram_10_1.m0_s 
* net 3556 = rbit_0_1.ram_10_1.m1_s 
* net 3557 = rbit_0_1.ram_10_0.m0_s 
* net 3558 = rbit_0_1.ram_10_0.m1_s 
* net 3559 = rbit_0_1.ram_9_1.m0_s 
* net 3560 = rbit_0_1.ram_9_1.m1_s 
* net 3561 = rbit_0_1.ram_9_0.m0_s 
* net 3562 = rbit_0_1.ram_9_0.m1_s 
* net 3563 = rbit_0_1.ram_8_1.m0_s 
* net 3564 = rbit_0_1.ram_8_1.m1_s 
* net 3565 = rbit_0_1.ram_8_0.m0_s 
* net 3566 = rbit_0_1.ram_8_0.m1_s 
* net 3567 = rbit_0_1.ram_7_1.m0_s 
* net 3568 = rbit_0_1.ram_7_1.m1_s 
* net 3569 = rbit_0_1.ram_7_0.m0_s 
* net 3570 = rbit_0_1.ram_7_0.m1_s 
* net 3571 = rbit_0_1.ram_6_1.m0_s 
* net 3572 = rbit_0_1.ram_6_1.m1_s 
* net 3573 = rbit_0_1.ram_6_0.m0_s 
* net 3574 = rbit_0_1.ram_6_0.m1_s 
* net 3575 = rbit_0_1.ram_5_1.m0_s 
* net 3576 = rbit_0_1.ram_5_1.m1_s 
* net 3577 = rbit_0_1.ram_5_0.m0_s 
* net 3578 = rbit_0_1.ram_5_0.m1_s 
* net 3579 = rbit_0_1.ram_4_1.m0_s 
* net 3580 = rbit_0_1.ram_4_1.m1_s 
* net 3581 = rbit_0_1.ram_4_0.m0_s 
* net 3582 = rbit_0_1.ram_4_0.m1_s 
* net 3583 = rbit_0_1.ram_3_1.m0_s 
* net 3584 = rbit_0_1.ram_3_1.m1_s 
* net 3585 = rbit_0_1.ram_3_0.m0_s 
* net 3586 = rbit_0_1.ram_3_0.m1_s 
* net 3587 = rbit_0_1.ram_2_1.m0_s 
* net 3588 = rbit_0_1.ram_2_1.m1_s 
* net 3589 = rbit_0_1.ram_2_0.m0_s 
* net 3590 = rbit_0_1.ram_2_0.m1_s 
* net 3591 = rbit_0_1.ram_1_1.m0_s 
* net 3592 = rbit_0_1.ram_1_1.m1_s 
* net 3593 = rbit_0_1.ram_1_0.m0_s 
* net 3594 = rbit_0_1.ram_1_0.m1_s 
* net 3595 = rbit_0_1.ram_0_1.m0_s 
* net 3596 = rbit_0_1.ram_0_1.m1_s 
* net 3597 = rbit_0_1.ram_0_0.m0_s 
* net 3598 = rbit_0_1.ram_0_0.m1_s 
* net 3599 = mbk_sig147 
* net 3600 = mbk_sig125 
* net 3601 = mbk_sig169 
* net 3602 = mbk_sig124 
* net 3603 = mbk_sig188 
* net 3604 = mbk_sig40 
* net 3605 = mbk_sig43 
* net 3606 = mbk_sig76 
* net 3607 = mbk_sig102 
* net 3608 = mbk_sig94 
* net 3609 = mbk_sig86 
* net 3610 = rbit_1_1.ram_127_1.m0_s 
* net 3611 = rbit_1_1.ram_127_1.m1_s 
* net 3612 = rbit_1_1.ram_127_0.m0_s 
* net 3613 = rbit_1_1.ram_127_0.m1_s 
* net 3614 = rbit_1_1.ram_126_1.m0_s 
* net 3615 = rbit_1_1.ram_126_1.m1_s 
* net 3616 = rbit_1_1.ram_126_0.m0_s 
* net 3617 = rbit_1_1.ram_126_0.m1_s 
* net 3618 = rbit_1_1.ram_125_1.m0_s 
* net 3619 = rbit_1_1.ram_125_1.m1_s 
* net 3620 = rbit_1_1.ram_125_0.m0_s 
* net 3621 = rbit_1_1.ram_125_0.m1_s 
* net 3622 = rbit_1_1.ram_124_1.m0_s 
* net 3623 = rbit_1_1.ram_124_1.m1_s 
* net 3624 = rbit_1_1.ram_124_0.m0_s 
* net 3625 = rbit_1_1.ram_124_0.m1_s 
* net 3626 = rbit_1_1.ram_123_1.m0_s 
* net 3627 = rbit_1_1.ram_123_1.m1_s 
* net 3628 = rbit_1_1.ram_123_0.m0_s 
* net 3629 = rbit_1_1.ram_123_0.m1_s 
* net 3630 = rbit_1_1.ram_122_1.m0_s 
* net 3631 = rbit_1_1.ram_122_1.m1_s 
* net 3632 = rbit_1_1.ram_122_0.m0_s 
* net 3633 = rbit_1_1.ram_122_0.m1_s 
* net 3634 = rbit_1_1.ram_121_1.m0_s 
* net 3635 = rbit_1_1.ram_121_1.m1_s 
* net 3636 = rbit_1_1.ram_121_0.m0_s 
* net 3637 = rbit_1_1.ram_121_0.m1_s 
* net 3638 = rbit_1_1.ram_120_1.m0_s 
* net 3639 = rbit_1_1.ram_120_1.m1_s 
* net 3640 = rbit_1_1.ram_120_0.m0_s 
* net 3641 = rbit_1_1.ram_120_0.m1_s 
* net 3642 = rbit_1_1.ram_119_1.m0_s 
* net 3643 = rbit_1_1.ram_119_1.m1_s 
* net 3644 = rbit_1_1.ram_119_0.m0_s 
* net 3645 = rbit_1_1.ram_119_0.m1_s 
* net 3646 = rbit_1_1.ram_118_1.m0_s 
* net 3647 = rbit_1_1.ram_118_1.m1_s 
* net 3648 = rbit_1_1.ram_118_0.m0_s 
* net 3649 = rbit_1_1.ram_118_0.m1_s 
* net 3650 = rbit_1_1.ram_117_1.m0_s 
* net 3651 = rbit_1_1.ram_117_1.m1_s 
* net 3652 = rbit_1_1.ram_117_0.m0_s 
* net 3653 = rbit_1_1.ram_117_0.m1_s 
* net 3654 = rbit_1_1.ram_116_1.m0_s 
* net 3655 = rbit_1_1.ram_116_1.m1_s 
* net 3656 = rbit_1_1.ram_116_0.m0_s 
* net 3657 = rbit_1_1.ram_116_0.m1_s 
* net 3658 = rbit_1_1.ram_115_1.m0_s 
* net 3659 = rbit_1_1.ram_115_1.m1_s 
* net 3660 = rbit_1_1.ram_115_0.m0_s 
* net 3661 = rbit_1_1.ram_115_0.m1_s 
* net 3662 = rbit_1_1.ram_114_1.m0_s 
* net 3663 = rbit_1_1.ram_114_1.m1_s 
* net 3664 = rbit_1_1.ram_114_0.m0_s 
* net 3665 = rbit_1_1.ram_114_0.m1_s 
* net 3666 = rbit_1_1.ram_113_1.m0_s 
* net 3667 = rbit_1_1.ram_113_1.m1_s 
* net 3668 = rbit_1_1.ram_113_0.m0_s 
* net 3669 = rbit_1_1.ram_113_0.m1_s 
* net 3670 = rbit_1_1.ram_112_1.m0_s 
* net 3671 = rbit_1_1.ram_112_1.m1_s 
* net 3672 = rbit_1_1.ram_112_0.m0_s 
* net 3673 = rbit_1_1.ram_112_0.m1_s 
* net 3674 = rbit_1_1.ram_111_1.m0_s 
* net 3675 = rbit_1_1.ram_111_1.m1_s 
* net 3676 = rbit_1_1.ram_111_0.m0_s 
* net 3677 = rbit_1_1.ram_111_0.m1_s 
* net 3678 = rbit_1_1.ram_110_1.m0_s 
* net 3679 = rbit_1_1.ram_110_1.m1_s 
* net 3680 = rbit_1_1.ram_110_0.m0_s 
* net 3681 = rbit_1_1.ram_110_0.m1_s 
* net 3682 = rbit_1_1.ram_109_1.m0_s 
* net 3683 = rbit_1_1.ram_109_1.m1_s 
* net 3684 = rbit_1_1.ram_109_0.m0_s 
* net 3685 = rbit_1_1.ram_109_0.m1_s 
* net 3686 = rbit_1_1.ram_108_1.m0_s 
* net 3687 = rbit_1_1.ram_108_1.m1_s 
* net 3688 = rbit_1_1.ram_108_0.m0_s 
* net 3689 = rbit_1_1.ram_108_0.m1_s 
* net 3690 = rbit_1_1.ram_107_1.m0_s 
* net 3691 = rbit_1_1.ram_107_1.m1_s 
* net 3692 = rbit_1_1.ram_107_0.m0_s 
* net 3693 = rbit_1_1.ram_107_0.m1_s 
* net 3694 = rbit_1_1.ram_106_1.m0_s 
* net 3695 = rbit_1_1.ram_106_1.m1_s 
* net 3696 = rbit_1_1.ram_106_0.m0_s 
* net 3697 = rbit_1_1.ram_106_0.m1_s 
* net 3698 = rbit_1_1.ram_105_1.m0_s 
* net 3699 = rbit_1_1.ram_105_1.m1_s 
* net 3700 = rbit_1_1.ram_105_0.m0_s 
* net 3701 = rbit_1_1.ram_105_0.m1_s 
* net 3702 = rbit_1_1.ram_104_1.m0_s 
* net 3703 = rbit_1_1.ram_104_1.m1_s 
* net 3704 = rbit_1_1.ram_104_0.m0_s 
* net 3705 = rbit_1_1.ram_104_0.m1_s 
* net 3706 = rbit_1_1.ram_103_1.m0_s 
* net 3707 = rbit_1_1.ram_103_1.m1_s 
* net 3708 = rbit_1_1.ram_103_0.m0_s 
* net 3709 = rbit_1_1.ram_103_0.m1_s 
* net 3710 = rbit_1_1.ram_102_1.m0_s 
* net 3711 = rbit_1_1.ram_102_1.m1_s 
* net 3712 = rbit_1_1.ram_102_0.m0_s 
* net 3713 = rbit_1_1.ram_102_0.m1_s 
* net 3714 = rbit_1_1.ram_101_1.m0_s 
* net 3715 = rbit_1_1.ram_101_1.m1_s 
* net 3716 = rbit_1_1.ram_101_0.m0_s 
* net 3717 = rbit_1_1.ram_101_0.m1_s 
* net 3718 = rbit_1_1.ram_100_1.m0_s 
* net 3719 = rbit_1_1.ram_100_1.m1_s 
* net 3720 = rbit_1_1.ram_100_0.m0_s 
* net 3721 = rbit_1_1.ram_100_0.m1_s 
* net 3722 = rbit_1_1.ram_99_1.m0_s 
* net 3723 = rbit_1_1.ram_99_1.m1_s 
* net 3724 = rbit_1_1.ram_99_0.m0_s 
* net 3725 = rbit_1_1.ram_99_0.m1_s 
* net 3726 = rbit_1_1.ram_98_1.m0_s 
* net 3727 = rbit_1_1.ram_98_1.m1_s 
* net 3728 = rbit_1_1.ram_98_0.m0_s 
* net 3729 = rbit_1_1.ram_98_0.m1_s 
* net 3730 = rbit_1_1.ram_97_1.m0_s 
* net 3731 = rbit_1_1.ram_97_1.m1_s 
* net 3732 = rbit_1_1.ram_97_0.m0_s 
* net 3733 = rbit_1_1.ram_97_0.m1_s 
* net 3734 = rbit_1_1.ram_96_1.m0_s 
* net 3735 = rbit_1_1.ram_96_1.m1_s 
* net 3736 = rbit_1_1.ram_96_0.m0_s 
* net 3737 = rbit_1_1.ram_96_0.m1_s 
* net 3738 = rbit_1_1.ram_95_1.m0_s 
* net 3739 = rbit_1_1.ram_95_1.m1_s 
* net 3740 = rbit_1_1.ram_95_0.m0_s 
* net 3741 = rbit_1_1.ram_95_0.m1_s 
* net 3742 = rbit_1_1.ram_94_1.m0_s 
* net 3743 = rbit_1_1.ram_94_1.m1_s 
* net 3744 = rbit_1_1.ram_94_0.m0_s 
* net 3745 = rbit_1_1.ram_94_0.m1_s 
* net 3746 = rbit_1_1.ram_93_1.m0_s 
* net 3747 = rbit_1_1.ram_93_1.m1_s 
* net 3748 = rbit_1_1.ram_93_0.m0_s 
* net 3749 = rbit_1_1.ram_93_0.m1_s 
* net 3750 = rbit_1_1.ram_92_1.m0_s 
* net 3751 = rbit_1_1.ram_92_1.m1_s 
* net 3752 = rbit_1_1.ram_92_0.m0_s 
* net 3753 = rbit_1_1.ram_92_0.m1_s 
* net 3754 = rbit_1_1.ram_91_1.m0_s 
* net 3755 = rbit_1_1.ram_91_1.m1_s 
* net 3756 = rbit_1_1.ram_91_0.m0_s 
* net 3757 = rbit_1_1.ram_91_0.m1_s 
* net 3758 = rbit_1_1.ram_90_1.m0_s 
* net 3759 = rbit_1_1.ram_90_1.m1_s 
* net 3760 = rbit_1_1.ram_90_0.m0_s 
* net 3761 = rbit_1_1.ram_90_0.m1_s 
* net 3762 = rbit_1_1.ram_89_1.m0_s 
* net 3763 = rbit_1_1.ram_89_1.m1_s 
* net 3764 = rbit_1_1.ram_89_0.m0_s 
* net 3765 = rbit_1_1.ram_89_0.m1_s 
* net 3766 = rbit_1_1.ram_88_1.m0_s 
* net 3767 = rbit_1_1.ram_88_1.m1_s 
* net 3768 = rbit_1_1.ram_88_0.m0_s 
* net 3769 = rbit_1_1.ram_88_0.m1_s 
* net 3770 = rbit_1_1.ram_87_1.m0_s 
* net 3771 = rbit_1_1.ram_87_1.m1_s 
* net 3772 = rbit_1_1.ram_87_0.m0_s 
* net 3773 = rbit_1_1.ram_87_0.m1_s 
* net 3774 = rbit_1_1.ram_86_1.m0_s 
* net 3775 = rbit_1_1.ram_86_1.m1_s 
* net 3776 = rbit_1_1.ram_86_0.m0_s 
* net 3777 = rbit_1_1.ram_86_0.m1_s 
* net 3778 = rbit_1_1.ram_85_1.m0_s 
* net 3779 = rbit_1_1.ram_85_1.m1_s 
* net 3780 = rbit_1_1.ram_85_0.m0_s 
* net 3781 = rbit_1_1.ram_85_0.m1_s 
* net 3782 = rbit_1_1.ram_84_1.m0_s 
* net 3783 = rbit_1_1.ram_84_1.m1_s 
* net 3784 = rbit_1_1.ram_84_0.m0_s 
* net 3785 = rbit_1_1.ram_84_0.m1_s 
* net 3786 = rbit_1_1.ram_83_1.m0_s 
* net 3787 = rbit_1_1.ram_83_1.m1_s 
* net 3788 = rbit_1_1.ram_83_0.m0_s 
* net 3789 = rbit_1_1.ram_83_0.m1_s 
* net 3790 = rbit_1_1.ram_82_1.m0_s 
* net 3791 = rbit_1_1.ram_82_1.m1_s 
* net 3792 = rbit_1_1.ram_82_0.m0_s 
* net 3793 = rbit_1_1.ram_82_0.m1_s 
* net 3794 = rbit_1_1.ram_81_1.m0_s 
* net 3795 = rbit_1_1.ram_81_1.m1_s 
* net 3796 = rbit_1_1.ram_81_0.m0_s 
* net 3797 = rbit_1_1.ram_81_0.m1_s 
* net 3798 = rbit_1_1.ram_80_1.m0_s 
* net 3799 = rbit_1_1.ram_80_1.m1_s 
* net 3800 = rbit_1_1.ram_80_0.m0_s 
* net 3801 = rbit_1_1.ram_80_0.m1_s 
* net 3802 = rbit_1_1.ram_79_1.m0_s 
* net 3803 = rbit_1_1.ram_79_1.m1_s 
* net 3804 = rbit_1_1.ram_79_0.m0_s 
* net 3805 = rbit_1_1.ram_79_0.m1_s 
* net 3806 = rbit_1_1.ram_78_1.m0_s 
* net 3807 = rbit_1_1.ram_78_1.m1_s 
* net 3808 = rbit_1_1.ram_78_0.m0_s 
* net 3809 = rbit_1_1.ram_78_0.m1_s 
* net 3810 = rbit_1_1.ram_77_1.m0_s 
* net 3811 = rbit_1_1.ram_77_1.m1_s 
* net 3812 = rbit_1_1.ram_77_0.m0_s 
* net 3813 = rbit_1_1.ram_77_0.m1_s 
* net 3814 = rbit_1_1.ram_76_1.m0_s 
* net 3815 = rbit_1_1.ram_76_1.m1_s 
* net 3816 = rbit_1_1.ram_76_0.m0_s 
* net 3817 = rbit_1_1.ram_76_0.m1_s 
* net 3818 = rbit_1_1.ram_75_1.m0_s 
* net 3819 = rbit_1_1.ram_75_1.m1_s 
* net 3820 = rbit_1_1.ram_75_0.m0_s 
* net 3821 = rbit_1_1.ram_75_0.m1_s 
* net 3822 = rbit_1_1.ram_74_1.m0_s 
* net 3823 = rbit_1_1.ram_74_1.m1_s 
* net 3824 = rbit_1_1.ram_74_0.m0_s 
* net 3825 = rbit_1_1.ram_74_0.m1_s 
* net 3826 = rbit_1_1.ram_73_1.m0_s 
* net 3827 = rbit_1_1.ram_73_1.m1_s 
* net 3828 = rbit_1_1.ram_73_0.m0_s 
* net 3829 = rbit_1_1.ram_73_0.m1_s 
* net 3830 = rbit_1_1.ram_72_1.m0_s 
* net 3831 = rbit_1_1.ram_72_1.m1_s 
* net 3832 = rbit_1_1.ram_72_0.m0_s 
* net 3833 = rbit_1_1.ram_72_0.m1_s 
* net 3834 = rbit_1_1.ram_71_1.m0_s 
* net 3835 = rbit_1_1.ram_71_1.m1_s 
* net 3836 = rbit_1_1.ram_71_0.m0_s 
* net 3837 = rbit_1_1.ram_71_0.m1_s 
* net 3838 = rbit_1_1.ram_70_1.m0_s 
* net 3839 = rbit_1_1.ram_70_1.m1_s 
* net 3840 = rbit_1_1.ram_70_0.m0_s 
* net 3841 = rbit_1_1.ram_70_0.m1_s 
* net 3842 = rbit_1_1.ram_69_1.m0_s 
* net 3843 = rbit_1_1.ram_69_1.m1_s 
* net 3844 = rbit_1_1.ram_69_0.m0_s 
* net 3845 = rbit_1_1.ram_69_0.m1_s 
* net 3846 = rbit_1_1.ram_68_1.m0_s 
* net 3847 = rbit_1_1.ram_68_1.m1_s 
* net 3848 = rbit_1_1.ram_68_0.m0_s 
* net 3849 = rbit_1_1.ram_68_0.m1_s 
* net 3850 = rbit_1_1.ram_67_1.m0_s 
* net 3851 = rbit_1_1.ram_67_1.m1_s 
* net 3852 = rbit_1_1.ram_67_0.m0_s 
* net 3853 = rbit_1_1.ram_67_0.m1_s 
* net 3854 = rbit_1_1.ram_66_1.m0_s 
* net 3855 = rbit_1_1.ram_66_1.m1_s 
* net 3856 = rbit_1_1.ram_66_0.m0_s 
* net 3857 = rbit_1_1.ram_66_0.m1_s 
* net 3858 = rbit_1_1.ram_65_1.m0_s 
* net 3859 = rbit_1_1.ram_65_1.m1_s 
* net 3860 = rbit_1_1.ram_65_0.m0_s 
* net 3861 = rbit_1_1.ram_65_0.m1_s 
* net 3862 = rbit_1_1.ram_64_1.m0_s 
* net 3863 = rbit_1_1.ram_64_1.m1_s 
* net 3864 = rbit_1_1.ram_64_0.m0_s 
* net 3865 = rbit_1_1.ram_64_0.m1_s 
* net 3866 = rbit_1_1.ram_63_1.m0_s 
* net 3867 = rbit_1_1.ram_63_1.m1_s 
* net 3868 = rbit_1_1.ram_63_0.m0_s 
* net 3869 = rbit_1_1.ram_63_0.m1_s 
* net 3870 = rbit_1_1.ram_62_1.m0_s 
* net 3871 = rbit_1_1.ram_62_1.m1_s 
* net 3872 = rbit_1_1.ram_62_0.m0_s 
* net 3873 = rbit_1_1.ram_62_0.m1_s 
* net 3874 = rbit_1_1.ram_61_1.m0_s 
* net 3875 = rbit_1_1.ram_61_1.m1_s 
* net 3876 = rbit_1_1.ram_61_0.m0_s 
* net 3877 = rbit_1_1.ram_61_0.m1_s 
* net 3878 = rbit_1_1.ram_60_1.m0_s 
* net 3879 = rbit_1_1.ram_60_1.m1_s 
* net 3880 = rbit_1_1.ram_60_0.m0_s 
* net 3881 = rbit_1_1.ram_60_0.m1_s 
* net 3882 = rbit_1_1.ram_59_1.m0_s 
* net 3883 = rbit_1_1.ram_59_1.m1_s 
* net 3884 = rbit_1_1.ram_59_0.m0_s 
* net 3885 = rbit_1_1.ram_59_0.m1_s 
* net 3886 = rbit_1_1.ram_58_1.m0_s 
* net 3887 = rbit_1_1.ram_58_1.m1_s 
* net 3888 = rbit_1_1.ram_58_0.m0_s 
* net 3889 = rbit_1_1.ram_58_0.m1_s 
* net 3890 = rbit_1_1.ram_57_1.m0_s 
* net 3891 = rbit_1_1.ram_57_1.m1_s 
* net 3892 = rbit_1_1.ram_57_0.m0_s 
* net 3893 = rbit_1_1.ram_57_0.m1_s 
* net 3894 = rbit_1_1.ram_56_1.m0_s 
* net 3895 = rbit_1_1.ram_56_1.m1_s 
* net 3896 = rbit_1_1.ram_56_0.m0_s 
* net 3897 = rbit_1_1.ram_56_0.m1_s 
* net 3898 = rbit_1_1.ram_55_1.m0_s 
* net 3899 = rbit_1_1.ram_55_1.m1_s 
* net 3900 = rbit_1_1.ram_55_0.m0_s 
* net 3901 = rbit_1_1.ram_55_0.m1_s 
* net 3902 = rbit_1_1.ram_54_1.m0_s 
* net 3903 = rbit_1_1.ram_54_1.m1_s 
* net 3904 = rbit_1_1.ram_54_0.m0_s 
* net 3905 = rbit_1_1.ram_54_0.m1_s 
* net 3906 = rbit_1_1.ram_53_1.m0_s 
* net 3907 = rbit_1_1.ram_53_1.m1_s 
* net 3908 = rbit_1_1.ram_53_0.m0_s 
* net 3909 = rbit_1_1.ram_53_0.m1_s 
* net 3910 = rbit_1_1.ram_52_1.m0_s 
* net 3911 = rbit_1_1.ram_52_1.m1_s 
* net 3912 = rbit_1_1.ram_52_0.m0_s 
* net 3913 = rbit_1_1.ram_52_0.m1_s 
* net 3914 = rbit_1_1.ram_51_1.m0_s 
* net 3915 = rbit_1_1.ram_51_1.m1_s 
* net 3916 = rbit_1_1.ram_51_0.m0_s 
* net 3917 = rbit_1_1.ram_51_0.m1_s 
* net 3918 = rbit_1_1.ram_50_1.m0_s 
* net 3919 = rbit_1_1.ram_50_1.m1_s 
* net 3920 = rbit_1_1.ram_50_0.m0_s 
* net 3921 = rbit_1_1.ram_50_0.m1_s 
* net 3922 = rbit_1_1.ram_49_1.m0_s 
* net 3923 = rbit_1_1.ram_49_1.m1_s 
* net 3924 = rbit_1_1.ram_49_0.m0_s 
* net 3925 = rbit_1_1.ram_49_0.m1_s 
* net 3926 = rbit_1_1.ram_48_1.m0_s 
* net 3927 = rbit_1_1.ram_48_1.m1_s 
* net 3928 = rbit_1_1.ram_48_0.m0_s 
* net 3929 = rbit_1_1.ram_48_0.m1_s 
* net 3930 = rbit_1_1.ram_47_1.m0_s 
* net 3931 = rbit_1_1.ram_47_1.m1_s 
* net 3932 = rbit_1_1.ram_47_0.m0_s 
* net 3933 = rbit_1_1.ram_47_0.m1_s 
* net 3934 = rbit_1_1.ram_46_1.m0_s 
* net 3935 = rbit_1_1.ram_46_1.m1_s 
* net 3936 = rbit_1_1.ram_46_0.m0_s 
* net 3937 = rbit_1_1.ram_46_0.m1_s 
* net 3938 = rbit_1_1.ram_45_1.m0_s 
* net 3939 = rbit_1_1.ram_45_1.m1_s 
* net 3940 = rbit_1_1.ram_45_0.m0_s 
* net 3941 = rbit_1_1.ram_45_0.m1_s 
* net 3942 = rbit_1_1.ram_44_1.m0_s 
* net 3943 = rbit_1_1.ram_44_1.m1_s 
* net 3944 = rbit_1_1.ram_44_0.m0_s 
* net 3945 = rbit_1_1.ram_44_0.m1_s 
* net 3946 = rbit_1_1.ram_43_1.m0_s 
* net 3947 = rbit_1_1.ram_43_1.m1_s 
* net 3948 = rbit_1_1.ram_43_0.m0_s 
* net 3949 = rbit_1_1.ram_43_0.m1_s 
* net 3950 = rbit_1_1.ram_42_1.m0_s 
* net 3951 = rbit_1_1.ram_42_1.m1_s 
* net 3952 = rbit_1_1.ram_42_0.m0_s 
* net 3953 = rbit_1_1.ram_42_0.m1_s 
* net 3954 = rbit_1_1.ram_41_1.m0_s 
* net 3955 = rbit_1_1.ram_41_1.m1_s 
* net 3956 = rbit_1_1.ram_41_0.m0_s 
* net 3957 = rbit_1_1.ram_41_0.m1_s 
* net 3958 = rbit_1_1.ram_40_1.m0_s 
* net 3959 = rbit_1_1.ram_40_1.m1_s 
* net 3960 = rbit_1_1.ram_40_0.m0_s 
* net 3961 = rbit_1_1.ram_40_0.m1_s 
* net 3962 = rbit_1_1.ram_39_1.m0_s 
* net 3963 = rbit_1_1.ram_39_1.m1_s 
* net 3964 = rbit_1_1.ram_39_0.m0_s 
* net 3965 = rbit_1_1.ram_39_0.m1_s 
* net 3966 = rbit_1_1.ram_38_1.m0_s 
* net 3967 = rbit_1_1.ram_38_1.m1_s 
* net 3968 = rbit_1_1.ram_38_0.m0_s 
* net 3969 = rbit_1_1.ram_38_0.m1_s 
* net 3970 = rbit_1_1.ram_37_1.m0_s 
* net 3971 = rbit_1_1.ram_37_1.m1_s 
* net 3972 = rbit_1_1.ram_37_0.m0_s 
* net 3973 = rbit_1_1.ram_37_0.m1_s 
* net 3974 = rbit_1_1.ram_36_1.m0_s 
* net 3975 = rbit_1_1.ram_36_1.m1_s 
* net 3976 = rbit_1_1.ram_36_0.m0_s 
* net 3977 = rbit_1_1.ram_36_0.m1_s 
* net 3978 = rbit_1_1.ram_35_1.m0_s 
* net 3979 = rbit_1_1.ram_35_1.m1_s 
* net 3980 = rbit_1_1.ram_35_0.m0_s 
* net 3981 = rbit_1_1.ram_35_0.m1_s 
* net 3982 = rbit_1_1.ram_34_1.m0_s 
* net 3983 = rbit_1_1.ram_34_1.m1_s 
* net 3984 = rbit_1_1.ram_34_0.m0_s 
* net 3985 = rbit_1_1.ram_34_0.m1_s 
* net 3986 = rbit_1_1.ram_33_1.m0_s 
* net 3987 = rbit_1_1.ram_33_1.m1_s 
* net 3988 = rbit_1_1.ram_33_0.m0_s 
* net 3989 = rbit_1_1.ram_33_0.m1_s 
* net 3990 = rbit_1_1.ram_32_1.m0_s 
* net 3991 = rbit_1_1.ram_32_1.m1_s 
* net 3992 = rbit_1_1.ram_32_0.m0_s 
* net 3993 = rbit_1_1.ram_32_0.m1_s 
* net 3994 = rbit_1_1.ram_31_1.m0_s 
* net 3995 = rbit_1_1.ram_31_1.m1_s 
* net 3996 = rbit_1_1.ram_31_0.m0_s 
* net 3997 = rbit_1_1.ram_31_0.m1_s 
* net 3998 = rbit_1_1.ram_30_1.m0_s 
* net 3999 = rbit_1_1.ram_30_1.m1_s 
* net 4000 = rbit_1_1.ram_30_0.m0_s 
* net 4001 = rbit_1_1.ram_30_0.m1_s 
* net 4002 = rbit_1_1.ram_29_1.m0_s 
* net 4003 = rbit_1_1.ram_29_1.m1_s 
* net 4004 = rbit_1_1.ram_29_0.m0_s 
* net 4005 = rbit_1_1.ram_29_0.m1_s 
* net 4006 = rbit_1_1.ram_28_1.m0_s 
* net 4007 = rbit_1_1.ram_28_1.m1_s 
* net 4008 = rbit_1_1.ram_28_0.m0_s 
* net 4009 = rbit_1_1.ram_28_0.m1_s 
* net 4010 = rbit_1_1.ram_27_1.m0_s 
* net 4011 = rbit_1_1.ram_27_1.m1_s 
* net 4012 = rbit_1_1.ram_27_0.m0_s 
* net 4013 = rbit_1_1.ram_27_0.m1_s 
* net 4014 = rbit_1_1.ram_26_1.m0_s 
* net 4015 = rbit_1_1.ram_26_1.m1_s 
* net 4016 = rbit_1_1.ram_26_0.m0_s 
* net 4017 = rbit_1_1.ram_26_0.m1_s 
* net 4018 = rbit_1_1.ram_25_1.m0_s 
* net 4019 = rbit_1_1.ram_25_1.m1_s 
* net 4020 = rbit_1_1.ram_25_0.m0_s 
* net 4021 = rbit_1_1.ram_25_0.m1_s 
* net 4022 = rbit_1_1.ram_24_1.m0_s 
* net 4023 = rbit_1_1.ram_24_1.m1_s 
* net 4024 = rbit_1_1.ram_24_0.m0_s 
* net 4025 = rbit_1_1.ram_24_0.m1_s 
* net 4026 = rbit_1_1.ram_23_1.m0_s 
* net 4027 = rbit_1_1.ram_23_1.m1_s 
* net 4028 = rbit_1_1.ram_23_0.m0_s 
* net 4029 = rbit_1_1.ram_23_0.m1_s 
* net 4030 = rbit_1_1.ram_22_1.m0_s 
* net 4031 = rbit_1_1.ram_22_1.m1_s 
* net 4032 = rbit_1_1.ram_22_0.m0_s 
* net 4033 = rbit_1_1.ram_22_0.m1_s 
* net 4034 = rbit_1_1.ram_21_1.m0_s 
* net 4035 = rbit_1_1.ram_21_1.m1_s 
* net 4036 = rbit_1_1.ram_21_0.m0_s 
* net 4037 = rbit_1_1.ram_21_0.m1_s 
* net 4038 = rbit_1_1.ram_20_1.m0_s 
* net 4039 = rbit_1_1.ram_20_1.m1_s 
* net 4040 = rbit_1_1.ram_20_0.m0_s 
* net 4041 = rbit_1_1.ram_20_0.m1_s 
* net 4042 = rbit_1_1.ram_19_1.m0_s 
* net 4043 = rbit_1_1.ram_19_1.m1_s 
* net 4044 = rbit_1_1.ram_19_0.m0_s 
* net 4045 = rbit_1_1.ram_19_0.m1_s 
* net 4046 = rbit_1_1.ram_18_1.m0_s 
* net 4047 = rbit_1_1.ram_18_1.m1_s 
* net 4048 = rbit_1_1.ram_18_0.m0_s 
* net 4049 = rbit_1_1.ram_18_0.m1_s 
* net 4050 = rbit_1_1.ram_17_1.m0_s 
* net 4051 = rbit_1_1.ram_17_1.m1_s 
* net 4052 = rbit_1_1.ram_17_0.m0_s 
* net 4053 = rbit_1_1.ram_17_0.m1_s 
* net 4054 = rbit_1_1.ram_16_1.m0_s 
* net 4055 = rbit_1_1.ram_16_1.m1_s 
* net 4056 = rbit_1_1.ram_16_0.m0_s 
* net 4057 = rbit_1_1.ram_16_0.m1_s 
* net 4058 = rbit_1_1.ram_15_1.m0_s 
* net 4059 = rbit_1_1.ram_15_1.m1_s 
* net 4060 = rbit_1_1.ram_15_0.m0_s 
* net 4061 = rbit_1_1.ram_15_0.m1_s 
* net 4062 = rbit_1_1.ram_14_1.m0_s 
* net 4063 = rbit_1_1.ram_14_1.m1_s 
* net 4064 = rbit_1_1.ram_14_0.m0_s 
* net 4065 = rbit_1_1.ram_14_0.m1_s 
* net 4066 = rbit_1_1.ram_13_1.m0_s 
* net 4067 = rbit_1_1.ram_13_1.m1_s 
* net 4068 = rbit_1_1.ram_13_0.m0_s 
* net 4069 = rbit_1_1.ram_13_0.m1_s 
* net 4070 = rbit_1_1.ram_12_1.m0_s 
* net 4071 = rbit_1_1.ram_12_1.m1_s 
* net 4072 = rbit_1_1.ram_12_0.m0_s 
* net 4073 = rbit_1_1.ram_12_0.m1_s 
* net 4074 = rbit_1_1.ram_11_1.m0_s 
* net 4075 = rbit_1_1.ram_11_1.m1_s 
* net 4076 = rbit_1_1.ram_11_0.m0_s 
* net 4077 = rbit_1_1.ram_11_0.m1_s 
* net 4078 = rbit_1_1.ram_10_1.m0_s 
* net 4079 = rbit_1_1.ram_10_1.m1_s 
* net 4080 = rbit_1_1.ram_10_0.m0_s 
* net 4081 = rbit_1_1.ram_10_0.m1_s 
* net 4082 = rbit_1_1.ram_9_1.m0_s 
* net 4083 = rbit_1_1.ram_9_1.m1_s 
* net 4084 = rbit_1_1.ram_9_0.m0_s 
* net 4085 = rbit_1_1.ram_9_0.m1_s 
* net 4086 = rbit_1_1.ram_8_1.m0_s 
* net 4087 = rbit_1_1.ram_8_1.m1_s 
* net 4088 = rbit_1_1.ram_8_0.m0_s 
* net 4089 = rbit_1_1.ram_8_0.m1_s 
* net 4090 = rbit_1_1.ram_7_1.m0_s 
* net 4091 = rbit_1_1.ram_7_1.m1_s 
* net 4092 = rbit_1_1.ram_7_0.m0_s 
* net 4093 = rbit_1_1.ram_7_0.m1_s 
* net 4094 = rbit_1_1.ram_6_1.m0_s 
* net 4095 = rbit_1_1.ram_6_1.m1_s 
* net 4096 = rbit_1_1.ram_6_0.m0_s 
* net 4097 = rbit_1_1.ram_6_0.m1_s 
* net 4098 = rbit_1_1.ram_5_1.m0_s 
* net 4099 = rbit_1_1.ram_5_1.m1_s 
* net 4100 = rbit_1_1.ram_5_0.m0_s 
* net 4101 = rbit_1_1.ram_5_0.m1_s 
* net 4102 = rbit_1_1.ram_4_1.m0_s 
* net 4103 = rbit_1_1.ram_4_1.m1_s 
* net 4104 = rbit_1_1.ram_4_0.m0_s 
* net 4105 = rbit_1_1.ram_4_0.m1_s 
* net 4106 = rbit_1_1.ram_3_1.m0_s 
* net 4107 = rbit_1_1.ram_3_1.m1_s 
* net 4108 = rbit_1_1.ram_3_0.m0_s 
* net 4109 = rbit_1_1.ram_3_0.m1_s 
* net 4110 = rbit_1_1.ram_2_1.m0_s 
* net 4111 = rbit_1_1.ram_2_1.m1_s 
* net 4112 = rbit_1_1.ram_2_0.m0_s 
* net 4113 = rbit_1_1.ram_2_0.m1_s 
* net 4114 = rbit_1_1.ram_1_1.m0_s 
* net 4115 = rbit_1_1.ram_1_1.m1_s 
* net 4116 = rbit_1_1.ram_1_0.m0_s 
* net 4117 = rbit_1_1.ram_1_0.m1_s 
* net 4118 = rbit_1_1.ram_0_1.m0_s 
* net 4119 = rbit_1_1.ram_0_1.m1_s 
* net 4120 = rbit_1_1.ram_0_0.m0_s 
* net 4121 = rbit_1_1.ram_0_0.m1_s 
* net 4122 = mbk_sig149 
* net 4123 = mbk_sig127 
* net 4124 = mbk_sig172 
* net 4125 = mbk_sig126 
* net 4126 = mbk_sig189 
* net 4127 = mbk_sig49 
* net 4128 = mbk_sig47 
* net 4129 = mbk_sig77 
* net 4130 = mbk_sig103 
* net 4131 = mbk_sig95 
* net 4132 = mbk_sig87 
* net 4133 = rbit_2_1.ram_127_1.m0_s 
* net 4134 = rbit_2_1.ram_127_1.m1_s 
* net 4135 = rbit_2_1.ram_127_0.m0_s 
* net 4136 = rbit_2_1.ram_127_0.m1_s 
* net 4137 = rbit_2_1.ram_126_1.m0_s 
* net 4138 = rbit_2_1.ram_126_1.m1_s 
* net 4139 = rbit_2_1.ram_126_0.m0_s 
* net 4140 = rbit_2_1.ram_126_0.m1_s 
* net 4141 = rbit_2_1.ram_125_1.m0_s 
* net 4142 = rbit_2_1.ram_125_1.m1_s 
* net 4143 = rbit_2_1.ram_125_0.m0_s 
* net 4144 = rbit_2_1.ram_125_0.m1_s 
* net 4145 = rbit_2_1.ram_124_1.m0_s 
* net 4146 = rbit_2_1.ram_124_1.m1_s 
* net 4147 = rbit_2_1.ram_124_0.m0_s 
* net 4148 = rbit_2_1.ram_124_0.m1_s 
* net 4149 = rbit_2_1.ram_123_1.m0_s 
* net 4150 = rbit_2_1.ram_123_1.m1_s 
* net 4151 = rbit_2_1.ram_123_0.m0_s 
* net 4152 = rbit_2_1.ram_123_0.m1_s 
* net 4153 = rbit_2_1.ram_122_1.m0_s 
* net 4154 = rbit_2_1.ram_122_1.m1_s 
* net 4155 = rbit_2_1.ram_122_0.m0_s 
* net 4156 = rbit_2_1.ram_122_0.m1_s 
* net 4157 = rbit_2_1.ram_121_1.m0_s 
* net 4158 = rbit_2_1.ram_121_1.m1_s 
* net 4159 = rbit_2_1.ram_121_0.m0_s 
* net 4160 = rbit_2_1.ram_121_0.m1_s 
* net 4161 = rbit_2_1.ram_120_1.m0_s 
* net 4162 = rbit_2_1.ram_120_1.m1_s 
* net 4163 = rbit_2_1.ram_120_0.m0_s 
* net 4164 = rbit_2_1.ram_120_0.m1_s 
* net 4165 = rbit_2_1.ram_119_1.m0_s 
* net 4166 = rbit_2_1.ram_119_1.m1_s 
* net 4167 = rbit_2_1.ram_119_0.m0_s 
* net 4168 = rbit_2_1.ram_119_0.m1_s 
* net 4169 = rbit_2_1.ram_118_1.m0_s 
* net 4170 = rbit_2_1.ram_118_1.m1_s 
* net 4171 = rbit_2_1.ram_118_0.m0_s 
* net 4172 = rbit_2_1.ram_118_0.m1_s 
* net 4173 = rbit_2_1.ram_117_1.m0_s 
* net 4174 = rbit_2_1.ram_117_1.m1_s 
* net 4175 = rbit_2_1.ram_117_0.m0_s 
* net 4176 = rbit_2_1.ram_117_0.m1_s 
* net 4177 = rbit_2_1.ram_116_1.m0_s 
* net 4178 = rbit_2_1.ram_116_1.m1_s 
* net 4179 = rbit_2_1.ram_116_0.m0_s 
* net 4180 = rbit_2_1.ram_116_0.m1_s 
* net 4181 = rbit_2_1.ram_115_1.m0_s 
* net 4182 = rbit_2_1.ram_115_1.m1_s 
* net 4183 = rbit_2_1.ram_115_0.m0_s 
* net 4184 = rbit_2_1.ram_115_0.m1_s 
* net 4185 = rbit_2_1.ram_114_1.m0_s 
* net 4186 = rbit_2_1.ram_114_1.m1_s 
* net 4187 = rbit_2_1.ram_114_0.m0_s 
* net 4188 = rbit_2_1.ram_114_0.m1_s 
* net 4189 = rbit_2_1.ram_113_1.m0_s 
* net 4190 = rbit_2_1.ram_113_1.m1_s 
* net 4191 = rbit_2_1.ram_113_0.m0_s 
* net 4192 = rbit_2_1.ram_113_0.m1_s 
* net 4193 = rbit_2_1.ram_112_1.m0_s 
* net 4194 = rbit_2_1.ram_112_1.m1_s 
* net 4195 = rbit_2_1.ram_112_0.m0_s 
* net 4196 = rbit_2_1.ram_112_0.m1_s 
* net 4197 = rbit_2_1.ram_111_1.m0_s 
* net 4198 = rbit_2_1.ram_111_1.m1_s 
* net 4199 = rbit_2_1.ram_111_0.m0_s 
* net 4200 = rbit_2_1.ram_111_0.m1_s 
* net 4201 = rbit_2_1.ram_110_1.m0_s 
* net 4202 = rbit_2_1.ram_110_1.m1_s 
* net 4203 = rbit_2_1.ram_110_0.m0_s 
* net 4204 = rbit_2_1.ram_110_0.m1_s 
* net 4205 = rbit_2_1.ram_109_1.m0_s 
* net 4206 = rbit_2_1.ram_109_1.m1_s 
* net 4207 = rbit_2_1.ram_109_0.m0_s 
* net 4208 = rbit_2_1.ram_109_0.m1_s 
* net 4209 = rbit_2_1.ram_108_1.m0_s 
* net 4210 = rbit_2_1.ram_108_1.m1_s 
* net 4211 = rbit_2_1.ram_108_0.m0_s 
* net 4212 = rbit_2_1.ram_108_0.m1_s 
* net 4213 = rbit_2_1.ram_107_1.m0_s 
* net 4214 = rbit_2_1.ram_107_1.m1_s 
* net 4215 = rbit_2_1.ram_107_0.m0_s 
* net 4216 = rbit_2_1.ram_107_0.m1_s 
* net 4217 = rbit_2_1.ram_106_1.m0_s 
* net 4218 = rbit_2_1.ram_106_1.m1_s 
* net 4219 = rbit_2_1.ram_106_0.m0_s 
* net 4220 = rbit_2_1.ram_106_0.m1_s 
* net 4221 = rbit_2_1.ram_105_1.m0_s 
* net 4222 = rbit_2_1.ram_105_1.m1_s 
* net 4223 = rbit_2_1.ram_105_0.m0_s 
* net 4224 = rbit_2_1.ram_105_0.m1_s 
* net 4225 = rbit_2_1.ram_104_1.m0_s 
* net 4226 = rbit_2_1.ram_104_1.m1_s 
* net 4227 = rbit_2_1.ram_104_0.m0_s 
* net 4228 = rbit_2_1.ram_104_0.m1_s 
* net 4229 = rbit_2_1.ram_103_1.m0_s 
* net 4230 = rbit_2_1.ram_103_1.m1_s 
* net 4231 = rbit_2_1.ram_103_0.m0_s 
* net 4232 = rbit_2_1.ram_103_0.m1_s 
* net 4233 = rbit_2_1.ram_102_1.m0_s 
* net 4234 = rbit_2_1.ram_102_1.m1_s 
* net 4235 = rbit_2_1.ram_102_0.m0_s 
* net 4236 = rbit_2_1.ram_102_0.m1_s 
* net 4237 = rbit_2_1.ram_101_1.m0_s 
* net 4238 = rbit_2_1.ram_101_1.m1_s 
* net 4239 = rbit_2_1.ram_101_0.m0_s 
* net 4240 = rbit_2_1.ram_101_0.m1_s 
* net 4241 = rbit_2_1.ram_100_1.m0_s 
* net 4242 = rbit_2_1.ram_100_1.m1_s 
* net 4243 = rbit_2_1.ram_100_0.m0_s 
* net 4244 = rbit_2_1.ram_100_0.m1_s 
* net 4245 = rbit_2_1.ram_99_1.m0_s 
* net 4246 = rbit_2_1.ram_99_1.m1_s 
* net 4247 = rbit_2_1.ram_99_0.m0_s 
* net 4248 = rbit_2_1.ram_99_0.m1_s 
* net 4249 = rbit_2_1.ram_98_1.m0_s 
* net 4250 = rbit_2_1.ram_98_1.m1_s 
* net 4251 = rbit_2_1.ram_98_0.m0_s 
* net 4252 = rbit_2_1.ram_98_0.m1_s 
* net 4253 = rbit_2_1.ram_97_1.m0_s 
* net 4254 = rbit_2_1.ram_97_1.m1_s 
* net 4255 = rbit_2_1.ram_97_0.m0_s 
* net 4256 = rbit_2_1.ram_97_0.m1_s 
* net 4257 = rbit_2_1.ram_96_1.m0_s 
* net 4258 = rbit_2_1.ram_96_1.m1_s 
* net 4259 = rbit_2_1.ram_96_0.m0_s 
* net 4260 = rbit_2_1.ram_96_0.m1_s 
* net 4261 = rbit_2_1.ram_95_1.m0_s 
* net 4262 = rbit_2_1.ram_95_1.m1_s 
* net 4263 = rbit_2_1.ram_95_0.m0_s 
* net 4264 = rbit_2_1.ram_95_0.m1_s 
* net 4265 = rbit_2_1.ram_94_1.m0_s 
* net 4266 = rbit_2_1.ram_94_1.m1_s 
* net 4267 = rbit_2_1.ram_94_0.m0_s 
* net 4268 = rbit_2_1.ram_94_0.m1_s 
* net 4269 = rbit_2_1.ram_93_1.m0_s 
* net 4270 = rbit_2_1.ram_93_1.m1_s 
* net 4271 = rbit_2_1.ram_93_0.m0_s 
* net 4272 = rbit_2_1.ram_93_0.m1_s 
* net 4273 = rbit_2_1.ram_92_1.m0_s 
* net 4274 = rbit_2_1.ram_92_1.m1_s 
* net 4275 = rbit_2_1.ram_92_0.m0_s 
* net 4276 = rbit_2_1.ram_92_0.m1_s 
* net 4277 = rbit_2_1.ram_91_1.m0_s 
* net 4278 = rbit_2_1.ram_91_1.m1_s 
* net 4279 = rbit_2_1.ram_91_0.m0_s 
* net 4280 = rbit_2_1.ram_91_0.m1_s 
* net 4281 = rbit_2_1.ram_90_1.m0_s 
* net 4282 = rbit_2_1.ram_90_1.m1_s 
* net 4283 = rbit_2_1.ram_90_0.m0_s 
* net 4284 = rbit_2_1.ram_90_0.m1_s 
* net 4285 = rbit_2_1.ram_89_1.m0_s 
* net 4286 = rbit_2_1.ram_89_1.m1_s 
* net 4287 = rbit_2_1.ram_89_0.m0_s 
* net 4288 = rbit_2_1.ram_89_0.m1_s 
* net 4289 = rbit_2_1.ram_88_1.m0_s 
* net 4290 = rbit_2_1.ram_88_1.m1_s 
* net 4291 = rbit_2_1.ram_88_0.m0_s 
* net 4292 = rbit_2_1.ram_88_0.m1_s 
* net 4293 = rbit_2_1.ram_87_1.m0_s 
* net 4294 = rbit_2_1.ram_87_1.m1_s 
* net 4295 = rbit_2_1.ram_87_0.m0_s 
* net 4296 = rbit_2_1.ram_87_0.m1_s 
* net 4297 = rbit_2_1.ram_86_1.m0_s 
* net 4298 = rbit_2_1.ram_86_1.m1_s 
* net 4299 = rbit_2_1.ram_86_0.m0_s 
* net 4300 = rbit_2_1.ram_86_0.m1_s 
* net 4301 = rbit_2_1.ram_85_1.m0_s 
* net 4302 = rbit_2_1.ram_85_1.m1_s 
* net 4303 = rbit_2_1.ram_85_0.m0_s 
* net 4304 = rbit_2_1.ram_85_0.m1_s 
* net 4305 = rbit_2_1.ram_84_1.m0_s 
* net 4306 = rbit_2_1.ram_84_1.m1_s 
* net 4307 = rbit_2_1.ram_84_0.m0_s 
* net 4308 = rbit_2_1.ram_84_0.m1_s 
* net 4309 = rbit_2_1.ram_83_1.m0_s 
* net 4310 = rbit_2_1.ram_83_1.m1_s 
* net 4311 = rbit_2_1.ram_83_0.m0_s 
* net 4312 = rbit_2_1.ram_83_0.m1_s 
* net 4313 = rbit_2_1.ram_82_1.m0_s 
* net 4314 = rbit_2_1.ram_82_1.m1_s 
* net 4315 = rbit_2_1.ram_82_0.m0_s 
* net 4316 = rbit_2_1.ram_82_0.m1_s 
* net 4317 = rbit_2_1.ram_81_1.m0_s 
* net 4318 = rbit_2_1.ram_81_1.m1_s 
* net 4319 = rbit_2_1.ram_81_0.m0_s 
* net 4320 = rbit_2_1.ram_81_0.m1_s 
* net 4321 = rbit_2_1.ram_80_1.m0_s 
* net 4322 = rbit_2_1.ram_80_1.m1_s 
* net 4323 = rbit_2_1.ram_80_0.m0_s 
* net 4324 = rbit_2_1.ram_80_0.m1_s 
* net 4325 = rbit_2_1.ram_79_1.m0_s 
* net 4326 = rbit_2_1.ram_79_1.m1_s 
* net 4327 = rbit_2_1.ram_79_0.m0_s 
* net 4328 = rbit_2_1.ram_79_0.m1_s 
* net 4329 = rbit_2_1.ram_78_1.m0_s 
* net 4330 = rbit_2_1.ram_78_1.m1_s 
* net 4331 = rbit_2_1.ram_78_0.m0_s 
* net 4332 = rbit_2_1.ram_78_0.m1_s 
* net 4333 = rbit_2_1.ram_77_1.m0_s 
* net 4334 = rbit_2_1.ram_77_1.m1_s 
* net 4335 = rbit_2_1.ram_77_0.m0_s 
* net 4336 = rbit_2_1.ram_77_0.m1_s 
* net 4337 = rbit_2_1.ram_76_1.m0_s 
* net 4338 = rbit_2_1.ram_76_1.m1_s 
* net 4339 = rbit_2_1.ram_76_0.m0_s 
* net 4340 = rbit_2_1.ram_76_0.m1_s 
* net 4341 = rbit_2_1.ram_75_1.m0_s 
* net 4342 = rbit_2_1.ram_75_1.m1_s 
* net 4343 = rbit_2_1.ram_75_0.m0_s 
* net 4344 = rbit_2_1.ram_75_0.m1_s 
* net 4345 = rbit_2_1.ram_74_1.m0_s 
* net 4346 = rbit_2_1.ram_74_1.m1_s 
* net 4347 = rbit_2_1.ram_74_0.m0_s 
* net 4348 = rbit_2_1.ram_74_0.m1_s 
* net 4349 = rbit_2_1.ram_73_1.m0_s 
* net 4350 = rbit_2_1.ram_73_1.m1_s 
* net 4351 = rbit_2_1.ram_73_0.m0_s 
* net 4352 = rbit_2_1.ram_73_0.m1_s 
* net 4353 = rbit_2_1.ram_72_1.m0_s 
* net 4354 = rbit_2_1.ram_72_1.m1_s 
* net 4355 = rbit_2_1.ram_72_0.m0_s 
* net 4356 = rbit_2_1.ram_72_0.m1_s 
* net 4357 = rbit_2_1.ram_71_1.m0_s 
* net 4358 = rbit_2_1.ram_71_1.m1_s 
* net 4359 = rbit_2_1.ram_71_0.m0_s 
* net 4360 = rbit_2_1.ram_71_0.m1_s 
* net 4361 = rbit_2_1.ram_70_1.m0_s 
* net 4362 = rbit_2_1.ram_70_1.m1_s 
* net 4363 = rbit_2_1.ram_70_0.m0_s 
* net 4364 = rbit_2_1.ram_70_0.m1_s 
* net 4365 = rbit_2_1.ram_69_1.m0_s 
* net 4366 = rbit_2_1.ram_69_1.m1_s 
* net 4367 = rbit_2_1.ram_69_0.m0_s 
* net 4368 = rbit_2_1.ram_69_0.m1_s 
* net 4369 = rbit_2_1.ram_68_1.m0_s 
* net 4370 = rbit_2_1.ram_68_1.m1_s 
* net 4371 = rbit_2_1.ram_68_0.m0_s 
* net 4372 = rbit_2_1.ram_68_0.m1_s 
* net 4373 = rbit_2_1.ram_67_1.m0_s 
* net 4374 = rbit_2_1.ram_67_1.m1_s 
* net 4375 = rbit_2_1.ram_67_0.m0_s 
* net 4376 = rbit_2_1.ram_67_0.m1_s 
* net 4377 = rbit_2_1.ram_66_1.m0_s 
* net 4378 = rbit_2_1.ram_66_1.m1_s 
* net 4379 = rbit_2_1.ram_66_0.m0_s 
* net 4380 = rbit_2_1.ram_66_0.m1_s 
* net 4381 = rbit_2_1.ram_65_1.m0_s 
* net 4382 = rbit_2_1.ram_65_1.m1_s 
* net 4383 = rbit_2_1.ram_65_0.m0_s 
* net 4384 = rbit_2_1.ram_65_0.m1_s 
* net 4385 = rbit_2_1.ram_64_1.m0_s 
* net 4386 = rbit_2_1.ram_64_1.m1_s 
* net 4387 = rbit_2_1.ram_64_0.m0_s 
* net 4388 = rbit_2_1.ram_64_0.m1_s 
* net 4389 = rbit_2_1.ram_63_1.m0_s 
* net 4390 = rbit_2_1.ram_63_1.m1_s 
* net 4391 = rbit_2_1.ram_63_0.m0_s 
* net 4392 = rbit_2_1.ram_63_0.m1_s 
* net 4393 = rbit_2_1.ram_62_1.m0_s 
* net 4394 = rbit_2_1.ram_62_1.m1_s 
* net 4395 = rbit_2_1.ram_62_0.m0_s 
* net 4396 = rbit_2_1.ram_62_0.m1_s 
* net 4397 = rbit_2_1.ram_61_1.m0_s 
* net 4398 = rbit_2_1.ram_61_1.m1_s 
* net 4399 = rbit_2_1.ram_61_0.m0_s 
* net 4400 = rbit_2_1.ram_61_0.m1_s 
* net 4401 = rbit_2_1.ram_60_1.m0_s 
* net 4402 = rbit_2_1.ram_60_1.m1_s 
* net 4403 = rbit_2_1.ram_60_0.m0_s 
* net 4404 = rbit_2_1.ram_60_0.m1_s 
* net 4405 = rbit_2_1.ram_59_1.m0_s 
* net 4406 = rbit_2_1.ram_59_1.m1_s 
* net 4407 = rbit_2_1.ram_59_0.m0_s 
* net 4408 = rbit_2_1.ram_59_0.m1_s 
* net 4409 = rbit_2_1.ram_58_1.m0_s 
* net 4410 = rbit_2_1.ram_58_1.m1_s 
* net 4411 = rbit_2_1.ram_58_0.m0_s 
* net 4412 = rbit_2_1.ram_58_0.m1_s 
* net 4413 = rbit_2_1.ram_57_1.m0_s 
* net 4414 = rbit_2_1.ram_57_1.m1_s 
* net 4415 = rbit_2_1.ram_57_0.m0_s 
* net 4416 = rbit_2_1.ram_57_0.m1_s 
* net 4417 = rbit_2_1.ram_56_1.m0_s 
* net 4418 = rbit_2_1.ram_56_1.m1_s 
* net 4419 = rbit_2_1.ram_56_0.m0_s 
* net 4420 = rbit_2_1.ram_56_0.m1_s 
* net 4421 = rbit_2_1.ram_55_1.m0_s 
* net 4422 = rbit_2_1.ram_55_1.m1_s 
* net 4423 = rbit_2_1.ram_55_0.m0_s 
* net 4424 = rbit_2_1.ram_55_0.m1_s 
* net 4425 = rbit_2_1.ram_54_1.m0_s 
* net 4426 = rbit_2_1.ram_54_1.m1_s 
* net 4427 = rbit_2_1.ram_54_0.m0_s 
* net 4428 = rbit_2_1.ram_54_0.m1_s 
* net 4429 = rbit_2_1.ram_53_1.m0_s 
* net 4430 = rbit_2_1.ram_53_1.m1_s 
* net 4431 = rbit_2_1.ram_53_0.m0_s 
* net 4432 = rbit_2_1.ram_53_0.m1_s 
* net 4433 = rbit_2_1.ram_52_1.m0_s 
* net 4434 = rbit_2_1.ram_52_1.m1_s 
* net 4435 = rbit_2_1.ram_52_0.m0_s 
* net 4436 = rbit_2_1.ram_52_0.m1_s 
* net 4437 = rbit_2_1.ram_51_1.m0_s 
* net 4438 = rbit_2_1.ram_51_1.m1_s 
* net 4439 = rbit_2_1.ram_51_0.m0_s 
* net 4440 = rbit_2_1.ram_51_0.m1_s 
* net 4441 = rbit_2_1.ram_50_1.m0_s 
* net 4442 = rbit_2_1.ram_50_1.m1_s 
* net 4443 = rbit_2_1.ram_50_0.m0_s 
* net 4444 = rbit_2_1.ram_50_0.m1_s 
* net 4445 = rbit_2_1.ram_49_1.m0_s 
* net 4446 = rbit_2_1.ram_49_1.m1_s 
* net 4447 = rbit_2_1.ram_49_0.m0_s 
* net 4448 = rbit_2_1.ram_49_0.m1_s 
* net 4449 = rbit_2_1.ram_48_1.m0_s 
* net 4450 = rbit_2_1.ram_48_1.m1_s 
* net 4451 = rbit_2_1.ram_48_0.m0_s 
* net 4452 = rbit_2_1.ram_48_0.m1_s 
* net 4453 = rbit_2_1.ram_47_1.m0_s 
* net 4454 = rbit_2_1.ram_47_1.m1_s 
* net 4455 = rbit_2_1.ram_47_0.m0_s 
* net 4456 = rbit_2_1.ram_47_0.m1_s 
* net 4457 = rbit_2_1.ram_46_1.m0_s 
* net 4458 = rbit_2_1.ram_46_1.m1_s 
* net 4459 = rbit_2_1.ram_46_0.m0_s 
* net 4460 = rbit_2_1.ram_46_0.m1_s 
* net 4461 = rbit_2_1.ram_45_1.m0_s 
* net 4462 = rbit_2_1.ram_45_1.m1_s 
* net 4463 = rbit_2_1.ram_45_0.m0_s 
* net 4464 = rbit_2_1.ram_45_0.m1_s 
* net 4465 = rbit_2_1.ram_44_1.m0_s 
* net 4466 = rbit_2_1.ram_44_1.m1_s 
* net 4467 = rbit_2_1.ram_44_0.m0_s 
* net 4468 = rbit_2_1.ram_44_0.m1_s 
* net 4469 = rbit_2_1.ram_43_1.m0_s 
* net 4470 = rbit_2_1.ram_43_1.m1_s 
* net 4471 = rbit_2_1.ram_43_0.m0_s 
* net 4472 = rbit_2_1.ram_43_0.m1_s 
* net 4473 = rbit_2_1.ram_42_1.m0_s 
* net 4474 = rbit_2_1.ram_42_1.m1_s 
* net 4475 = rbit_2_1.ram_42_0.m0_s 
* net 4476 = rbit_2_1.ram_42_0.m1_s 
* net 4477 = rbit_2_1.ram_41_1.m0_s 
* net 4478 = rbit_2_1.ram_41_1.m1_s 
* net 4479 = rbit_2_1.ram_41_0.m0_s 
* net 4480 = rbit_2_1.ram_41_0.m1_s 
* net 4481 = rbit_2_1.ram_40_1.m0_s 
* net 4482 = rbit_2_1.ram_40_1.m1_s 
* net 4483 = rbit_2_1.ram_40_0.m0_s 
* net 4484 = rbit_2_1.ram_40_0.m1_s 
* net 4485 = rbit_2_1.ram_39_1.m0_s 
* net 4486 = rbit_2_1.ram_39_1.m1_s 
* net 4487 = rbit_2_1.ram_39_0.m0_s 
* net 4488 = rbit_2_1.ram_39_0.m1_s 
* net 4489 = rbit_2_1.ram_38_1.m0_s 
* net 4490 = rbit_2_1.ram_38_1.m1_s 
* net 4491 = rbit_2_1.ram_38_0.m0_s 
* net 4492 = rbit_2_1.ram_38_0.m1_s 
* net 4493 = rbit_2_1.ram_37_1.m0_s 
* net 4494 = rbit_2_1.ram_37_1.m1_s 
* net 4495 = rbit_2_1.ram_37_0.m0_s 
* net 4496 = rbit_2_1.ram_37_0.m1_s 
* net 4497 = rbit_2_1.ram_36_1.m0_s 
* net 4498 = rbit_2_1.ram_36_1.m1_s 
* net 4499 = rbit_2_1.ram_36_0.m0_s 
* net 4500 = rbit_2_1.ram_36_0.m1_s 
* net 4501 = rbit_2_1.ram_35_1.m0_s 
* net 4502 = rbit_2_1.ram_35_1.m1_s 
* net 4503 = rbit_2_1.ram_35_0.m0_s 
* net 4504 = rbit_2_1.ram_35_0.m1_s 
* net 4505 = rbit_2_1.ram_34_1.m0_s 
* net 4506 = rbit_2_1.ram_34_1.m1_s 
* net 4507 = rbit_2_1.ram_34_0.m0_s 
* net 4508 = rbit_2_1.ram_34_0.m1_s 
* net 4509 = rbit_2_1.ram_33_1.m0_s 
* net 4510 = rbit_2_1.ram_33_1.m1_s 
* net 4511 = rbit_2_1.ram_33_0.m0_s 
* net 4512 = rbit_2_1.ram_33_0.m1_s 
* net 4513 = rbit_2_1.ram_32_1.m0_s 
* net 4514 = rbit_2_1.ram_32_1.m1_s 
* net 4515 = rbit_2_1.ram_32_0.m0_s 
* net 4516 = rbit_2_1.ram_32_0.m1_s 
* net 4517 = rbit_2_1.ram_31_1.m0_s 
* net 4518 = rbit_2_1.ram_31_1.m1_s 
* net 4519 = rbit_2_1.ram_31_0.m0_s 
* net 4520 = rbit_2_1.ram_31_0.m1_s 
* net 4521 = rbit_2_1.ram_30_1.m0_s 
* net 4522 = rbit_2_1.ram_30_1.m1_s 
* net 4523 = rbit_2_1.ram_30_0.m0_s 
* net 4524 = rbit_2_1.ram_30_0.m1_s 
* net 4525 = rbit_2_1.ram_29_1.m0_s 
* net 4526 = rbit_2_1.ram_29_1.m1_s 
* net 4527 = rbit_2_1.ram_29_0.m0_s 
* net 4528 = rbit_2_1.ram_29_0.m1_s 
* net 4529 = rbit_2_1.ram_28_1.m0_s 
* net 4530 = rbit_2_1.ram_28_1.m1_s 
* net 4531 = rbit_2_1.ram_28_0.m0_s 
* net 4532 = rbit_2_1.ram_28_0.m1_s 
* net 4533 = rbit_2_1.ram_27_1.m0_s 
* net 4534 = rbit_2_1.ram_27_1.m1_s 
* net 4535 = rbit_2_1.ram_27_0.m0_s 
* net 4536 = rbit_2_1.ram_27_0.m1_s 
* net 4537 = rbit_2_1.ram_26_1.m0_s 
* net 4538 = rbit_2_1.ram_26_1.m1_s 
* net 4539 = rbit_2_1.ram_26_0.m0_s 
* net 4540 = rbit_2_1.ram_26_0.m1_s 
* net 4541 = rbit_2_1.ram_25_1.m0_s 
* net 4542 = rbit_2_1.ram_25_1.m1_s 
* net 4543 = rbit_2_1.ram_25_0.m0_s 
* net 4544 = rbit_2_1.ram_25_0.m1_s 
* net 4545 = rbit_2_1.ram_24_1.m0_s 
* net 4546 = rbit_2_1.ram_24_1.m1_s 
* net 4547 = rbit_2_1.ram_24_0.m0_s 
* net 4548 = rbit_2_1.ram_24_0.m1_s 
* net 4549 = rbit_2_1.ram_23_1.m0_s 
* net 4550 = rbit_2_1.ram_23_1.m1_s 
* net 4551 = rbit_2_1.ram_23_0.m0_s 
* net 4552 = rbit_2_1.ram_23_0.m1_s 
* net 4553 = rbit_2_1.ram_22_1.m0_s 
* net 4554 = rbit_2_1.ram_22_1.m1_s 
* net 4555 = rbit_2_1.ram_22_0.m0_s 
* net 4556 = rbit_2_1.ram_22_0.m1_s 
* net 4557 = rbit_2_1.ram_21_1.m0_s 
* net 4558 = rbit_2_1.ram_21_1.m1_s 
* net 4559 = rbit_2_1.ram_21_0.m0_s 
* net 4560 = rbit_2_1.ram_21_0.m1_s 
* net 4561 = rbit_2_1.ram_20_1.m0_s 
* net 4562 = rbit_2_1.ram_20_1.m1_s 
* net 4563 = rbit_2_1.ram_20_0.m0_s 
* net 4564 = rbit_2_1.ram_20_0.m1_s 
* net 4565 = rbit_2_1.ram_19_1.m0_s 
* net 4566 = rbit_2_1.ram_19_1.m1_s 
* net 4567 = rbit_2_1.ram_19_0.m0_s 
* net 4568 = rbit_2_1.ram_19_0.m1_s 
* net 4569 = rbit_2_1.ram_18_1.m0_s 
* net 4570 = rbit_2_1.ram_18_1.m1_s 
* net 4571 = rbit_2_1.ram_18_0.m0_s 
* net 4572 = rbit_2_1.ram_18_0.m1_s 
* net 4573 = rbit_2_1.ram_17_1.m0_s 
* net 4574 = rbit_2_1.ram_17_1.m1_s 
* net 4575 = rbit_2_1.ram_17_0.m0_s 
* net 4576 = rbit_2_1.ram_17_0.m1_s 
* net 4577 = rbit_2_1.ram_16_1.m0_s 
* net 4578 = rbit_2_1.ram_16_1.m1_s 
* net 4579 = rbit_2_1.ram_16_0.m0_s 
* net 4580 = rbit_2_1.ram_16_0.m1_s 
* net 4581 = rbit_2_1.ram_15_1.m0_s 
* net 4582 = rbit_2_1.ram_15_1.m1_s 
* net 4583 = rbit_2_1.ram_15_0.m0_s 
* net 4584 = rbit_2_1.ram_15_0.m1_s 
* net 4585 = rbit_2_1.ram_14_1.m0_s 
* net 4586 = rbit_2_1.ram_14_1.m1_s 
* net 4587 = rbit_2_1.ram_14_0.m0_s 
* net 4588 = rbit_2_1.ram_14_0.m1_s 
* net 4589 = rbit_2_1.ram_13_1.m0_s 
* net 4590 = rbit_2_1.ram_13_1.m1_s 
* net 4591 = rbit_2_1.ram_13_0.m0_s 
* net 4592 = rbit_2_1.ram_13_0.m1_s 
* net 4593 = rbit_2_1.ram_12_1.m0_s 
* net 4594 = rbit_2_1.ram_12_1.m1_s 
* net 4595 = rbit_2_1.ram_12_0.m0_s 
* net 4596 = rbit_2_1.ram_12_0.m1_s 
* net 4597 = rbit_2_1.ram_11_1.m0_s 
* net 4598 = rbit_2_1.ram_11_1.m1_s 
* net 4599 = rbit_2_1.ram_11_0.m0_s 
* net 4600 = rbit_2_1.ram_11_0.m1_s 
* net 4601 = rbit_2_1.ram_10_1.m0_s 
* net 4602 = rbit_2_1.ram_10_1.m1_s 
* net 4603 = rbit_2_1.ram_10_0.m0_s 
* net 4604 = rbit_2_1.ram_10_0.m1_s 
* net 4605 = rbit_2_1.ram_9_1.m0_s 
* net 4606 = rbit_2_1.ram_9_1.m1_s 
* net 4607 = rbit_2_1.ram_9_0.m0_s 
* net 4608 = rbit_2_1.ram_9_0.m1_s 
* net 4609 = rbit_2_1.ram_8_1.m0_s 
* net 4610 = rbit_2_1.ram_8_1.m1_s 
* net 4611 = rbit_2_1.ram_8_0.m0_s 
* net 4612 = rbit_2_1.ram_8_0.m1_s 
* net 4613 = rbit_2_1.ram_7_1.m0_s 
* net 4614 = rbit_2_1.ram_7_1.m1_s 
* net 4615 = rbit_2_1.ram_7_0.m0_s 
* net 4616 = rbit_2_1.ram_7_0.m1_s 
* net 4617 = rbit_2_1.ram_6_1.m0_s 
* net 4618 = rbit_2_1.ram_6_1.m1_s 
* net 4619 = rbit_2_1.ram_6_0.m0_s 
* net 4620 = rbit_2_1.ram_6_0.m1_s 
* net 4621 = rbit_2_1.ram_5_1.m0_s 
* net 4622 = rbit_2_1.ram_5_1.m1_s 
* net 4623 = rbit_2_1.ram_5_0.m0_s 
* net 4624 = rbit_2_1.ram_5_0.m1_s 
* net 4625 = rbit_2_1.ram_4_1.m0_s 
* net 4626 = rbit_2_1.ram_4_1.m1_s 
* net 4627 = rbit_2_1.ram_4_0.m0_s 
* net 4628 = rbit_2_1.ram_4_0.m1_s 
* net 4629 = rbit_2_1.ram_3_1.m0_s 
* net 4630 = rbit_2_1.ram_3_1.m1_s 
* net 4631 = rbit_2_1.ram_3_0.m0_s 
* net 4632 = rbit_2_1.ram_3_0.m1_s 
* net 4633 = rbit_2_1.ram_2_1.m0_s 
* net 4634 = rbit_2_1.ram_2_1.m1_s 
* net 4635 = rbit_2_1.ram_2_0.m0_s 
* net 4636 = rbit_2_1.ram_2_0.m1_s 
* net 4637 = rbit_2_1.ram_1_1.m0_s 
* net 4638 = rbit_2_1.ram_1_1.m1_s 
* net 4639 = rbit_2_1.ram_1_0.m0_s 
* net 4640 = rbit_2_1.ram_1_0.m1_s 
* net 4641 = rbit_2_1.ram_0_1.m0_s 
* net 4642 = rbit_2_1.ram_0_1.m1_s 
* net 4643 = rbit_2_1.ram_0_0.m0_s 
* net 4644 = rbit_2_1.ram_0_0.m1_s 
* net 4645 = mbk_sig150 
* net 4646 = mbk_sig129 
* net 4647 = mbk_sig173 
* net 4648 = mbk_sig128 
* net 4649 = mbk_sig190 
* net 4650 = mbk_sig52 
* net 4651 = mbk_sig53 
* net 4652 = mbk_sig78 
* net 4653 = mbk_sig104 
* net 4654 = mbk_sig96 
* net 4655 = mbk_sig88 
* net 4656 = rbit_3_1.ram_127_1.m0_s 
* net 4657 = rbit_3_1.ram_127_1.m1_s 
* net 4658 = rbit_3_1.ram_127_0.m0_s 
* net 4659 = rbit_3_1.ram_127_0.m1_s 
* net 4660 = rbit_3_1.ram_126_1.m0_s 
* net 4661 = rbit_3_1.ram_126_1.m1_s 
* net 4662 = rbit_3_1.ram_126_0.m0_s 
* net 4663 = rbit_3_1.ram_126_0.m1_s 
* net 4664 = rbit_3_1.ram_125_1.m0_s 
* net 4665 = rbit_3_1.ram_125_1.m1_s 
* net 4666 = rbit_3_1.ram_125_0.m0_s 
* net 4667 = rbit_3_1.ram_125_0.m1_s 
* net 4668 = rbit_3_1.ram_124_1.m0_s 
* net 4669 = rbit_3_1.ram_124_1.m1_s 
* net 4670 = rbit_3_1.ram_124_0.m0_s 
* net 4671 = rbit_3_1.ram_124_0.m1_s 
* net 4672 = rbit_3_1.ram_123_1.m0_s 
* net 4673 = rbit_3_1.ram_123_1.m1_s 
* net 4674 = rbit_3_1.ram_123_0.m0_s 
* net 4675 = rbit_3_1.ram_123_0.m1_s 
* net 4676 = rbit_3_1.ram_122_1.m0_s 
* net 4677 = rbit_3_1.ram_122_1.m1_s 
* net 4678 = rbit_3_1.ram_122_0.m0_s 
* net 4679 = rbit_3_1.ram_122_0.m1_s 
* net 4680 = rbit_3_1.ram_121_1.m0_s 
* net 4681 = rbit_3_1.ram_121_1.m1_s 
* net 4682 = rbit_3_1.ram_121_0.m0_s 
* net 4683 = rbit_3_1.ram_121_0.m1_s 
* net 4684 = rbit_3_1.ram_120_1.m0_s 
* net 4685 = rbit_3_1.ram_120_1.m1_s 
* net 4686 = rbit_3_1.ram_120_0.m0_s 
* net 4687 = rbit_3_1.ram_120_0.m1_s 
* net 4688 = rbit_3_1.ram_119_1.m0_s 
* net 4689 = rbit_3_1.ram_119_1.m1_s 
* net 4690 = rbit_3_1.ram_119_0.m0_s 
* net 4691 = rbit_3_1.ram_119_0.m1_s 
* net 4692 = rbit_3_1.ram_118_1.m0_s 
* net 4693 = rbit_3_1.ram_118_1.m1_s 
* net 4694 = rbit_3_1.ram_118_0.m0_s 
* net 4695 = rbit_3_1.ram_118_0.m1_s 
* net 4696 = rbit_3_1.ram_117_1.m0_s 
* net 4697 = rbit_3_1.ram_117_1.m1_s 
* net 4698 = rbit_3_1.ram_117_0.m0_s 
* net 4699 = rbit_3_1.ram_117_0.m1_s 
* net 4700 = rbit_3_1.ram_116_1.m0_s 
* net 4701 = rbit_3_1.ram_116_1.m1_s 
* net 4702 = rbit_3_1.ram_116_0.m0_s 
* net 4703 = rbit_3_1.ram_116_0.m1_s 
* net 4704 = rbit_3_1.ram_115_1.m0_s 
* net 4705 = rbit_3_1.ram_115_1.m1_s 
* net 4706 = rbit_3_1.ram_115_0.m0_s 
* net 4707 = rbit_3_1.ram_115_0.m1_s 
* net 4708 = rbit_3_1.ram_114_1.m0_s 
* net 4709 = rbit_3_1.ram_114_1.m1_s 
* net 4710 = rbit_3_1.ram_114_0.m0_s 
* net 4711 = rbit_3_1.ram_114_0.m1_s 
* net 4712 = rbit_3_1.ram_113_1.m0_s 
* net 4713 = rbit_3_1.ram_113_1.m1_s 
* net 4714 = rbit_3_1.ram_113_0.m0_s 
* net 4715 = rbit_3_1.ram_113_0.m1_s 
* net 4716 = rbit_3_1.ram_112_1.m0_s 
* net 4717 = rbit_3_1.ram_112_1.m1_s 
* net 4718 = rbit_3_1.ram_112_0.m0_s 
* net 4719 = rbit_3_1.ram_112_0.m1_s 
* net 4720 = rbit_3_1.ram_111_1.m0_s 
* net 4721 = rbit_3_1.ram_111_1.m1_s 
* net 4722 = rbit_3_1.ram_111_0.m0_s 
* net 4723 = rbit_3_1.ram_111_0.m1_s 
* net 4724 = rbit_3_1.ram_110_1.m0_s 
* net 4725 = rbit_3_1.ram_110_1.m1_s 
* net 4726 = rbit_3_1.ram_110_0.m0_s 
* net 4727 = rbit_3_1.ram_110_0.m1_s 
* net 4728 = rbit_3_1.ram_109_1.m0_s 
* net 4729 = rbit_3_1.ram_109_1.m1_s 
* net 4730 = rbit_3_1.ram_109_0.m0_s 
* net 4731 = rbit_3_1.ram_109_0.m1_s 
* net 4732 = rbit_3_1.ram_108_1.m0_s 
* net 4733 = rbit_3_1.ram_108_1.m1_s 
* net 4734 = rbit_3_1.ram_108_0.m0_s 
* net 4735 = rbit_3_1.ram_108_0.m1_s 
* net 4736 = rbit_3_1.ram_107_1.m0_s 
* net 4737 = rbit_3_1.ram_107_1.m1_s 
* net 4738 = rbit_3_1.ram_107_0.m0_s 
* net 4739 = rbit_3_1.ram_107_0.m1_s 
* net 4740 = rbit_3_1.ram_106_1.m0_s 
* net 4741 = rbit_3_1.ram_106_1.m1_s 
* net 4742 = rbit_3_1.ram_106_0.m0_s 
* net 4743 = rbit_3_1.ram_106_0.m1_s 
* net 4744 = rbit_3_1.ram_105_1.m0_s 
* net 4745 = rbit_3_1.ram_105_1.m1_s 
* net 4746 = rbit_3_1.ram_105_0.m0_s 
* net 4747 = rbit_3_1.ram_105_0.m1_s 
* net 4748 = rbit_3_1.ram_104_1.m0_s 
* net 4749 = rbit_3_1.ram_104_1.m1_s 
* net 4750 = rbit_3_1.ram_104_0.m0_s 
* net 4751 = rbit_3_1.ram_104_0.m1_s 
* net 4752 = rbit_3_1.ram_103_1.m0_s 
* net 4753 = rbit_3_1.ram_103_1.m1_s 
* net 4754 = rbit_3_1.ram_103_0.m0_s 
* net 4755 = rbit_3_1.ram_103_0.m1_s 
* net 4756 = rbit_3_1.ram_102_1.m0_s 
* net 4757 = rbit_3_1.ram_102_1.m1_s 
* net 4758 = rbit_3_1.ram_102_0.m0_s 
* net 4759 = rbit_3_1.ram_102_0.m1_s 
* net 4760 = rbit_3_1.ram_101_1.m0_s 
* net 4761 = rbit_3_1.ram_101_1.m1_s 
* net 4762 = rbit_3_1.ram_101_0.m0_s 
* net 4763 = rbit_3_1.ram_101_0.m1_s 
* net 4764 = rbit_3_1.ram_100_1.m0_s 
* net 4765 = rbit_3_1.ram_100_1.m1_s 
* net 4766 = rbit_3_1.ram_100_0.m0_s 
* net 4767 = rbit_3_1.ram_100_0.m1_s 
* net 4768 = rbit_3_1.ram_99_1.m0_s 
* net 4769 = rbit_3_1.ram_99_1.m1_s 
* net 4770 = rbit_3_1.ram_99_0.m0_s 
* net 4771 = rbit_3_1.ram_99_0.m1_s 
* net 4772 = rbit_3_1.ram_98_1.m0_s 
* net 4773 = rbit_3_1.ram_98_1.m1_s 
* net 4774 = rbit_3_1.ram_98_0.m0_s 
* net 4775 = rbit_3_1.ram_98_0.m1_s 
* net 4776 = rbit_3_1.ram_97_1.m0_s 
* net 4777 = rbit_3_1.ram_97_1.m1_s 
* net 4778 = rbit_3_1.ram_97_0.m0_s 
* net 4779 = rbit_3_1.ram_97_0.m1_s 
* net 4780 = rbit_3_1.ram_96_1.m0_s 
* net 4781 = rbit_3_1.ram_96_1.m1_s 
* net 4782 = rbit_3_1.ram_96_0.m0_s 
* net 4783 = rbit_3_1.ram_96_0.m1_s 
* net 4784 = rbit_3_1.ram_95_1.m0_s 
* net 4785 = rbit_3_1.ram_95_1.m1_s 
* net 4786 = rbit_3_1.ram_95_0.m0_s 
* net 4787 = rbit_3_1.ram_95_0.m1_s 
* net 4788 = rbit_3_1.ram_94_1.m0_s 
* net 4789 = rbit_3_1.ram_94_1.m1_s 
* net 4790 = rbit_3_1.ram_94_0.m0_s 
* net 4791 = rbit_3_1.ram_94_0.m1_s 
* net 4792 = rbit_3_1.ram_93_1.m0_s 
* net 4793 = rbit_3_1.ram_93_1.m1_s 
* net 4794 = rbit_3_1.ram_93_0.m0_s 
* net 4795 = rbit_3_1.ram_93_0.m1_s 
* net 4796 = rbit_3_1.ram_92_1.m0_s 
* net 4797 = rbit_3_1.ram_92_1.m1_s 
* net 4798 = rbit_3_1.ram_92_0.m0_s 
* net 4799 = rbit_3_1.ram_92_0.m1_s 
* net 4800 = rbit_3_1.ram_91_1.m0_s 
* net 4801 = rbit_3_1.ram_91_1.m1_s 
* net 4802 = rbit_3_1.ram_91_0.m0_s 
* net 4803 = rbit_3_1.ram_91_0.m1_s 
* net 4804 = rbit_3_1.ram_90_1.m0_s 
* net 4805 = rbit_3_1.ram_90_1.m1_s 
* net 4806 = rbit_3_1.ram_90_0.m0_s 
* net 4807 = rbit_3_1.ram_90_0.m1_s 
* net 4808 = rbit_3_1.ram_89_1.m0_s 
* net 4809 = rbit_3_1.ram_89_1.m1_s 
* net 4810 = rbit_3_1.ram_89_0.m0_s 
* net 4811 = rbit_3_1.ram_89_0.m1_s 
* net 4812 = rbit_3_1.ram_88_1.m0_s 
* net 4813 = rbit_3_1.ram_88_1.m1_s 
* net 4814 = rbit_3_1.ram_88_0.m0_s 
* net 4815 = rbit_3_1.ram_88_0.m1_s 
* net 4816 = rbit_3_1.ram_87_1.m0_s 
* net 4817 = rbit_3_1.ram_87_1.m1_s 
* net 4818 = rbit_3_1.ram_87_0.m0_s 
* net 4819 = rbit_3_1.ram_87_0.m1_s 
* net 4820 = rbit_3_1.ram_86_1.m0_s 
* net 4821 = rbit_3_1.ram_86_1.m1_s 
* net 4822 = rbit_3_1.ram_86_0.m0_s 
* net 4823 = rbit_3_1.ram_86_0.m1_s 
* net 4824 = rbit_3_1.ram_85_1.m0_s 
* net 4825 = rbit_3_1.ram_85_1.m1_s 
* net 4826 = rbit_3_1.ram_85_0.m0_s 
* net 4827 = rbit_3_1.ram_85_0.m1_s 
* net 4828 = rbit_3_1.ram_84_1.m0_s 
* net 4829 = rbit_3_1.ram_84_1.m1_s 
* net 4830 = rbit_3_1.ram_84_0.m0_s 
* net 4831 = rbit_3_1.ram_84_0.m1_s 
* net 4832 = rbit_3_1.ram_83_1.m0_s 
* net 4833 = rbit_3_1.ram_83_1.m1_s 
* net 4834 = rbit_3_1.ram_83_0.m0_s 
* net 4835 = rbit_3_1.ram_83_0.m1_s 
* net 4836 = rbit_3_1.ram_82_1.m0_s 
* net 4837 = rbit_3_1.ram_82_1.m1_s 
* net 4838 = rbit_3_1.ram_82_0.m0_s 
* net 4839 = rbit_3_1.ram_82_0.m1_s 
* net 4840 = rbit_3_1.ram_81_1.m0_s 
* net 4841 = rbit_3_1.ram_81_1.m1_s 
* net 4842 = rbit_3_1.ram_81_0.m0_s 
* net 4843 = rbit_3_1.ram_81_0.m1_s 
* net 4844 = rbit_3_1.ram_80_1.m0_s 
* net 4845 = rbit_3_1.ram_80_1.m1_s 
* net 4846 = rbit_3_1.ram_80_0.m0_s 
* net 4847 = rbit_3_1.ram_80_0.m1_s 
* net 4848 = rbit_3_1.ram_79_1.m0_s 
* net 4849 = rbit_3_1.ram_79_1.m1_s 
* net 4850 = rbit_3_1.ram_79_0.m0_s 
* net 4851 = rbit_3_1.ram_79_0.m1_s 
* net 4852 = rbit_3_1.ram_78_1.m0_s 
* net 4853 = rbit_3_1.ram_78_1.m1_s 
* net 4854 = rbit_3_1.ram_78_0.m0_s 
* net 4855 = rbit_3_1.ram_78_0.m1_s 
* net 4856 = rbit_3_1.ram_77_1.m0_s 
* net 4857 = rbit_3_1.ram_77_1.m1_s 
* net 4858 = rbit_3_1.ram_77_0.m0_s 
* net 4859 = rbit_3_1.ram_77_0.m1_s 
* net 4860 = rbit_3_1.ram_76_1.m0_s 
* net 4861 = rbit_3_1.ram_76_1.m1_s 
* net 4862 = rbit_3_1.ram_76_0.m0_s 
* net 4863 = rbit_3_1.ram_76_0.m1_s 
* net 4864 = rbit_3_1.ram_75_1.m0_s 
* net 4865 = rbit_3_1.ram_75_1.m1_s 
* net 4866 = rbit_3_1.ram_75_0.m0_s 
* net 4867 = rbit_3_1.ram_75_0.m1_s 
* net 4868 = rbit_3_1.ram_74_1.m0_s 
* net 4869 = rbit_3_1.ram_74_1.m1_s 
* net 4870 = rbit_3_1.ram_74_0.m0_s 
* net 4871 = rbit_3_1.ram_74_0.m1_s 
* net 4872 = rbit_3_1.ram_73_1.m0_s 
* net 4873 = rbit_3_1.ram_73_1.m1_s 
* net 4874 = rbit_3_1.ram_73_0.m0_s 
* net 4875 = rbit_3_1.ram_73_0.m1_s 
* net 4876 = rbit_3_1.ram_72_1.m0_s 
* net 4877 = rbit_3_1.ram_72_1.m1_s 
* net 4878 = rbit_3_1.ram_72_0.m0_s 
* net 4879 = rbit_3_1.ram_72_0.m1_s 
* net 4880 = rbit_3_1.ram_71_1.m0_s 
* net 4881 = rbit_3_1.ram_71_1.m1_s 
* net 4882 = rbit_3_1.ram_71_0.m0_s 
* net 4883 = rbit_3_1.ram_71_0.m1_s 
* net 4884 = rbit_3_1.ram_70_1.m0_s 
* net 4885 = rbit_3_1.ram_70_1.m1_s 
* net 4886 = rbit_3_1.ram_70_0.m0_s 
* net 4887 = rbit_3_1.ram_70_0.m1_s 
* net 4888 = rbit_3_1.ram_69_1.m0_s 
* net 4889 = rbit_3_1.ram_69_1.m1_s 
* net 4890 = rbit_3_1.ram_69_0.m0_s 
* net 4891 = rbit_3_1.ram_69_0.m1_s 
* net 4892 = rbit_3_1.ram_68_1.m0_s 
* net 4893 = rbit_3_1.ram_68_1.m1_s 
* net 4894 = rbit_3_1.ram_68_0.m0_s 
* net 4895 = rbit_3_1.ram_68_0.m1_s 
* net 4896 = rbit_3_1.ram_67_1.m0_s 
* net 4897 = rbit_3_1.ram_67_1.m1_s 
* net 4898 = rbit_3_1.ram_67_0.m0_s 
* net 4899 = rbit_3_1.ram_67_0.m1_s 
* net 4900 = rbit_3_1.ram_66_1.m0_s 
* net 4901 = rbit_3_1.ram_66_1.m1_s 
* net 4902 = rbit_3_1.ram_66_0.m0_s 
* net 4903 = rbit_3_1.ram_66_0.m1_s 
* net 4904 = rbit_3_1.ram_65_1.m0_s 
* net 4905 = rbit_3_1.ram_65_1.m1_s 
* net 4906 = rbit_3_1.ram_65_0.m0_s 
* net 4907 = rbit_3_1.ram_65_0.m1_s 
* net 4908 = rbit_3_1.ram_64_1.m0_s 
* net 4909 = rbit_3_1.ram_64_1.m1_s 
* net 4910 = rbit_3_1.ram_64_0.m0_s 
* net 4911 = rbit_3_1.ram_64_0.m1_s 
* net 4912 = rbit_3_1.ram_63_1.m0_s 
* net 4913 = rbit_3_1.ram_63_1.m1_s 
* net 4914 = rbit_3_1.ram_63_0.m0_s 
* net 4915 = rbit_3_1.ram_63_0.m1_s 
* net 4916 = rbit_3_1.ram_62_1.m0_s 
* net 4917 = rbit_3_1.ram_62_1.m1_s 
* net 4918 = rbit_3_1.ram_62_0.m0_s 
* net 4919 = rbit_3_1.ram_62_0.m1_s 
* net 4920 = rbit_3_1.ram_61_1.m0_s 
* net 4921 = rbit_3_1.ram_61_1.m1_s 
* net 4922 = rbit_3_1.ram_61_0.m0_s 
* net 4923 = rbit_3_1.ram_61_0.m1_s 
* net 4924 = rbit_3_1.ram_60_1.m0_s 
* net 4925 = rbit_3_1.ram_60_1.m1_s 
* net 4926 = rbit_3_1.ram_60_0.m0_s 
* net 4927 = rbit_3_1.ram_60_0.m1_s 
* net 4928 = rbit_3_1.ram_59_1.m0_s 
* net 4929 = rbit_3_1.ram_59_1.m1_s 
* net 4930 = rbit_3_1.ram_59_0.m0_s 
* net 4931 = rbit_3_1.ram_59_0.m1_s 
* net 4932 = rbit_3_1.ram_58_1.m0_s 
* net 4933 = rbit_3_1.ram_58_1.m1_s 
* net 4934 = rbit_3_1.ram_58_0.m0_s 
* net 4935 = rbit_3_1.ram_58_0.m1_s 
* net 4936 = rbit_3_1.ram_57_1.m0_s 
* net 4937 = rbit_3_1.ram_57_1.m1_s 
* net 4938 = rbit_3_1.ram_57_0.m0_s 
* net 4939 = rbit_3_1.ram_57_0.m1_s 
* net 4940 = rbit_3_1.ram_56_1.m0_s 
* net 4941 = rbit_3_1.ram_56_1.m1_s 
* net 4942 = rbit_3_1.ram_56_0.m0_s 
* net 4943 = rbit_3_1.ram_56_0.m1_s 
* net 4944 = rbit_3_1.ram_55_1.m0_s 
* net 4945 = rbit_3_1.ram_55_1.m1_s 
* net 4946 = rbit_3_1.ram_55_0.m0_s 
* net 4947 = rbit_3_1.ram_55_0.m1_s 
* net 4948 = rbit_3_1.ram_54_1.m0_s 
* net 4949 = rbit_3_1.ram_54_1.m1_s 
* net 4950 = rbit_3_1.ram_54_0.m0_s 
* net 4951 = rbit_3_1.ram_54_0.m1_s 
* net 4952 = rbit_3_1.ram_53_1.m0_s 
* net 4953 = rbit_3_1.ram_53_1.m1_s 
* net 4954 = rbit_3_1.ram_53_0.m0_s 
* net 4955 = rbit_3_1.ram_53_0.m1_s 
* net 4956 = rbit_3_1.ram_52_1.m0_s 
* net 4957 = rbit_3_1.ram_52_1.m1_s 
* net 4958 = rbit_3_1.ram_52_0.m0_s 
* net 4959 = rbit_3_1.ram_52_0.m1_s 
* net 4960 = rbit_3_1.ram_51_1.m0_s 
* net 4961 = rbit_3_1.ram_51_1.m1_s 
* net 4962 = rbit_3_1.ram_51_0.m0_s 
* net 4963 = rbit_3_1.ram_51_0.m1_s 
* net 4964 = rbit_3_1.ram_50_1.m0_s 
* net 4965 = rbit_3_1.ram_50_1.m1_s 
* net 4966 = rbit_3_1.ram_50_0.m0_s 
* net 4967 = rbit_3_1.ram_50_0.m1_s 
* net 4968 = rbit_3_1.ram_49_1.m0_s 
* net 4969 = rbit_3_1.ram_49_1.m1_s 
* net 4970 = rbit_3_1.ram_49_0.m0_s 
* net 4971 = rbit_3_1.ram_49_0.m1_s 
* net 4972 = rbit_3_1.ram_48_1.m0_s 
* net 4973 = rbit_3_1.ram_48_1.m1_s 
* net 4974 = rbit_3_1.ram_48_0.m0_s 
* net 4975 = rbit_3_1.ram_48_0.m1_s 
* net 4976 = rbit_3_1.ram_47_1.m0_s 
* net 4977 = rbit_3_1.ram_47_1.m1_s 
* net 4978 = rbit_3_1.ram_47_0.m0_s 
* net 4979 = rbit_3_1.ram_47_0.m1_s 
* net 4980 = rbit_3_1.ram_46_1.m0_s 
* net 4981 = rbit_3_1.ram_46_1.m1_s 
* net 4982 = rbit_3_1.ram_46_0.m0_s 
* net 4983 = rbit_3_1.ram_46_0.m1_s 
* net 4984 = rbit_3_1.ram_45_1.m0_s 
* net 4985 = rbit_3_1.ram_45_1.m1_s 
* net 4986 = rbit_3_1.ram_45_0.m0_s 
* net 4987 = rbit_3_1.ram_45_0.m1_s 
* net 4988 = rbit_3_1.ram_44_1.m0_s 
* net 4989 = rbit_3_1.ram_44_1.m1_s 
* net 4990 = rbit_3_1.ram_44_0.m0_s 
* net 4991 = rbit_3_1.ram_44_0.m1_s 
* net 4992 = rbit_3_1.ram_43_1.m0_s 
* net 4993 = rbit_3_1.ram_43_1.m1_s 
* net 4994 = rbit_3_1.ram_43_0.m0_s 
* net 4995 = rbit_3_1.ram_43_0.m1_s 
* net 4996 = rbit_3_1.ram_42_1.m0_s 
* net 4997 = rbit_3_1.ram_42_1.m1_s 
* net 4998 = rbit_3_1.ram_42_0.m0_s 
* net 4999 = rbit_3_1.ram_42_0.m1_s 
* net 5000 = rbit_3_1.ram_41_1.m0_s 
* net 5001 = rbit_3_1.ram_41_1.m1_s 
* net 5002 = rbit_3_1.ram_41_0.m0_s 
* net 5003 = rbit_3_1.ram_41_0.m1_s 
* net 5004 = rbit_3_1.ram_40_1.m0_s 
* net 5005 = rbit_3_1.ram_40_1.m1_s 
* net 5006 = rbit_3_1.ram_40_0.m0_s 
* net 5007 = rbit_3_1.ram_40_0.m1_s 
* net 5008 = rbit_3_1.ram_39_1.m0_s 
* net 5009 = rbit_3_1.ram_39_1.m1_s 
* net 5010 = rbit_3_1.ram_39_0.m0_s 
* net 5011 = rbit_3_1.ram_39_0.m1_s 
* net 5012 = rbit_3_1.ram_38_1.m0_s 
* net 5013 = rbit_3_1.ram_38_1.m1_s 
* net 5014 = rbit_3_1.ram_38_0.m0_s 
* net 5015 = rbit_3_1.ram_38_0.m1_s 
* net 5016 = rbit_3_1.ram_37_1.m0_s 
* net 5017 = rbit_3_1.ram_37_1.m1_s 
* net 5018 = rbit_3_1.ram_37_0.m0_s 
* net 5019 = rbit_3_1.ram_37_0.m1_s 
* net 5020 = rbit_3_1.ram_36_1.m0_s 
* net 5021 = rbit_3_1.ram_36_1.m1_s 
* net 5022 = rbit_3_1.ram_36_0.m0_s 
* net 5023 = rbit_3_1.ram_36_0.m1_s 
* net 5024 = rbit_3_1.ram_35_1.m0_s 
* net 5025 = rbit_3_1.ram_35_1.m1_s 
* net 5026 = rbit_3_1.ram_35_0.m0_s 
* net 5027 = rbit_3_1.ram_35_0.m1_s 
* net 5028 = rbit_3_1.ram_34_1.m0_s 
* net 5029 = rbit_3_1.ram_34_1.m1_s 
* net 5030 = rbit_3_1.ram_34_0.m0_s 
* net 5031 = rbit_3_1.ram_34_0.m1_s 
* net 5032 = rbit_3_1.ram_33_1.m0_s 
* net 5033 = rbit_3_1.ram_33_1.m1_s 
* net 5034 = rbit_3_1.ram_33_0.m0_s 
* net 5035 = rbit_3_1.ram_33_0.m1_s 
* net 5036 = rbit_3_1.ram_32_1.m0_s 
* net 5037 = rbit_3_1.ram_32_1.m1_s 
* net 5038 = rbit_3_1.ram_32_0.m0_s 
* net 5039 = rbit_3_1.ram_32_0.m1_s 
* net 5040 = rbit_3_1.ram_31_1.m0_s 
* net 5041 = rbit_3_1.ram_31_1.m1_s 
* net 5042 = rbit_3_1.ram_31_0.m0_s 
* net 5043 = rbit_3_1.ram_31_0.m1_s 
* net 5044 = rbit_3_1.ram_30_1.m0_s 
* net 5045 = rbit_3_1.ram_30_1.m1_s 
* net 5046 = rbit_3_1.ram_30_0.m0_s 
* net 5047 = rbit_3_1.ram_30_0.m1_s 
* net 5048 = rbit_3_1.ram_29_1.m0_s 
* net 5049 = rbit_3_1.ram_29_1.m1_s 
* net 5050 = rbit_3_1.ram_29_0.m0_s 
* net 5051 = rbit_3_1.ram_29_0.m1_s 
* net 5052 = rbit_3_1.ram_28_1.m0_s 
* net 5053 = rbit_3_1.ram_28_1.m1_s 
* net 5054 = rbit_3_1.ram_28_0.m0_s 
* net 5055 = rbit_3_1.ram_28_0.m1_s 
* net 5056 = rbit_3_1.ram_27_1.m0_s 
* net 5057 = rbit_3_1.ram_27_1.m1_s 
* net 5058 = rbit_3_1.ram_27_0.m0_s 
* net 5059 = rbit_3_1.ram_27_0.m1_s 
* net 5060 = rbit_3_1.ram_26_1.m0_s 
* net 5061 = rbit_3_1.ram_26_1.m1_s 
* net 5062 = rbit_3_1.ram_26_0.m0_s 
* net 5063 = rbit_3_1.ram_26_0.m1_s 
* net 5064 = rbit_3_1.ram_25_1.m0_s 
* net 5065 = rbit_3_1.ram_25_1.m1_s 
* net 5066 = rbit_3_1.ram_25_0.m0_s 
* net 5067 = rbit_3_1.ram_25_0.m1_s 
* net 5068 = rbit_3_1.ram_24_1.m0_s 
* net 5069 = rbit_3_1.ram_24_1.m1_s 
* net 5070 = rbit_3_1.ram_24_0.m0_s 
* net 5071 = rbit_3_1.ram_24_0.m1_s 
* net 5072 = rbit_3_1.ram_23_1.m0_s 
* net 5073 = rbit_3_1.ram_23_1.m1_s 
* net 5074 = rbit_3_1.ram_23_0.m0_s 
* net 5075 = rbit_3_1.ram_23_0.m1_s 
* net 5076 = rbit_3_1.ram_22_1.m0_s 
* net 5077 = rbit_3_1.ram_22_1.m1_s 
* net 5078 = rbit_3_1.ram_22_0.m0_s 
* net 5079 = rbit_3_1.ram_22_0.m1_s 
* net 5080 = rbit_3_1.ram_21_1.m0_s 
* net 5081 = rbit_3_1.ram_21_1.m1_s 
* net 5082 = rbit_3_1.ram_21_0.m0_s 
* net 5083 = rbit_3_1.ram_21_0.m1_s 
* net 5084 = rbit_3_1.ram_20_1.m0_s 
* net 5085 = rbit_3_1.ram_20_1.m1_s 
* net 5086 = rbit_3_1.ram_20_0.m0_s 
* net 5087 = rbit_3_1.ram_20_0.m1_s 
* net 5088 = rbit_3_1.ram_19_1.m0_s 
* net 5089 = rbit_3_1.ram_19_1.m1_s 
* net 5090 = rbit_3_1.ram_19_0.m0_s 
* net 5091 = rbit_3_1.ram_19_0.m1_s 
* net 5092 = rbit_3_1.ram_18_1.m0_s 
* net 5093 = rbit_3_1.ram_18_1.m1_s 
* net 5094 = rbit_3_1.ram_18_0.m0_s 
* net 5095 = rbit_3_1.ram_18_0.m1_s 
* net 5096 = rbit_3_1.ram_17_1.m0_s 
* net 5097 = rbit_3_1.ram_17_1.m1_s 
* net 5098 = rbit_3_1.ram_17_0.m0_s 
* net 5099 = rbit_3_1.ram_17_0.m1_s 
* net 5100 = rbit_3_1.ram_16_1.m0_s 
* net 5101 = rbit_3_1.ram_16_1.m1_s 
* net 5102 = rbit_3_1.ram_16_0.m0_s 
* net 5103 = rbit_3_1.ram_16_0.m1_s 
* net 5104 = rbit_3_1.ram_15_1.m0_s 
* net 5105 = rbit_3_1.ram_15_1.m1_s 
* net 5106 = rbit_3_1.ram_15_0.m0_s 
* net 5107 = rbit_3_1.ram_15_0.m1_s 
* net 5108 = rbit_3_1.ram_14_1.m0_s 
* net 5109 = rbit_3_1.ram_14_1.m1_s 
* net 5110 = rbit_3_1.ram_14_0.m0_s 
* net 5111 = rbit_3_1.ram_14_0.m1_s 
* net 5112 = rbit_3_1.ram_13_1.m0_s 
* net 5113 = rbit_3_1.ram_13_1.m1_s 
* net 5114 = rbit_3_1.ram_13_0.m0_s 
* net 5115 = rbit_3_1.ram_13_0.m1_s 
* net 5116 = rbit_3_1.ram_12_1.m0_s 
* net 5117 = rbit_3_1.ram_12_1.m1_s 
* net 5118 = rbit_3_1.ram_12_0.m0_s 
* net 5119 = rbit_3_1.ram_12_0.m1_s 
* net 5120 = rbit_3_1.ram_11_1.m0_s 
* net 5121 = rbit_3_1.ram_11_1.m1_s 
* net 5122 = rbit_3_1.ram_11_0.m0_s 
* net 5123 = rbit_3_1.ram_11_0.m1_s 
* net 5124 = rbit_3_1.ram_10_1.m0_s 
* net 5125 = rbit_3_1.ram_10_1.m1_s 
* net 5126 = rbit_3_1.ram_10_0.m0_s 
* net 5127 = rbit_3_1.ram_10_0.m1_s 
* net 5128 = rbit_3_1.ram_9_1.m0_s 
* net 5129 = rbit_3_1.ram_9_1.m1_s 
* net 5130 = rbit_3_1.ram_9_0.m0_s 
* net 5131 = rbit_3_1.ram_9_0.m1_s 
* net 5132 = rbit_3_1.ram_8_1.m0_s 
* net 5133 = rbit_3_1.ram_8_1.m1_s 
* net 5134 = rbit_3_1.ram_8_0.m0_s 
* net 5135 = rbit_3_1.ram_8_0.m1_s 
* net 5136 = rbit_3_1.ram_7_1.m0_s 
* net 5137 = rbit_3_1.ram_7_1.m1_s 
* net 5138 = rbit_3_1.ram_7_0.m0_s 
* net 5139 = rbit_3_1.ram_7_0.m1_s 
* net 5140 = rbit_3_1.ram_6_1.m0_s 
* net 5141 = rbit_3_1.ram_6_1.m1_s 
* net 5142 = rbit_3_1.ram_6_0.m0_s 
* net 5143 = rbit_3_1.ram_6_0.m1_s 
* net 5144 = rbit_3_1.ram_5_1.m0_s 
* net 5145 = rbit_3_1.ram_5_1.m1_s 
* net 5146 = rbit_3_1.ram_5_0.m0_s 
* net 5147 = rbit_3_1.ram_5_0.m1_s 
* net 5148 = rbit_3_1.ram_4_1.m0_s 
* net 5149 = rbit_3_1.ram_4_1.m1_s 
* net 5150 = rbit_3_1.ram_4_0.m0_s 
* net 5151 = rbit_3_1.ram_4_0.m1_s 
* net 5152 = rbit_3_1.ram_3_1.m0_s 
* net 5153 = rbit_3_1.ram_3_1.m1_s 
* net 5154 = rbit_3_1.ram_3_0.m0_s 
* net 5155 = rbit_3_1.ram_3_0.m1_s 
* net 5156 = rbit_3_1.ram_2_1.m0_s 
* net 5157 = rbit_3_1.ram_2_1.m1_s 
* net 5158 = rbit_3_1.ram_2_0.m0_s 
* net 5159 = rbit_3_1.ram_2_0.m1_s 
* net 5160 = rbit_3_1.ram_1_1.m0_s 
* net 5161 = rbit_3_1.ram_1_1.m1_s 
* net 5162 = rbit_3_1.ram_1_0.m0_s 
* net 5163 = rbit_3_1.ram_1_0.m1_s 
* net 5164 = rbit_3_1.ram_0_1.m0_s 
* net 5165 = rbit_3_1.ram_0_1.m1_s 
* net 5166 = rbit_3_1.ram_0_0.m0_s 
* net 5167 = rbit_3_1.ram_0_0.m1_s 
* net 5168 = mbk_sig153 
* net 5169 = mbk_sig131 
* net 5170 = mbk_sig176 
* net 5171 = mbk_sig130 
* net 5172 = mbk_sig191 
* net 5173 = mbk_sig59 
* net 5174 = mbk_sig57 
* net 5175 = mbk_sig79 
* net 5176 = mbk_sig81 
* net 5177 = mbk_sig105 
* net 5178 = mbk_sig97 
* net 5179 = mbk_sig39 
* net 5180 = mbk_sig89 
* net 5181 = write 
* net 5182 = vss 
* net 5183 = vdd 
* net 5184 = en 
* net 5185 = dout[7] 
* net 5186 = dout[6] 
* net 5187 = dout[5] 
* net 5188 = dout[4] 
* net 5189 = dout[3] 
* net 5190 = dout[2] 
* net 5191 = dout[1] 
* net 5192 = dout[0] 
* net 5193 = ck 
* net 5194 = adr[7] 
* net 5195 = adr[6] 
* net 5196 = adr[5] 
* net 5197 = adr[4] 
* net 5198 = adr[3] 
* net 5199 = adr[2] 
* net 5200 = adr[1] 
* net 5201 = adr[0] 
Mtr_00001 4 2529 2 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00002 4 2529 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00003 2 2529 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00004 3 2529 1 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00005 5183 2529 3 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00006 5183 2529 1 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00007 5182 437 436 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00008 437 436 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00009 4 2547 436 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00010 2 2547 437 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00011 5182 439 438 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00012 439 438 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00013 3 2547 438 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00014 1 2547 439 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00015 5182 441 440 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00016 441 440 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00017 4 2541 440 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00018 2 2541 441 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00019 5182 443 442 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00020 443 442 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00021 3 2541 442 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00022 1 2541 443 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00023 5182 445 444 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00024 445 444 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00025 4 2543 444 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00026 2 2543 445 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00027 5182 447 446 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00028 447 446 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00029 3 2543 446 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00030 1 2543 447 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00031 5182 449 448 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00032 449 448 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00033 4 2545 448 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00034 2 2545 449 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00035 5182 451 450 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00036 451 450 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00037 3 2545 450 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00038 1 2545 451 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00039 5182 453 452 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00040 453 452 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00041 4 2563 452 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00042 2 2563 453 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00043 5182 455 454 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00044 455 454 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00045 3 2563 454 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00046 1 2563 455 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00047 5182 457 456 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00048 457 456 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00049 4 2557 456 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00050 2 2557 457 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00051 5182 459 458 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00052 459 458 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00053 3 2557 458 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00054 1 2557 459 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00055 5182 461 460 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00056 461 460 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00057 4 2559 460 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00058 2 2559 461 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00059 5182 463 462 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00060 463 462 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00061 3 2559 462 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00062 1 2559 463 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00063 5182 465 464 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00064 465 464 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00065 4 2561 464 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00066 2 2561 465 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00067 5182 467 466 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00068 467 466 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00069 3 2561 466 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00070 1 2561 467 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00071 5182 469 468 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00072 469 468 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00073 4 2579 468 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00074 2 2579 469 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00075 5182 471 470 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00076 471 470 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00077 3 2579 470 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00078 1 2579 471 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00079 5182 473 472 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00080 473 472 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00081 4 2573 472 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00082 2 2573 473 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00083 5182 475 474 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00084 475 474 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00085 3 2573 474 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00086 1 2573 475 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00087 5182 477 476 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00088 477 476 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00089 4 2575 476 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00090 2 2575 477 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00091 5182 479 478 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00092 479 478 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00093 3 2575 478 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00094 1 2575 479 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00095 5182 481 480 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00096 481 480 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00097 4 2577 480 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00098 2 2577 481 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00099 5182 483 482 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00100 483 482 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00101 3 2577 482 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00102 1 2577 483 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00103 5182 485 484 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00104 485 484 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00105 4 2595 484 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00106 2 2595 485 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00107 5182 487 486 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00108 487 486 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00109 3 2595 486 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00110 1 2595 487 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00111 5182 489 488 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00112 489 488 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00113 4 2589 488 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00114 2 2589 489 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00115 5182 491 490 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00116 491 490 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00117 3 2589 490 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00118 1 2589 491 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00119 5182 493 492 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00120 493 492 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00121 4 2591 492 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00122 2 2591 493 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00123 5182 495 494 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00124 495 494 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00125 3 2591 494 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00126 1 2591 495 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00127 5182 497 496 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00128 497 496 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00129 4 2593 496 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00130 2 2593 497 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00131 5182 499 498 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00132 499 498 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00133 3 2593 498 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00134 1 2593 499 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00135 5182 501 500 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00136 501 500 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00137 4 2611 500 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00138 2 2611 501 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00139 5182 503 502 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00140 503 502 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00141 3 2611 502 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00142 1 2611 503 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00143 5182 505 504 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00144 505 504 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00145 4 2605 504 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00146 2 2605 505 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00147 5182 507 506 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00148 507 506 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00149 3 2605 506 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00150 1 2605 507 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00151 5182 509 508 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00152 509 508 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00153 4 2607 508 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00154 2 2607 509 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00155 5182 511 510 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00156 511 510 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00157 3 2607 510 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00158 1 2607 511 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00159 5182 513 512 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00160 513 512 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00161 4 2609 512 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00162 2 2609 513 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00163 5182 515 514 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00164 515 514 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00165 3 2609 514 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00166 1 2609 515 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00167 5182 517 516 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00168 517 516 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00169 4 2627 516 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00170 2 2627 517 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00171 5182 519 518 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00172 519 518 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00173 3 2627 518 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00174 1 2627 519 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00175 5182 521 520 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00176 521 520 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00177 4 2621 520 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00178 2 2621 521 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00179 5182 523 522 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00180 523 522 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00181 3 2621 522 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00182 1 2621 523 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00183 5182 525 524 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00184 525 524 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00185 4 2623 524 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00186 2 2623 525 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00187 5182 527 526 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00188 527 526 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00189 3 2623 526 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00190 1 2623 527 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00191 5182 529 528 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00192 529 528 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00193 4 2625 528 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00194 2 2625 529 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00195 5182 531 530 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00196 531 530 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00197 3 2625 530 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00198 1 2625 531 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00199 5182 533 532 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00200 533 532 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00201 4 2643 532 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00202 2 2643 533 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00203 5182 535 534 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00204 535 534 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00205 3 2643 534 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00206 1 2643 535 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00207 5182 537 536 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00208 537 536 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00209 4 2637 536 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00210 2 2637 537 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00211 5182 539 538 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00212 539 538 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00213 3 2637 538 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00214 1 2637 539 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00215 5182 541 540 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00216 541 540 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00217 4 2639 540 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00218 2 2639 541 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00219 5182 543 542 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00220 543 542 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00221 3 2639 542 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00222 1 2639 543 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00223 5182 545 544 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00224 545 544 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00225 4 2641 544 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00226 2 2641 545 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00227 5182 547 546 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00228 547 546 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00229 3 2641 546 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00230 1 2641 547 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00231 5182 549 548 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00232 549 548 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00233 4 2659 548 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00234 2 2659 549 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00235 5182 551 550 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00236 551 550 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00237 3 2659 550 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00238 1 2659 551 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00239 5182 553 552 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00240 553 552 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00241 4 2653 552 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00242 2 2653 553 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00243 5182 555 554 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00244 555 554 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00245 3 2653 554 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00246 1 2653 555 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00247 5182 557 556 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00248 557 556 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00249 4 2655 556 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00250 2 2655 557 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00251 5182 559 558 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00252 559 558 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00253 3 2655 558 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00254 1 2655 559 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00255 5182 561 560 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00256 561 560 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00257 4 2657 560 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00258 2 2657 561 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00259 5182 563 562 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00260 563 562 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00261 3 2657 562 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00262 1 2657 563 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00263 5182 565 564 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00264 565 564 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00265 4 2675 564 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00266 2 2675 565 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00267 5182 567 566 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00268 567 566 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00269 3 2675 566 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00270 1 2675 567 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00271 5182 569 568 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00272 569 568 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00273 4 2669 568 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00274 2 2669 569 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00275 5182 571 570 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00276 571 570 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00277 3 2669 570 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00278 1 2669 571 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00279 5182 573 572 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00280 573 572 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00281 4 2671 572 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00282 2 2671 573 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00283 5182 575 574 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00284 575 574 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00285 3 2671 574 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00286 1 2671 575 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00287 5182 577 576 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00288 577 576 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00289 4 2673 576 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00290 2 2673 577 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00291 5182 579 578 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00292 579 578 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00293 3 2673 578 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00294 1 2673 579 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00295 5182 581 580 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00296 581 580 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00297 4 2691 580 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00298 2 2691 581 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00299 5182 583 582 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00300 583 582 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00301 3 2691 582 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00302 1 2691 583 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00303 5182 585 584 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00304 585 584 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00305 4 2685 584 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00306 2 2685 585 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00307 5182 587 586 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00308 587 586 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00309 3 2685 586 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00310 1 2685 587 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00311 5182 589 588 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00312 589 588 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00313 4 2687 588 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00314 2 2687 589 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00315 5182 591 590 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00316 591 590 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00317 3 2687 590 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00318 1 2687 591 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00319 5182 593 592 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00320 593 592 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00321 4 2689 592 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00322 2 2689 593 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00323 5182 595 594 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00324 595 594 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00325 3 2689 594 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00326 1 2689 595 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00327 5182 597 596 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00328 597 596 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00329 4 2707 596 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00330 2 2707 597 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00331 5182 599 598 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00332 599 598 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00333 3 2707 598 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00334 1 2707 599 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00335 5182 601 600 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00336 601 600 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00337 4 2701 600 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00338 2 2701 601 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00339 5182 603 602 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00340 603 602 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00341 3 2701 602 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00342 1 2701 603 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00343 5182 605 604 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00344 605 604 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00345 4 2703 604 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00346 2 2703 605 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00347 5182 607 606 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00348 607 606 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00349 3 2703 606 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00350 1 2703 607 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00351 5182 609 608 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00352 609 608 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00353 4 2705 608 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00354 2 2705 609 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00355 5182 611 610 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00356 611 610 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00357 3 2705 610 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00358 1 2705 611 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00359 5182 613 612 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00360 613 612 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00361 4 2723 612 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00362 2 2723 613 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00363 5182 615 614 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00364 615 614 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00365 3 2723 614 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00366 1 2723 615 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00367 5182 617 616 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00368 617 616 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00369 4 2717 616 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00370 2 2717 617 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00371 5182 619 618 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00372 619 618 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00373 3 2717 618 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00374 1 2717 619 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00375 5182 621 620 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00376 621 620 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00377 4 2719 620 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00378 2 2719 621 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00379 5182 623 622 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00380 623 622 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00381 3 2719 622 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00382 1 2719 623 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00383 5182 625 624 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00384 625 624 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00385 4 2721 624 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00386 2 2721 625 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00387 5182 627 626 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00388 627 626 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00389 3 2721 626 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00390 1 2721 627 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00391 5182 629 628 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00392 629 628 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00393 4 2739 628 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00394 2 2739 629 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00395 5182 631 630 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00396 631 630 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00397 3 2739 630 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00398 1 2739 631 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00399 5182 633 632 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00400 633 632 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00401 4 2733 632 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00402 2 2733 633 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00403 5182 635 634 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00404 635 634 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00405 3 2733 634 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00406 1 2733 635 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00407 5182 637 636 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00408 637 636 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00409 4 2735 636 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00410 2 2735 637 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00411 5182 639 638 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00412 639 638 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00413 3 2735 638 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00414 1 2735 639 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00415 5182 641 640 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00416 641 640 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00417 4 2737 640 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00418 2 2737 641 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00419 5182 643 642 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00420 643 642 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00421 3 2737 642 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00422 1 2737 643 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00423 5182 645 644 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00424 645 644 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00425 4 2755 644 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00426 2 2755 645 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00427 5182 647 646 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00428 647 646 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00429 3 2755 646 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00430 1 2755 647 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00431 5182 649 648 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00432 649 648 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00433 4 2749 648 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00434 2 2749 649 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00435 5182 651 650 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00436 651 650 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00437 3 2749 650 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00438 1 2749 651 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00439 5182 653 652 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00440 653 652 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00441 4 2751 652 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00442 2 2751 653 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00443 5182 655 654 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00444 655 654 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00445 3 2751 654 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00446 1 2751 655 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00447 5182 657 656 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00448 657 656 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00449 4 2753 656 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00450 2 2753 657 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00451 5182 659 658 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00452 659 658 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00453 3 2753 658 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00454 1 2753 659 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00455 5182 661 660 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00456 661 660 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00457 4 2771 660 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00458 2 2771 661 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00459 5182 663 662 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00460 663 662 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00461 3 2771 662 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00462 1 2771 663 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00463 5182 665 664 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00464 665 664 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00465 4 2765 664 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00466 2 2765 665 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00467 5182 667 666 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00468 667 666 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00469 3 2765 666 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00470 1 2765 667 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00471 5182 669 668 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00472 669 668 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00473 4 2767 668 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00474 2 2767 669 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00475 5182 671 670 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00476 671 670 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00477 3 2767 670 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00478 1 2767 671 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00479 5182 673 672 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00480 673 672 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00481 4 2769 672 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00482 2 2769 673 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00483 5182 675 674 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00484 675 674 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00485 3 2769 674 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00486 1 2769 675 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00487 5182 677 676 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00488 677 676 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00489 4 2787 676 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00490 2 2787 677 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00491 5182 679 678 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00492 679 678 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00493 3 2787 678 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00494 1 2787 679 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00495 5182 681 680 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00496 681 680 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00497 4 2781 680 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00498 2 2781 681 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00499 5182 683 682 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00500 683 682 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00501 3 2781 682 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00502 1 2781 683 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00503 5182 685 684 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00504 685 684 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00505 4 2783 684 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00506 2 2783 685 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00507 5182 687 686 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00508 687 686 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00509 3 2783 686 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00510 1 2783 687 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00511 5182 689 688 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00512 689 688 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00513 4 2785 688 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00514 2 2785 689 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00515 5182 691 690 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00516 691 690 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00517 3 2785 690 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00518 1 2785 691 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00519 5182 693 692 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00520 693 692 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00521 4 2803 692 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00522 2 2803 693 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00523 5182 695 694 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00524 695 694 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00525 3 2803 694 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00526 1 2803 695 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00527 5182 697 696 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00528 697 696 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00529 4 2797 696 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00530 2 2797 697 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00531 5182 699 698 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00532 699 698 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00533 3 2797 698 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00534 1 2797 699 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00535 5182 701 700 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00536 701 700 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00537 4 2799 700 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00538 2 2799 701 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00539 5182 703 702 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00540 703 702 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00541 3 2799 702 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00542 1 2799 703 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00543 5182 705 704 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00544 705 704 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00545 4 2801 704 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00546 2 2801 705 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00547 5182 707 706 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00548 707 706 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00549 3 2801 706 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00550 1 2801 707 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00551 5182 709 708 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00552 709 708 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00553 4 2819 708 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00554 2 2819 709 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00555 5182 711 710 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00556 711 710 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00557 3 2819 710 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00558 1 2819 711 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00559 5182 713 712 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00560 713 712 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00561 4 2813 712 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00562 2 2813 713 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00563 5182 715 714 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00564 715 714 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00565 3 2813 714 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00566 1 2813 715 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00567 5182 717 716 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00568 717 716 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00569 4 2815 716 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00570 2 2815 717 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00571 5182 719 718 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00572 719 718 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00573 3 2815 718 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00574 1 2815 719 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00575 5182 721 720 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00576 721 720 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00577 4 2817 720 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00578 2 2817 721 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00579 5182 723 722 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00580 723 722 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00581 3 2817 722 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00582 1 2817 723 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00583 5182 725 724 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00584 725 724 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00585 4 2835 724 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00586 2 2835 725 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00587 5182 727 726 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00588 727 726 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00589 3 2835 726 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00590 1 2835 727 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00591 5182 729 728 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00592 729 728 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00593 4 2829 728 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00594 2 2829 729 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00595 5182 731 730 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00596 731 730 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00597 3 2829 730 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00598 1 2829 731 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00599 5182 733 732 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00600 733 732 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00601 4 2831 732 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00602 2 2831 733 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00603 5182 735 734 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00604 735 734 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00605 3 2831 734 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00606 1 2831 735 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00607 5182 737 736 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00608 737 736 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00609 4 2833 736 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00610 2 2833 737 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00611 5182 739 738 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00612 739 738 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00613 3 2833 738 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00614 1 2833 739 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00615 5182 741 740 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00616 741 740 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00617 4 2851 740 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00618 2 2851 741 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00619 5182 743 742 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00620 743 742 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00621 3 2851 742 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00622 1 2851 743 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00623 5182 745 744 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00624 745 744 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00625 4 2845 744 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00626 2 2845 745 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00627 5182 747 746 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00628 747 746 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00629 3 2845 746 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00630 1 2845 747 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00631 5182 749 748 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00632 749 748 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00633 4 2847 748 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00634 2 2847 749 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00635 5182 751 750 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00636 751 750 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00637 3 2847 750 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00638 1 2847 751 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00639 5182 753 752 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00640 753 752 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00641 4 2849 752 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00642 2 2849 753 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00643 5182 755 754 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00644 755 754 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00645 3 2849 754 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00646 1 2849 755 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00647 5182 757 756 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00648 757 756 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00649 4 2867 756 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00650 2 2867 757 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00651 5182 759 758 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00652 759 758 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00653 3 2867 758 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00654 1 2867 759 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00655 5182 761 760 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00656 761 760 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00657 4 2861 760 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00658 2 2861 761 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00659 5182 763 762 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00660 763 762 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00661 3 2861 762 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00662 1 2861 763 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00663 5182 765 764 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00664 765 764 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00665 4 2863 764 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00666 2 2863 765 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00667 5182 767 766 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00668 767 766 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00669 3 2863 766 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00670 1 2863 767 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00671 5182 769 768 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00672 769 768 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00673 4 2865 768 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00674 2 2865 769 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00675 5182 771 770 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00676 771 770 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00677 3 2865 770 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00678 1 2865 771 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00679 5182 773 772 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00680 773 772 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00681 4 2883 772 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00682 2 2883 773 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00683 5182 775 774 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00684 775 774 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00685 3 2883 774 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00686 1 2883 775 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00687 5182 777 776 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00688 777 776 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00689 4 2877 776 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00690 2 2877 777 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00691 5182 779 778 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00692 779 778 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00693 3 2877 778 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00694 1 2877 779 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00695 5182 781 780 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00696 781 780 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00697 4 2879 780 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00698 2 2879 781 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00699 5182 783 782 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00700 783 782 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00701 3 2879 782 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00702 1 2879 783 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00703 5182 785 784 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00704 785 784 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00705 4 2881 784 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00706 2 2881 785 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00707 5182 787 786 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00708 787 786 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00709 3 2881 786 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00710 1 2881 787 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00711 5182 789 788 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00712 789 788 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00713 4 2899 788 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00714 2 2899 789 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00715 5182 791 790 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00716 791 790 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00717 3 2899 790 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00718 1 2899 791 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00719 5182 793 792 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00720 793 792 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00721 4 2893 792 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00722 2 2893 793 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00723 5182 795 794 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00724 795 794 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00725 3 2893 794 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00726 1 2893 795 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00727 5182 797 796 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00728 797 796 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00729 4 2895 796 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00730 2 2895 797 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00731 5182 799 798 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00732 799 798 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00733 3 2895 798 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00734 1 2895 799 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00735 5182 801 800 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00736 801 800 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00737 4 2897 800 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00738 2 2897 801 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00739 5182 803 802 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00740 803 802 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00741 3 2897 802 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00742 1 2897 803 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00743 5182 805 804 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00744 805 804 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00745 4 2915 804 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00746 2 2915 805 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00747 5182 807 806 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00748 807 806 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00749 3 2915 806 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00750 1 2915 807 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00751 5182 809 808 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00752 809 808 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00753 4 2909 808 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00754 2 2909 809 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00755 5182 811 810 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00756 811 810 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00757 3 2909 810 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00758 1 2909 811 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00759 5182 813 812 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00760 813 812 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00761 4 2911 812 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00762 2 2911 813 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00763 5182 815 814 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00764 815 814 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00765 3 2911 814 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00766 1 2911 815 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00767 5182 817 816 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00768 817 816 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00769 4 2913 816 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00770 2 2913 817 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00771 5182 819 818 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00772 819 818 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00773 3 2913 818 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00774 1 2913 819 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00775 5182 821 820 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00776 821 820 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00777 4 2931 820 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00778 2 2931 821 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00779 5182 823 822 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00780 823 822 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00781 3 2931 822 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00782 1 2931 823 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00783 5182 825 824 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00784 825 824 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00785 4 2925 824 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00786 2 2925 825 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00787 5182 827 826 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00788 827 826 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00789 3 2925 826 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00790 1 2925 827 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00791 5182 829 828 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00792 829 828 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00793 4 2927 828 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00794 2 2927 829 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00795 5182 831 830 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00796 831 830 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00797 3 2927 830 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00798 1 2927 831 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00799 5182 833 832 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00800 833 832 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00801 4 2929 832 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00802 2 2929 833 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00803 5182 835 834 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00804 835 834 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00805 3 2929 834 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00806 1 2929 835 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00807 5182 837 836 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00808 837 836 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00809 4 2947 836 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00810 2 2947 837 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00811 5182 839 838 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00812 839 838 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00813 3 2947 838 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00814 1 2947 839 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00815 5182 841 840 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00816 841 840 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00817 4 2941 840 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00818 2 2941 841 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00819 5182 843 842 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00820 843 842 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00821 3 2941 842 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00822 1 2941 843 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00823 5182 845 844 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00824 845 844 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00825 4 2943 844 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00826 2 2943 845 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00827 5182 847 846 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00828 847 846 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00829 3 2943 846 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00830 1 2943 847 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00831 5182 849 848 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00832 849 848 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00833 4 2945 848 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00834 2 2945 849 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00835 5182 851 850 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00836 851 850 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00837 3 2945 850 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00838 1 2945 851 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00839 5182 853 852 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00840 853 852 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00841 4 2963 852 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00842 2 2963 853 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00843 5182 855 854 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00844 855 854 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00845 3 2963 854 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00846 1 2963 855 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00847 5182 857 856 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00848 857 856 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00849 4 2957 856 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00850 2 2957 857 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00851 5182 859 858 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00852 859 858 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00853 3 2957 858 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00854 1 2957 859 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00855 5182 861 860 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00856 861 860 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00857 4 2959 860 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00858 2 2959 861 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00859 5182 863 862 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00860 863 862 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00861 3 2959 862 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00862 1 2959 863 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00863 5182 865 864 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00864 865 864 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00865 4 2961 864 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00866 2 2961 865 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00867 5182 867 866 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00868 867 866 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00869 3 2961 866 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00870 1 2961 867 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00871 5182 869 868 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00872 869 868 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00873 4 2979 868 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00874 2 2979 869 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00875 5182 871 870 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00876 871 870 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00877 3 2979 870 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00878 1 2979 871 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00879 5182 873 872 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00880 873 872 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00881 4 2973 872 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00882 2 2973 873 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00883 5182 875 874 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00884 875 874 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00885 3 2973 874 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00886 1 2973 875 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00887 5182 877 876 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00888 877 876 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00889 4 2975 876 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00890 2 2975 877 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00891 5182 879 878 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00892 879 878 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00893 3 2975 878 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00894 1 2975 879 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00895 5182 881 880 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00896 881 880 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00897 4 2977 880 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00898 2 2977 881 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00899 5182 883 882 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00900 883 882 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00901 3 2977 882 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00902 1 2977 883 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00903 5182 885 884 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00904 885 884 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00905 4 2995 884 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00906 2 2995 885 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00907 5182 887 886 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00908 887 886 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00909 3 2995 886 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00910 1 2995 887 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00911 5182 889 888 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00912 889 888 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00913 4 2989 888 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00914 2 2989 889 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00915 5182 891 890 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00916 891 890 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00917 3 2989 890 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00918 1 2989 891 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00919 5182 893 892 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00920 893 892 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00921 4 2991 892 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00922 2 2991 893 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00923 5182 895 894 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00924 895 894 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00925 3 2991 894 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00926 1 2991 895 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00927 5182 897 896 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00928 897 896 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00929 4 2993 896 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00930 2 2993 897 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00931 5182 899 898 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00932 899 898 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00933 3 2993 898 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00934 1 2993 899 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00935 5182 901 900 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00936 901 900 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00937 4 3011 900 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00938 2 3011 901 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00939 5182 903 902 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00940 903 902 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00941 3 3011 902 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00942 1 3011 903 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00943 5182 905 904 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00944 905 904 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00945 4 3005 904 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00946 2 3005 905 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00947 5182 907 906 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00948 907 906 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00949 3 3005 906 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00950 1 3005 907 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00951 5182 909 908 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00952 909 908 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00953 4 3007 908 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00954 2 3007 909 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00955 5182 911 910 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00956 911 910 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00957 3 3007 910 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00958 1 3007 911 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00959 5182 913 912 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00960 913 912 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00961 4 3009 912 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00962 2 3009 913 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00963 5182 915 914 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00964 915 914 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00965 3 3009 914 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00966 1 3009 915 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00967 5182 917 916 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00968 917 916 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00969 4 3027 916 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00970 2 3027 917 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00971 5182 919 918 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00972 919 918 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00973 3 3027 918 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00974 1 3027 919 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00975 5182 921 920 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00976 921 920 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00977 4 3021 920 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00978 2 3021 921 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00979 5182 923 922 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00980 923 922 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00981 3 3021 922 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00982 1 3021 923 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00983 5182 925 924 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00984 925 924 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00985 4 3023 924 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00986 2 3023 925 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00987 5182 927 926 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00988 927 926 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00989 3 3023 926 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00990 1 3023 927 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00991 5182 929 928 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00992 929 928 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00993 4 3025 928 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00994 2 3025 929 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00995 5182 931 930 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00996 931 930 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00997 3 3025 930 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00998 1 3025 931 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00999 5182 933 932 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01000 933 932 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01001 4 3043 932 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01002 2 3043 933 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01003 5182 935 934 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01004 935 934 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01005 3 3043 934 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01006 1 3043 935 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01007 5182 937 936 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01008 937 936 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01009 4 3037 936 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01010 2 3037 937 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01011 5182 939 938 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01012 939 938 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01013 3 3037 938 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01014 1 3037 939 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01015 5182 941 940 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01016 941 940 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01017 4 3039 940 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01018 2 3039 941 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01019 5182 943 942 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01020 943 942 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01021 3 3039 942 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01022 1 3039 943 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01023 5182 945 944 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01024 945 944 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01025 4 3041 944 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01026 2 3041 945 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01027 5182 947 946 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01028 947 946 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01029 3 3041 946 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01030 1 3041 947 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01031 1 3045 8 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01032 8 3046 2 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01033 3 3045 9 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01034 9 3046 4 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01035 951 3083 949 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01036 956 951 5 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01037 5 3074 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01038 5 949 948 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01039 5182 3074 6 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01040 950 9 6 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01041 6 8 949 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01042 951 9 7 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01043 7 3074 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01044 7 8 952 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01045 5183 3083 9 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01046 9 3083 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01047 5183 3083 8 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01048 8 3083 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01049 953 3077 9 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_01050 8 3077 954 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_01051 9 3083 8 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_01052 5182 5192 953 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_01053 954 955 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_01054 953 5192 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_01055 5182 955 954 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_01056 5182 5192 955 5182 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01057 5192 957 5182 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01058 5182 957 5192 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01059 5182 3077 957 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01060 957 956 5182 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01061 957 3074 958 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01062 13 2529 11 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01063 13 2529 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01064 11 2529 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01065 12 2529 10 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01066 5183 2529 12 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01067 5183 2529 10 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01068 5182 960 959 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01069 960 959 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01070 13 2547 959 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01071 11 2547 960 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01072 5182 962 961 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01073 962 961 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01074 12 2547 961 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01075 10 2547 962 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01076 5182 964 963 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01077 964 963 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01078 13 2541 963 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01079 11 2541 964 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01080 5182 966 965 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01081 966 965 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01082 12 2541 965 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01083 10 2541 966 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01084 5182 968 967 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01085 968 967 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01086 13 2543 967 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01087 11 2543 968 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01088 5182 970 969 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01089 970 969 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01090 12 2543 969 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01091 10 2543 970 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01092 5182 972 971 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01093 972 971 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01094 13 2545 971 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01095 11 2545 972 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01096 5182 974 973 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01097 974 973 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01098 12 2545 973 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01099 10 2545 974 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01100 5182 976 975 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01101 976 975 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01102 13 2563 975 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01103 11 2563 976 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01104 5182 978 977 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01105 978 977 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01106 12 2563 977 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01107 10 2563 978 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01108 5182 980 979 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01109 980 979 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01110 13 2557 979 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01111 11 2557 980 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01112 5182 982 981 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01113 982 981 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01114 12 2557 981 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01115 10 2557 982 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01116 5182 984 983 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01117 984 983 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01118 13 2559 983 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01119 11 2559 984 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01120 5182 986 985 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01121 986 985 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01122 12 2559 985 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01123 10 2559 986 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01124 5182 988 987 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01125 988 987 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01126 13 2561 987 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01127 11 2561 988 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01128 5182 990 989 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01129 990 989 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01130 12 2561 989 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01131 10 2561 990 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01132 5182 992 991 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01133 992 991 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01134 13 2579 991 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01135 11 2579 992 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01136 5182 994 993 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01137 994 993 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01138 12 2579 993 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01139 10 2579 994 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01140 5182 996 995 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01141 996 995 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01142 13 2573 995 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01143 11 2573 996 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01144 5182 998 997 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01145 998 997 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01146 12 2573 997 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01147 10 2573 998 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01148 5182 1000 999 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01149 1000 999 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01150 13 2575 999 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01151 11 2575 1000 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01152 5182 1002 1001 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01153 1002 1001 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01154 12 2575 1001 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01155 10 2575 1002 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01156 5182 1004 1003 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01157 1004 1003 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01158 13 2577 1003 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01159 11 2577 1004 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01160 5182 1006 1005 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01161 1006 1005 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01162 12 2577 1005 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01163 10 2577 1006 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01164 5182 1008 1007 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01165 1008 1007 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01166 13 2595 1007 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01167 11 2595 1008 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01168 5182 1010 1009 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01169 1010 1009 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01170 12 2595 1009 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01171 10 2595 1010 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01172 5182 1012 1011 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01173 1012 1011 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01174 13 2589 1011 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01175 11 2589 1012 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01176 5182 1014 1013 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01177 1014 1013 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01178 12 2589 1013 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01179 10 2589 1014 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01180 5182 1016 1015 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01181 1016 1015 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01182 13 2591 1015 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01183 11 2591 1016 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01184 5182 1018 1017 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01185 1018 1017 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01186 12 2591 1017 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01187 10 2591 1018 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01188 5182 1020 1019 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01189 1020 1019 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01190 13 2593 1019 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01191 11 2593 1020 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01192 5182 1022 1021 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01193 1022 1021 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01194 12 2593 1021 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01195 10 2593 1022 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01196 5182 1024 1023 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01197 1024 1023 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01198 13 2611 1023 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01199 11 2611 1024 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01200 5182 1026 1025 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01201 1026 1025 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01202 12 2611 1025 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01203 10 2611 1026 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01204 5182 1028 1027 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01205 1028 1027 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01206 13 2605 1027 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01207 11 2605 1028 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01208 5182 1030 1029 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01209 1030 1029 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01210 12 2605 1029 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01211 10 2605 1030 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01212 5182 1032 1031 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01213 1032 1031 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01214 13 2607 1031 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01215 11 2607 1032 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01216 5182 1034 1033 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01217 1034 1033 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01218 12 2607 1033 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01219 10 2607 1034 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01220 5182 1036 1035 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01221 1036 1035 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01222 13 2609 1035 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01223 11 2609 1036 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01224 5182 1038 1037 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01225 1038 1037 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01226 12 2609 1037 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01227 10 2609 1038 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01228 5182 1040 1039 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01229 1040 1039 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01230 13 2627 1039 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01231 11 2627 1040 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01232 5182 1042 1041 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01233 1042 1041 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01234 12 2627 1041 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01235 10 2627 1042 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01236 5182 1044 1043 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01237 1044 1043 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01238 13 2621 1043 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01239 11 2621 1044 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01240 5182 1046 1045 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01241 1046 1045 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01242 12 2621 1045 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01243 10 2621 1046 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01244 5182 1048 1047 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01245 1048 1047 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01246 13 2623 1047 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01247 11 2623 1048 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01248 5182 1050 1049 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01249 1050 1049 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01250 12 2623 1049 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01251 10 2623 1050 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01252 5182 1052 1051 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01253 1052 1051 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01254 13 2625 1051 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01255 11 2625 1052 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01256 5182 1054 1053 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01257 1054 1053 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01258 12 2625 1053 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01259 10 2625 1054 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01260 5182 1056 1055 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01261 1056 1055 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01262 13 2643 1055 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01263 11 2643 1056 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01264 5182 1058 1057 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01265 1058 1057 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01266 12 2643 1057 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01267 10 2643 1058 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01268 5182 1060 1059 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01269 1060 1059 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01270 13 2637 1059 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01271 11 2637 1060 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01272 5182 1062 1061 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01273 1062 1061 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01274 12 2637 1061 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01275 10 2637 1062 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01276 5182 1064 1063 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01277 1064 1063 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01278 13 2639 1063 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01279 11 2639 1064 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01280 5182 1066 1065 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01281 1066 1065 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01282 12 2639 1065 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01283 10 2639 1066 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01284 5182 1068 1067 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01285 1068 1067 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01286 13 2641 1067 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01287 11 2641 1068 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01288 5182 1070 1069 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01289 1070 1069 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01290 12 2641 1069 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01291 10 2641 1070 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01292 5182 1072 1071 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01293 1072 1071 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01294 13 2659 1071 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01295 11 2659 1072 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01296 5182 1074 1073 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01297 1074 1073 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01298 12 2659 1073 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01299 10 2659 1074 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01300 5182 1076 1075 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01301 1076 1075 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01302 13 2653 1075 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01303 11 2653 1076 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01304 5182 1078 1077 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01305 1078 1077 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01306 12 2653 1077 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01307 10 2653 1078 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01308 5182 1080 1079 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01309 1080 1079 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01310 13 2655 1079 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01311 11 2655 1080 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01312 5182 1082 1081 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01313 1082 1081 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01314 12 2655 1081 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01315 10 2655 1082 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01316 5182 1084 1083 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01317 1084 1083 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01318 13 2657 1083 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01319 11 2657 1084 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01320 5182 1086 1085 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01321 1086 1085 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01322 12 2657 1085 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01323 10 2657 1086 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01324 5182 1088 1087 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01325 1088 1087 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01326 13 2675 1087 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01327 11 2675 1088 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01328 5182 1090 1089 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01329 1090 1089 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01330 12 2675 1089 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01331 10 2675 1090 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01332 5182 1092 1091 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01333 1092 1091 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01334 13 2669 1091 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01335 11 2669 1092 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01336 5182 1094 1093 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01337 1094 1093 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01338 12 2669 1093 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01339 10 2669 1094 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01340 5182 1096 1095 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01341 1096 1095 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01342 13 2671 1095 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01343 11 2671 1096 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01344 5182 1098 1097 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01345 1098 1097 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01346 12 2671 1097 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01347 10 2671 1098 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01348 5182 1100 1099 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01349 1100 1099 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01350 13 2673 1099 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01351 11 2673 1100 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01352 5182 1102 1101 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01353 1102 1101 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01354 12 2673 1101 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01355 10 2673 1102 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01356 5182 1104 1103 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01357 1104 1103 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01358 13 2691 1103 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01359 11 2691 1104 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01360 5182 1106 1105 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01361 1106 1105 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01362 12 2691 1105 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01363 10 2691 1106 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01364 5182 1108 1107 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01365 1108 1107 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01366 13 2685 1107 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01367 11 2685 1108 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01368 5182 1110 1109 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01369 1110 1109 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01370 12 2685 1109 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01371 10 2685 1110 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01372 5182 1112 1111 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01373 1112 1111 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01374 13 2687 1111 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01375 11 2687 1112 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01376 5182 1114 1113 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01377 1114 1113 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01378 12 2687 1113 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01379 10 2687 1114 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01380 5182 1116 1115 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01381 1116 1115 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01382 13 2689 1115 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01383 11 2689 1116 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01384 5182 1118 1117 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01385 1118 1117 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01386 12 2689 1117 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01387 10 2689 1118 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01388 5182 1120 1119 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01389 1120 1119 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01390 13 2707 1119 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01391 11 2707 1120 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01392 5182 1122 1121 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01393 1122 1121 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01394 12 2707 1121 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01395 10 2707 1122 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01396 5182 1124 1123 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01397 1124 1123 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01398 13 2701 1123 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01399 11 2701 1124 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01400 5182 1126 1125 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01401 1126 1125 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01402 12 2701 1125 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01403 10 2701 1126 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01404 5182 1128 1127 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01405 1128 1127 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01406 13 2703 1127 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01407 11 2703 1128 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01408 5182 1130 1129 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01409 1130 1129 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01410 12 2703 1129 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01411 10 2703 1130 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01412 5182 1132 1131 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01413 1132 1131 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01414 13 2705 1131 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01415 11 2705 1132 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01416 5182 1134 1133 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01417 1134 1133 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01418 12 2705 1133 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01419 10 2705 1134 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01420 5182 1136 1135 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01421 1136 1135 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01422 13 2723 1135 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01423 11 2723 1136 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01424 5182 1138 1137 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01425 1138 1137 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01426 12 2723 1137 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01427 10 2723 1138 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01428 5182 1140 1139 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01429 1140 1139 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01430 13 2717 1139 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01431 11 2717 1140 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01432 5182 1142 1141 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01433 1142 1141 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01434 12 2717 1141 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01435 10 2717 1142 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01436 5182 1144 1143 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01437 1144 1143 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01438 13 2719 1143 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01439 11 2719 1144 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01440 5182 1146 1145 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01441 1146 1145 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01442 12 2719 1145 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01443 10 2719 1146 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01444 5182 1148 1147 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01445 1148 1147 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01446 13 2721 1147 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01447 11 2721 1148 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01448 5182 1150 1149 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01449 1150 1149 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01450 12 2721 1149 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01451 10 2721 1150 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01452 5182 1152 1151 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01453 1152 1151 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01454 13 2739 1151 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01455 11 2739 1152 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01456 5182 1154 1153 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01457 1154 1153 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01458 12 2739 1153 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01459 10 2739 1154 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01460 5182 1156 1155 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01461 1156 1155 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01462 13 2733 1155 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01463 11 2733 1156 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01464 5182 1158 1157 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01465 1158 1157 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01466 12 2733 1157 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01467 10 2733 1158 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01468 5182 1160 1159 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01469 1160 1159 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01470 13 2735 1159 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01471 11 2735 1160 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01472 5182 1162 1161 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01473 1162 1161 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01474 12 2735 1161 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01475 10 2735 1162 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01476 5182 1164 1163 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01477 1164 1163 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01478 13 2737 1163 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01479 11 2737 1164 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01480 5182 1166 1165 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01481 1166 1165 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01482 12 2737 1165 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01483 10 2737 1166 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01484 5182 1168 1167 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01485 1168 1167 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01486 13 2755 1167 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01487 11 2755 1168 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01488 5182 1170 1169 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01489 1170 1169 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01490 12 2755 1169 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01491 10 2755 1170 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01492 5182 1172 1171 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01493 1172 1171 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01494 13 2749 1171 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01495 11 2749 1172 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01496 5182 1174 1173 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01497 1174 1173 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01498 12 2749 1173 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01499 10 2749 1174 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01500 5182 1176 1175 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01501 1176 1175 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01502 13 2751 1175 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01503 11 2751 1176 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01504 5182 1178 1177 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01505 1178 1177 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01506 12 2751 1177 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01507 10 2751 1178 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01508 5182 1180 1179 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01509 1180 1179 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01510 13 2753 1179 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01511 11 2753 1180 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01512 5182 1182 1181 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01513 1182 1181 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01514 12 2753 1181 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01515 10 2753 1182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01516 5182 1184 1183 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01517 1184 1183 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01518 13 2771 1183 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01519 11 2771 1184 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01520 5182 1186 1185 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01521 1186 1185 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01522 12 2771 1185 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01523 10 2771 1186 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01524 5182 1188 1187 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01525 1188 1187 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01526 13 2765 1187 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01527 11 2765 1188 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01528 5182 1190 1189 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01529 1190 1189 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01530 12 2765 1189 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01531 10 2765 1190 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01532 5182 1192 1191 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01533 1192 1191 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01534 13 2767 1191 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01535 11 2767 1192 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01536 5182 1194 1193 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01537 1194 1193 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01538 12 2767 1193 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01539 10 2767 1194 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01540 5182 1196 1195 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01541 1196 1195 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01542 13 2769 1195 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01543 11 2769 1196 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01544 5182 1198 1197 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01545 1198 1197 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01546 12 2769 1197 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01547 10 2769 1198 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01548 5182 1200 1199 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01549 1200 1199 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01550 13 2787 1199 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01551 11 2787 1200 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01552 5182 1202 1201 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01553 1202 1201 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01554 12 2787 1201 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01555 10 2787 1202 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01556 5182 1204 1203 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01557 1204 1203 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01558 13 2781 1203 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01559 11 2781 1204 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01560 5182 1206 1205 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01561 1206 1205 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01562 12 2781 1205 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01563 10 2781 1206 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01564 5182 1208 1207 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01565 1208 1207 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01566 13 2783 1207 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01567 11 2783 1208 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01568 5182 1210 1209 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01569 1210 1209 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01570 12 2783 1209 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01571 10 2783 1210 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01572 5182 1212 1211 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01573 1212 1211 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01574 13 2785 1211 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01575 11 2785 1212 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01576 5182 1214 1213 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01577 1214 1213 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01578 12 2785 1213 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01579 10 2785 1214 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01580 5182 1216 1215 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01581 1216 1215 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01582 13 2803 1215 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01583 11 2803 1216 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01584 5182 1218 1217 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01585 1218 1217 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01586 12 2803 1217 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01587 10 2803 1218 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01588 5182 1220 1219 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01589 1220 1219 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01590 13 2797 1219 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01591 11 2797 1220 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01592 5182 1222 1221 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01593 1222 1221 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01594 12 2797 1221 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01595 10 2797 1222 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01596 5182 1224 1223 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01597 1224 1223 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01598 13 2799 1223 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01599 11 2799 1224 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01600 5182 1226 1225 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01601 1226 1225 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01602 12 2799 1225 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01603 10 2799 1226 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01604 5182 1228 1227 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01605 1228 1227 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01606 13 2801 1227 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01607 11 2801 1228 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01608 5182 1230 1229 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01609 1230 1229 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01610 12 2801 1229 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01611 10 2801 1230 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01612 5182 1232 1231 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01613 1232 1231 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01614 13 2819 1231 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01615 11 2819 1232 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01616 5182 1234 1233 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01617 1234 1233 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01618 12 2819 1233 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01619 10 2819 1234 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01620 5182 1236 1235 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01621 1236 1235 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01622 13 2813 1235 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01623 11 2813 1236 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01624 5182 1238 1237 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01625 1238 1237 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01626 12 2813 1237 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01627 10 2813 1238 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01628 5182 1240 1239 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01629 1240 1239 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01630 13 2815 1239 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01631 11 2815 1240 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01632 5182 1242 1241 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01633 1242 1241 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01634 12 2815 1241 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01635 10 2815 1242 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01636 5182 1244 1243 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01637 1244 1243 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01638 13 2817 1243 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01639 11 2817 1244 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01640 5182 1246 1245 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01641 1246 1245 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01642 12 2817 1245 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01643 10 2817 1246 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01644 5182 1248 1247 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01645 1248 1247 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01646 13 2835 1247 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01647 11 2835 1248 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01648 5182 1250 1249 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01649 1250 1249 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01650 12 2835 1249 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01651 10 2835 1250 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01652 5182 1252 1251 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01653 1252 1251 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01654 13 2829 1251 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01655 11 2829 1252 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01656 5182 1254 1253 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01657 1254 1253 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01658 12 2829 1253 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01659 10 2829 1254 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01660 5182 1256 1255 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01661 1256 1255 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01662 13 2831 1255 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01663 11 2831 1256 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01664 5182 1258 1257 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01665 1258 1257 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01666 12 2831 1257 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01667 10 2831 1258 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01668 5182 1260 1259 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01669 1260 1259 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01670 13 2833 1259 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01671 11 2833 1260 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01672 5182 1262 1261 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01673 1262 1261 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01674 12 2833 1261 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01675 10 2833 1262 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01676 5182 1264 1263 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01677 1264 1263 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01678 13 2851 1263 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01679 11 2851 1264 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01680 5182 1266 1265 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01681 1266 1265 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01682 12 2851 1265 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01683 10 2851 1266 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01684 5182 1268 1267 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01685 1268 1267 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01686 13 2845 1267 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01687 11 2845 1268 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01688 5182 1270 1269 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01689 1270 1269 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01690 12 2845 1269 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01691 10 2845 1270 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01692 5182 1272 1271 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01693 1272 1271 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01694 13 2847 1271 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01695 11 2847 1272 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01696 5182 1274 1273 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01697 1274 1273 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01698 12 2847 1273 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01699 10 2847 1274 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01700 5182 1276 1275 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01701 1276 1275 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01702 13 2849 1275 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01703 11 2849 1276 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01704 5182 1278 1277 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01705 1278 1277 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01706 12 2849 1277 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01707 10 2849 1278 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01708 5182 1280 1279 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01709 1280 1279 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01710 13 2867 1279 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01711 11 2867 1280 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01712 5182 1282 1281 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01713 1282 1281 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01714 12 2867 1281 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01715 10 2867 1282 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01716 5182 1284 1283 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01717 1284 1283 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01718 13 2861 1283 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01719 11 2861 1284 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01720 5182 1286 1285 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01721 1286 1285 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01722 12 2861 1285 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01723 10 2861 1286 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01724 5182 1288 1287 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01725 1288 1287 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01726 13 2863 1287 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01727 11 2863 1288 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01728 5182 1290 1289 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01729 1290 1289 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01730 12 2863 1289 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01731 10 2863 1290 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01732 5182 1292 1291 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01733 1292 1291 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01734 13 2865 1291 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01735 11 2865 1292 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01736 5182 1294 1293 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01737 1294 1293 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01738 12 2865 1293 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01739 10 2865 1294 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01740 5182 1296 1295 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01741 1296 1295 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01742 13 2883 1295 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01743 11 2883 1296 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01744 5182 1298 1297 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01745 1298 1297 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01746 12 2883 1297 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01747 10 2883 1298 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01748 5182 1300 1299 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01749 1300 1299 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01750 13 2877 1299 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01751 11 2877 1300 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01752 5182 1302 1301 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01753 1302 1301 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01754 12 2877 1301 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01755 10 2877 1302 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01756 5182 1304 1303 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01757 1304 1303 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01758 13 2879 1303 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01759 11 2879 1304 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01760 5182 1306 1305 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01761 1306 1305 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01762 12 2879 1305 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01763 10 2879 1306 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01764 5182 1308 1307 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01765 1308 1307 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01766 13 2881 1307 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01767 11 2881 1308 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01768 5182 1310 1309 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01769 1310 1309 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01770 12 2881 1309 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01771 10 2881 1310 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01772 5182 1312 1311 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01773 1312 1311 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01774 13 2899 1311 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01775 11 2899 1312 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01776 5182 1314 1313 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01777 1314 1313 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01778 12 2899 1313 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01779 10 2899 1314 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01780 5182 1316 1315 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01781 1316 1315 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01782 13 2893 1315 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01783 11 2893 1316 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01784 5182 1318 1317 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01785 1318 1317 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01786 12 2893 1317 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01787 10 2893 1318 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01788 5182 1320 1319 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01789 1320 1319 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01790 13 2895 1319 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01791 11 2895 1320 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01792 5182 1322 1321 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01793 1322 1321 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01794 12 2895 1321 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01795 10 2895 1322 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01796 5182 1324 1323 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01797 1324 1323 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01798 13 2897 1323 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01799 11 2897 1324 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01800 5182 1326 1325 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01801 1326 1325 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01802 12 2897 1325 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01803 10 2897 1326 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01804 5182 1328 1327 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01805 1328 1327 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01806 13 2915 1327 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01807 11 2915 1328 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01808 5182 1330 1329 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01809 1330 1329 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01810 12 2915 1329 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01811 10 2915 1330 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01812 5182 1332 1331 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01813 1332 1331 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01814 13 2909 1331 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01815 11 2909 1332 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01816 5182 1334 1333 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01817 1334 1333 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01818 12 2909 1333 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01819 10 2909 1334 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01820 5182 1336 1335 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01821 1336 1335 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01822 13 2911 1335 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01823 11 2911 1336 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01824 5182 1338 1337 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01825 1338 1337 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01826 12 2911 1337 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01827 10 2911 1338 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01828 5182 1340 1339 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01829 1340 1339 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01830 13 2913 1339 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01831 11 2913 1340 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01832 5182 1342 1341 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01833 1342 1341 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01834 12 2913 1341 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01835 10 2913 1342 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01836 5182 1344 1343 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01837 1344 1343 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01838 13 2931 1343 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01839 11 2931 1344 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01840 5182 1346 1345 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01841 1346 1345 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01842 12 2931 1345 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01843 10 2931 1346 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01844 5182 1348 1347 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01845 1348 1347 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01846 13 2925 1347 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01847 11 2925 1348 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01848 5182 1350 1349 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01849 1350 1349 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01850 12 2925 1349 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01851 10 2925 1350 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01852 5182 1352 1351 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01853 1352 1351 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01854 13 2927 1351 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01855 11 2927 1352 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01856 5182 1354 1353 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01857 1354 1353 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01858 12 2927 1353 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01859 10 2927 1354 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01860 5182 1356 1355 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01861 1356 1355 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01862 13 2929 1355 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01863 11 2929 1356 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01864 5182 1358 1357 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01865 1358 1357 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01866 12 2929 1357 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01867 10 2929 1358 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01868 5182 1360 1359 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01869 1360 1359 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01870 13 2947 1359 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01871 11 2947 1360 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01872 5182 1362 1361 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01873 1362 1361 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01874 12 2947 1361 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01875 10 2947 1362 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01876 5182 1364 1363 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01877 1364 1363 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01878 13 2941 1363 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01879 11 2941 1364 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01880 5182 1366 1365 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01881 1366 1365 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01882 12 2941 1365 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01883 10 2941 1366 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01884 5182 1368 1367 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01885 1368 1367 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01886 13 2943 1367 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01887 11 2943 1368 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01888 5182 1370 1369 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01889 1370 1369 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01890 12 2943 1369 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01891 10 2943 1370 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01892 5182 1372 1371 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01893 1372 1371 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01894 13 2945 1371 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01895 11 2945 1372 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01896 5182 1374 1373 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01897 1374 1373 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01898 12 2945 1373 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01899 10 2945 1374 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01900 5182 1376 1375 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01901 1376 1375 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01902 13 2963 1375 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01903 11 2963 1376 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01904 5182 1378 1377 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01905 1378 1377 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01906 12 2963 1377 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01907 10 2963 1378 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01908 5182 1380 1379 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01909 1380 1379 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01910 13 2957 1379 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01911 11 2957 1380 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01912 5182 1382 1381 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01913 1382 1381 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01914 12 2957 1381 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01915 10 2957 1382 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01916 5182 1384 1383 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01917 1384 1383 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01918 13 2959 1383 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01919 11 2959 1384 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01920 5182 1386 1385 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01921 1386 1385 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01922 12 2959 1385 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01923 10 2959 1386 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01924 5182 1388 1387 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01925 1388 1387 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01926 13 2961 1387 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01927 11 2961 1388 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01928 5182 1390 1389 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01929 1390 1389 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01930 12 2961 1389 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01931 10 2961 1390 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01932 5182 1392 1391 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01933 1392 1391 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01934 13 2979 1391 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01935 11 2979 1392 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01936 5182 1394 1393 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01937 1394 1393 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01938 12 2979 1393 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01939 10 2979 1394 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01940 5182 1396 1395 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01941 1396 1395 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01942 13 2973 1395 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01943 11 2973 1396 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01944 5182 1398 1397 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01945 1398 1397 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01946 12 2973 1397 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01947 10 2973 1398 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01948 5182 1400 1399 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01949 1400 1399 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01950 13 2975 1399 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01951 11 2975 1400 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01952 5182 1402 1401 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01953 1402 1401 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01954 12 2975 1401 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01955 10 2975 1402 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01956 5182 1404 1403 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01957 1404 1403 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01958 13 2977 1403 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01959 11 2977 1404 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01960 5182 1406 1405 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01961 1406 1405 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01962 12 2977 1405 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01963 10 2977 1406 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01964 5182 1408 1407 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01965 1408 1407 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01966 13 2995 1407 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01967 11 2995 1408 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01968 5182 1410 1409 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01969 1410 1409 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01970 12 2995 1409 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01971 10 2995 1410 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01972 5182 1412 1411 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01973 1412 1411 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01974 13 2989 1411 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01975 11 2989 1412 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01976 5182 1414 1413 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01977 1414 1413 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01978 12 2989 1413 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01979 10 2989 1414 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01980 5182 1416 1415 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01981 1416 1415 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01982 13 2991 1415 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01983 11 2991 1416 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01984 5182 1418 1417 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01985 1418 1417 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01986 12 2991 1417 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01987 10 2991 1418 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01988 5182 1420 1419 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01989 1420 1419 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01990 13 2993 1419 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01991 11 2993 1420 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01992 5182 1422 1421 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01993 1422 1421 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01994 12 2993 1421 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01995 10 2993 1422 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01996 5182 1424 1423 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01997 1424 1423 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01998 13 3011 1423 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01999 11 3011 1424 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02000 5182 1426 1425 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02001 1426 1425 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02002 12 3011 1425 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02003 10 3011 1426 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02004 5182 1428 1427 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02005 1428 1427 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02006 13 3005 1427 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02007 11 3005 1428 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02008 5182 1430 1429 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02009 1430 1429 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02010 12 3005 1429 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02011 10 3005 1430 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02012 5182 1432 1431 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02013 1432 1431 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02014 13 3007 1431 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02015 11 3007 1432 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02016 5182 1434 1433 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02017 1434 1433 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02018 12 3007 1433 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02019 10 3007 1434 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02020 5182 1436 1435 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02021 1436 1435 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02022 13 3009 1435 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02023 11 3009 1436 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02024 5182 1438 1437 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02025 1438 1437 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02026 12 3009 1437 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02027 10 3009 1438 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02028 5182 1440 1439 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02029 1440 1439 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02030 13 3027 1439 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02031 11 3027 1440 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02032 5182 1442 1441 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02033 1442 1441 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02034 12 3027 1441 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02035 10 3027 1442 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02036 5182 1444 1443 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02037 1444 1443 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02038 13 3021 1443 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02039 11 3021 1444 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02040 5182 1446 1445 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02041 1446 1445 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02042 12 3021 1445 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02043 10 3021 1446 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02044 5182 1448 1447 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02045 1448 1447 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02046 13 3023 1447 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02047 11 3023 1448 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02048 5182 1450 1449 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02049 1450 1449 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02050 12 3023 1449 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02051 10 3023 1450 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02052 5182 1452 1451 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02053 1452 1451 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02054 13 3025 1451 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02055 11 3025 1452 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02056 5182 1454 1453 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02057 1454 1453 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02058 12 3025 1453 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02059 10 3025 1454 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02060 5182 1456 1455 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02061 1456 1455 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02062 13 3043 1455 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02063 11 3043 1456 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02064 5182 1458 1457 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02065 1458 1457 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02066 12 3043 1457 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02067 10 3043 1458 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02068 5182 1460 1459 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02069 1460 1459 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02070 13 3037 1459 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02071 11 3037 1460 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02072 5182 1462 1461 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02073 1462 1461 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02074 12 3037 1461 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02075 10 3037 1462 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02076 5182 1464 1463 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02077 1464 1463 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02078 13 3039 1463 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02079 11 3039 1464 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02080 5182 1466 1465 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02081 1466 1465 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02082 12 3039 1465 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02083 10 3039 1466 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02084 5182 1468 1467 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02085 1468 1467 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02086 13 3041 1467 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02087 11 3041 1468 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02088 5182 1470 1469 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02089 1470 1469 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02090 12 3041 1469 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02091 10 3041 1470 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02092 10 3045 17 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02093 17 3046 11 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02094 12 3045 18 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02095 18 3046 13 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02096 1474 3083 1472 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02097 1479 1474 14 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02098 14 3074 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02099 14 1472 1471 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02100 5182 3074 15 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02101 1473 18 15 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02102 15 17 1472 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02103 1474 18 16 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02104 16 3074 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02105 16 17 1475 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02106 5183 3083 18 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02107 18 3083 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02108 5183 3083 17 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02109 17 3083 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02110 1476 3077 18 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_02111 17 3077 1477 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_02112 18 3083 17 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_02113 5182 5191 1476 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_02114 1477 1478 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_02115 1476 5191 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_02116 5182 1478 1477 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_02117 5182 5191 1478 5182 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02118 5191 1480 5182 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02119 5182 1480 5191 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02120 5182 3077 1480 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02121 1480 1479 5182 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02122 1480 3074 1481 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02123 22 2529 20 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02124 22 2529 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02125 20 2529 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02126 21 2529 19 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02127 5183 2529 21 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02128 5183 2529 19 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02129 5182 1483 1482 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02130 1483 1482 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02131 22 2547 1482 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02132 20 2547 1483 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02133 5182 1485 1484 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02134 1485 1484 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02135 21 2547 1484 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02136 19 2547 1485 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02137 5182 1487 1486 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02138 1487 1486 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02139 22 2541 1486 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02140 20 2541 1487 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02141 5182 1489 1488 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02142 1489 1488 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02143 21 2541 1488 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02144 19 2541 1489 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02145 5182 1491 1490 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02146 1491 1490 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02147 22 2543 1490 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02148 20 2543 1491 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02149 5182 1493 1492 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02150 1493 1492 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02151 21 2543 1492 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02152 19 2543 1493 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02153 5182 1495 1494 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02154 1495 1494 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02155 22 2545 1494 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02156 20 2545 1495 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02157 5182 1497 1496 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02158 1497 1496 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02159 21 2545 1496 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02160 19 2545 1497 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02161 5182 1499 1498 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02162 1499 1498 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02163 22 2563 1498 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02164 20 2563 1499 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02165 5182 1501 1500 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02166 1501 1500 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02167 21 2563 1500 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02168 19 2563 1501 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02169 5182 1503 1502 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02170 1503 1502 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02171 22 2557 1502 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02172 20 2557 1503 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02173 5182 1505 1504 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02174 1505 1504 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02175 21 2557 1504 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02176 19 2557 1505 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02177 5182 1507 1506 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02178 1507 1506 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02179 22 2559 1506 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02180 20 2559 1507 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02181 5182 1509 1508 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02182 1509 1508 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02183 21 2559 1508 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02184 19 2559 1509 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02185 5182 1511 1510 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02186 1511 1510 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02187 22 2561 1510 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02188 20 2561 1511 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02189 5182 1513 1512 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02190 1513 1512 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02191 21 2561 1512 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02192 19 2561 1513 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02193 5182 1515 1514 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02194 1515 1514 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02195 22 2579 1514 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02196 20 2579 1515 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02197 5182 1517 1516 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02198 1517 1516 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02199 21 2579 1516 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02200 19 2579 1517 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02201 5182 1519 1518 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02202 1519 1518 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02203 22 2573 1518 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02204 20 2573 1519 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02205 5182 1521 1520 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02206 1521 1520 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02207 21 2573 1520 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02208 19 2573 1521 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02209 5182 1523 1522 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02210 1523 1522 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02211 22 2575 1522 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02212 20 2575 1523 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02213 5182 1525 1524 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02214 1525 1524 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02215 21 2575 1524 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02216 19 2575 1525 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02217 5182 1527 1526 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02218 1527 1526 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02219 22 2577 1526 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02220 20 2577 1527 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02221 5182 1529 1528 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02222 1529 1528 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02223 21 2577 1528 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02224 19 2577 1529 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02225 5182 1531 1530 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02226 1531 1530 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02227 22 2595 1530 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02228 20 2595 1531 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02229 5182 1533 1532 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02230 1533 1532 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02231 21 2595 1532 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02232 19 2595 1533 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02233 5182 1535 1534 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02234 1535 1534 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02235 22 2589 1534 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02236 20 2589 1535 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02237 5182 1537 1536 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02238 1537 1536 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02239 21 2589 1536 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02240 19 2589 1537 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02241 5182 1539 1538 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02242 1539 1538 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02243 22 2591 1538 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02244 20 2591 1539 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02245 5182 1541 1540 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02246 1541 1540 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02247 21 2591 1540 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02248 19 2591 1541 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02249 5182 1543 1542 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02250 1543 1542 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02251 22 2593 1542 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02252 20 2593 1543 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02253 5182 1545 1544 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02254 1545 1544 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02255 21 2593 1544 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02256 19 2593 1545 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02257 5182 1547 1546 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02258 1547 1546 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02259 22 2611 1546 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02260 20 2611 1547 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02261 5182 1549 1548 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02262 1549 1548 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02263 21 2611 1548 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02264 19 2611 1549 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02265 5182 1551 1550 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02266 1551 1550 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02267 22 2605 1550 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02268 20 2605 1551 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02269 5182 1553 1552 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02270 1553 1552 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02271 21 2605 1552 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02272 19 2605 1553 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02273 5182 1555 1554 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02274 1555 1554 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02275 22 2607 1554 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02276 20 2607 1555 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02277 5182 1557 1556 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02278 1557 1556 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02279 21 2607 1556 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02280 19 2607 1557 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02281 5182 1559 1558 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02282 1559 1558 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02283 22 2609 1558 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02284 20 2609 1559 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02285 5182 1561 1560 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02286 1561 1560 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02287 21 2609 1560 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02288 19 2609 1561 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02289 5182 1563 1562 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02290 1563 1562 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02291 22 2627 1562 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02292 20 2627 1563 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02293 5182 1565 1564 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02294 1565 1564 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02295 21 2627 1564 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02296 19 2627 1565 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02297 5182 1567 1566 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02298 1567 1566 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02299 22 2621 1566 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02300 20 2621 1567 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02301 5182 1569 1568 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02302 1569 1568 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02303 21 2621 1568 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02304 19 2621 1569 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02305 5182 1571 1570 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02306 1571 1570 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02307 22 2623 1570 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02308 20 2623 1571 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02309 5182 1573 1572 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02310 1573 1572 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02311 21 2623 1572 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02312 19 2623 1573 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02313 5182 1575 1574 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02314 1575 1574 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02315 22 2625 1574 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02316 20 2625 1575 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02317 5182 1577 1576 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02318 1577 1576 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02319 21 2625 1576 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02320 19 2625 1577 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02321 5182 1579 1578 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02322 1579 1578 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02323 22 2643 1578 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02324 20 2643 1579 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02325 5182 1581 1580 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02326 1581 1580 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02327 21 2643 1580 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02328 19 2643 1581 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02329 5182 1583 1582 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02330 1583 1582 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02331 22 2637 1582 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02332 20 2637 1583 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02333 5182 1585 1584 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02334 1585 1584 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02335 21 2637 1584 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02336 19 2637 1585 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02337 5182 1587 1586 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02338 1587 1586 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02339 22 2639 1586 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02340 20 2639 1587 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02341 5182 1589 1588 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02342 1589 1588 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02343 21 2639 1588 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02344 19 2639 1589 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02345 5182 1591 1590 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02346 1591 1590 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02347 22 2641 1590 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02348 20 2641 1591 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02349 5182 1593 1592 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02350 1593 1592 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02351 21 2641 1592 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02352 19 2641 1593 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02353 5182 1595 1594 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02354 1595 1594 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02355 22 2659 1594 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02356 20 2659 1595 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02357 5182 1597 1596 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02358 1597 1596 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02359 21 2659 1596 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02360 19 2659 1597 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02361 5182 1599 1598 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02362 1599 1598 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02363 22 2653 1598 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02364 20 2653 1599 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02365 5182 1601 1600 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02366 1601 1600 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02367 21 2653 1600 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02368 19 2653 1601 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02369 5182 1603 1602 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02370 1603 1602 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02371 22 2655 1602 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02372 20 2655 1603 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02373 5182 1605 1604 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02374 1605 1604 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02375 21 2655 1604 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02376 19 2655 1605 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02377 5182 1607 1606 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02378 1607 1606 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02379 22 2657 1606 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02380 20 2657 1607 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02381 5182 1609 1608 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02382 1609 1608 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02383 21 2657 1608 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02384 19 2657 1609 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02385 5182 1611 1610 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02386 1611 1610 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02387 22 2675 1610 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02388 20 2675 1611 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02389 5182 1613 1612 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02390 1613 1612 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02391 21 2675 1612 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02392 19 2675 1613 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02393 5182 1615 1614 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02394 1615 1614 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02395 22 2669 1614 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02396 20 2669 1615 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02397 5182 1617 1616 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02398 1617 1616 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02399 21 2669 1616 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02400 19 2669 1617 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02401 5182 1619 1618 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02402 1619 1618 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02403 22 2671 1618 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02404 20 2671 1619 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02405 5182 1621 1620 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02406 1621 1620 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02407 21 2671 1620 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02408 19 2671 1621 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02409 5182 1623 1622 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02410 1623 1622 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02411 22 2673 1622 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02412 20 2673 1623 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02413 5182 1625 1624 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02414 1625 1624 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02415 21 2673 1624 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02416 19 2673 1625 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02417 5182 1627 1626 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02418 1627 1626 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02419 22 2691 1626 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02420 20 2691 1627 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02421 5182 1629 1628 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02422 1629 1628 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02423 21 2691 1628 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02424 19 2691 1629 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02425 5182 1631 1630 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02426 1631 1630 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02427 22 2685 1630 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02428 20 2685 1631 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02429 5182 1633 1632 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02430 1633 1632 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02431 21 2685 1632 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02432 19 2685 1633 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02433 5182 1635 1634 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02434 1635 1634 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02435 22 2687 1634 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02436 20 2687 1635 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02437 5182 1637 1636 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02438 1637 1636 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02439 21 2687 1636 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02440 19 2687 1637 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02441 5182 1639 1638 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02442 1639 1638 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02443 22 2689 1638 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02444 20 2689 1639 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02445 5182 1641 1640 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02446 1641 1640 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02447 21 2689 1640 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02448 19 2689 1641 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02449 5182 1643 1642 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02450 1643 1642 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02451 22 2707 1642 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02452 20 2707 1643 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02453 5182 1645 1644 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02454 1645 1644 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02455 21 2707 1644 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02456 19 2707 1645 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02457 5182 1647 1646 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02458 1647 1646 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02459 22 2701 1646 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02460 20 2701 1647 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02461 5182 1649 1648 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02462 1649 1648 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02463 21 2701 1648 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02464 19 2701 1649 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02465 5182 1651 1650 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02466 1651 1650 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02467 22 2703 1650 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02468 20 2703 1651 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02469 5182 1653 1652 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02470 1653 1652 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02471 21 2703 1652 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02472 19 2703 1653 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02473 5182 1655 1654 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02474 1655 1654 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02475 22 2705 1654 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02476 20 2705 1655 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02477 5182 1657 1656 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02478 1657 1656 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02479 21 2705 1656 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02480 19 2705 1657 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02481 5182 1659 1658 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02482 1659 1658 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02483 22 2723 1658 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02484 20 2723 1659 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02485 5182 1661 1660 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02486 1661 1660 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02487 21 2723 1660 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02488 19 2723 1661 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02489 5182 1663 1662 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02490 1663 1662 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02491 22 2717 1662 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02492 20 2717 1663 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02493 5182 1665 1664 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02494 1665 1664 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02495 21 2717 1664 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02496 19 2717 1665 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02497 5182 1667 1666 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02498 1667 1666 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02499 22 2719 1666 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02500 20 2719 1667 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02501 5182 1669 1668 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02502 1669 1668 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02503 21 2719 1668 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02504 19 2719 1669 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02505 5182 1671 1670 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02506 1671 1670 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02507 22 2721 1670 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02508 20 2721 1671 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02509 5182 1673 1672 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02510 1673 1672 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02511 21 2721 1672 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02512 19 2721 1673 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02513 5182 1675 1674 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02514 1675 1674 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02515 22 2739 1674 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02516 20 2739 1675 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02517 5182 1677 1676 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02518 1677 1676 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02519 21 2739 1676 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02520 19 2739 1677 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02521 5182 1679 1678 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02522 1679 1678 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02523 22 2733 1678 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02524 20 2733 1679 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02525 5182 1681 1680 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02526 1681 1680 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02527 21 2733 1680 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02528 19 2733 1681 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02529 5182 1683 1682 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02530 1683 1682 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02531 22 2735 1682 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02532 20 2735 1683 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02533 5182 1685 1684 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02534 1685 1684 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02535 21 2735 1684 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02536 19 2735 1685 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02537 5182 1687 1686 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02538 1687 1686 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02539 22 2737 1686 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02540 20 2737 1687 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02541 5182 1689 1688 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02542 1689 1688 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02543 21 2737 1688 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02544 19 2737 1689 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02545 5182 1691 1690 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02546 1691 1690 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02547 22 2755 1690 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02548 20 2755 1691 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02549 5182 1693 1692 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02550 1693 1692 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02551 21 2755 1692 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02552 19 2755 1693 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02553 5182 1695 1694 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02554 1695 1694 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02555 22 2749 1694 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02556 20 2749 1695 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02557 5182 1697 1696 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02558 1697 1696 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02559 21 2749 1696 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02560 19 2749 1697 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02561 5182 1699 1698 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02562 1699 1698 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02563 22 2751 1698 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02564 20 2751 1699 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02565 5182 1701 1700 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02566 1701 1700 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02567 21 2751 1700 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02568 19 2751 1701 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02569 5182 1703 1702 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02570 1703 1702 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02571 22 2753 1702 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02572 20 2753 1703 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02573 5182 1705 1704 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02574 1705 1704 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02575 21 2753 1704 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02576 19 2753 1705 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02577 5182 1707 1706 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02578 1707 1706 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02579 22 2771 1706 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02580 20 2771 1707 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02581 5182 1709 1708 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02582 1709 1708 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02583 21 2771 1708 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02584 19 2771 1709 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02585 5182 1711 1710 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02586 1711 1710 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02587 22 2765 1710 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02588 20 2765 1711 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02589 5182 1713 1712 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02590 1713 1712 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02591 21 2765 1712 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02592 19 2765 1713 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02593 5182 1715 1714 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02594 1715 1714 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02595 22 2767 1714 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02596 20 2767 1715 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02597 5182 1717 1716 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02598 1717 1716 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02599 21 2767 1716 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02600 19 2767 1717 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02601 5182 1719 1718 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02602 1719 1718 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02603 22 2769 1718 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02604 20 2769 1719 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02605 5182 1721 1720 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02606 1721 1720 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02607 21 2769 1720 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02608 19 2769 1721 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02609 5182 1723 1722 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02610 1723 1722 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02611 22 2787 1722 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02612 20 2787 1723 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02613 5182 1725 1724 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02614 1725 1724 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02615 21 2787 1724 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02616 19 2787 1725 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02617 5182 1727 1726 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02618 1727 1726 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02619 22 2781 1726 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02620 20 2781 1727 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02621 5182 1729 1728 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02622 1729 1728 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02623 21 2781 1728 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02624 19 2781 1729 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02625 5182 1731 1730 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02626 1731 1730 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02627 22 2783 1730 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02628 20 2783 1731 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02629 5182 1733 1732 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02630 1733 1732 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02631 21 2783 1732 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02632 19 2783 1733 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02633 5182 1735 1734 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02634 1735 1734 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02635 22 2785 1734 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02636 20 2785 1735 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02637 5182 1737 1736 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02638 1737 1736 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02639 21 2785 1736 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02640 19 2785 1737 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02641 5182 1739 1738 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02642 1739 1738 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02643 22 2803 1738 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02644 20 2803 1739 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02645 5182 1741 1740 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02646 1741 1740 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02647 21 2803 1740 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02648 19 2803 1741 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02649 5182 1743 1742 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02650 1743 1742 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02651 22 2797 1742 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02652 20 2797 1743 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02653 5182 1745 1744 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02654 1745 1744 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02655 21 2797 1744 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02656 19 2797 1745 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02657 5182 1747 1746 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02658 1747 1746 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02659 22 2799 1746 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02660 20 2799 1747 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02661 5182 1749 1748 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02662 1749 1748 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02663 21 2799 1748 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02664 19 2799 1749 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02665 5182 1751 1750 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02666 1751 1750 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02667 22 2801 1750 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02668 20 2801 1751 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02669 5182 1753 1752 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02670 1753 1752 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02671 21 2801 1752 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02672 19 2801 1753 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02673 5182 1755 1754 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02674 1755 1754 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02675 22 2819 1754 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02676 20 2819 1755 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02677 5182 1757 1756 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02678 1757 1756 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02679 21 2819 1756 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02680 19 2819 1757 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02681 5182 1759 1758 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02682 1759 1758 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02683 22 2813 1758 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02684 20 2813 1759 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02685 5182 1761 1760 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02686 1761 1760 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02687 21 2813 1760 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02688 19 2813 1761 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02689 5182 1763 1762 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02690 1763 1762 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02691 22 2815 1762 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02692 20 2815 1763 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02693 5182 1765 1764 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02694 1765 1764 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02695 21 2815 1764 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02696 19 2815 1765 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02697 5182 1767 1766 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02698 1767 1766 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02699 22 2817 1766 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02700 20 2817 1767 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02701 5182 1769 1768 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02702 1769 1768 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02703 21 2817 1768 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02704 19 2817 1769 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02705 5182 1771 1770 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02706 1771 1770 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02707 22 2835 1770 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02708 20 2835 1771 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02709 5182 1773 1772 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02710 1773 1772 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02711 21 2835 1772 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02712 19 2835 1773 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02713 5182 1775 1774 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02714 1775 1774 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02715 22 2829 1774 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02716 20 2829 1775 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02717 5182 1777 1776 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02718 1777 1776 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02719 21 2829 1776 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02720 19 2829 1777 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02721 5182 1779 1778 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02722 1779 1778 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02723 22 2831 1778 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02724 20 2831 1779 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02725 5182 1781 1780 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02726 1781 1780 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02727 21 2831 1780 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02728 19 2831 1781 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02729 5182 1783 1782 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02730 1783 1782 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02731 22 2833 1782 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02732 20 2833 1783 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02733 5182 1785 1784 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02734 1785 1784 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02735 21 2833 1784 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02736 19 2833 1785 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02737 5182 1787 1786 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02738 1787 1786 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02739 22 2851 1786 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02740 20 2851 1787 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02741 5182 1789 1788 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02742 1789 1788 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02743 21 2851 1788 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02744 19 2851 1789 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02745 5182 1791 1790 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02746 1791 1790 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02747 22 2845 1790 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02748 20 2845 1791 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02749 5182 1793 1792 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02750 1793 1792 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02751 21 2845 1792 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02752 19 2845 1793 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02753 5182 1795 1794 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02754 1795 1794 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02755 22 2847 1794 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02756 20 2847 1795 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02757 5182 1797 1796 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02758 1797 1796 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02759 21 2847 1796 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02760 19 2847 1797 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02761 5182 1799 1798 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02762 1799 1798 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02763 22 2849 1798 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02764 20 2849 1799 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02765 5182 1801 1800 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02766 1801 1800 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02767 21 2849 1800 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02768 19 2849 1801 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02769 5182 1803 1802 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02770 1803 1802 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02771 22 2867 1802 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02772 20 2867 1803 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02773 5182 1805 1804 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02774 1805 1804 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02775 21 2867 1804 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02776 19 2867 1805 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02777 5182 1807 1806 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02778 1807 1806 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02779 22 2861 1806 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02780 20 2861 1807 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02781 5182 1809 1808 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02782 1809 1808 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02783 21 2861 1808 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02784 19 2861 1809 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02785 5182 1811 1810 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02786 1811 1810 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02787 22 2863 1810 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02788 20 2863 1811 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02789 5182 1813 1812 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02790 1813 1812 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02791 21 2863 1812 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02792 19 2863 1813 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02793 5182 1815 1814 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02794 1815 1814 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02795 22 2865 1814 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02796 20 2865 1815 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02797 5182 1817 1816 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02798 1817 1816 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02799 21 2865 1816 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02800 19 2865 1817 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02801 5182 1819 1818 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02802 1819 1818 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02803 22 2883 1818 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02804 20 2883 1819 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02805 5182 1821 1820 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02806 1821 1820 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02807 21 2883 1820 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02808 19 2883 1821 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02809 5182 1823 1822 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02810 1823 1822 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02811 22 2877 1822 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02812 20 2877 1823 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02813 5182 1825 1824 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02814 1825 1824 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02815 21 2877 1824 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02816 19 2877 1825 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02817 5182 1827 1826 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02818 1827 1826 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02819 22 2879 1826 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02820 20 2879 1827 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02821 5182 1829 1828 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02822 1829 1828 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02823 21 2879 1828 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02824 19 2879 1829 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02825 5182 1831 1830 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02826 1831 1830 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02827 22 2881 1830 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02828 20 2881 1831 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02829 5182 1833 1832 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02830 1833 1832 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02831 21 2881 1832 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02832 19 2881 1833 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02833 5182 1835 1834 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02834 1835 1834 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02835 22 2899 1834 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02836 20 2899 1835 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02837 5182 1837 1836 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02838 1837 1836 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02839 21 2899 1836 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02840 19 2899 1837 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02841 5182 1839 1838 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02842 1839 1838 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02843 22 2893 1838 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02844 20 2893 1839 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02845 5182 1841 1840 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02846 1841 1840 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02847 21 2893 1840 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02848 19 2893 1841 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02849 5182 1843 1842 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02850 1843 1842 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02851 22 2895 1842 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02852 20 2895 1843 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02853 5182 1845 1844 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02854 1845 1844 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02855 21 2895 1844 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02856 19 2895 1845 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02857 5182 1847 1846 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02858 1847 1846 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02859 22 2897 1846 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02860 20 2897 1847 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02861 5182 1849 1848 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02862 1849 1848 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02863 21 2897 1848 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02864 19 2897 1849 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02865 5182 1851 1850 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02866 1851 1850 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02867 22 2915 1850 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02868 20 2915 1851 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02869 5182 1853 1852 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02870 1853 1852 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02871 21 2915 1852 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02872 19 2915 1853 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02873 5182 1855 1854 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02874 1855 1854 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02875 22 2909 1854 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02876 20 2909 1855 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02877 5182 1857 1856 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02878 1857 1856 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02879 21 2909 1856 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02880 19 2909 1857 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02881 5182 1859 1858 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02882 1859 1858 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02883 22 2911 1858 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02884 20 2911 1859 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02885 5182 1861 1860 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02886 1861 1860 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02887 21 2911 1860 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02888 19 2911 1861 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02889 5182 1863 1862 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02890 1863 1862 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02891 22 2913 1862 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02892 20 2913 1863 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02893 5182 1865 1864 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02894 1865 1864 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02895 21 2913 1864 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02896 19 2913 1865 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02897 5182 1867 1866 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02898 1867 1866 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02899 22 2931 1866 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02900 20 2931 1867 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02901 5182 1869 1868 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02902 1869 1868 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02903 21 2931 1868 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02904 19 2931 1869 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02905 5182 1871 1870 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02906 1871 1870 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02907 22 2925 1870 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02908 20 2925 1871 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02909 5182 1873 1872 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02910 1873 1872 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02911 21 2925 1872 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02912 19 2925 1873 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02913 5182 1875 1874 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02914 1875 1874 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02915 22 2927 1874 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02916 20 2927 1875 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02917 5182 1877 1876 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02918 1877 1876 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02919 21 2927 1876 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02920 19 2927 1877 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02921 5182 1879 1878 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02922 1879 1878 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02923 22 2929 1878 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02924 20 2929 1879 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02925 5182 1881 1880 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02926 1881 1880 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02927 21 2929 1880 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02928 19 2929 1881 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02929 5182 1883 1882 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02930 1883 1882 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02931 22 2947 1882 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02932 20 2947 1883 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02933 5182 1885 1884 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02934 1885 1884 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02935 21 2947 1884 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02936 19 2947 1885 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02937 5182 1887 1886 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02938 1887 1886 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02939 22 2941 1886 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02940 20 2941 1887 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02941 5182 1889 1888 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02942 1889 1888 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02943 21 2941 1888 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02944 19 2941 1889 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02945 5182 1891 1890 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02946 1891 1890 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02947 22 2943 1890 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02948 20 2943 1891 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02949 5182 1893 1892 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02950 1893 1892 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02951 21 2943 1892 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02952 19 2943 1893 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02953 5182 1895 1894 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02954 1895 1894 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02955 22 2945 1894 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02956 20 2945 1895 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02957 5182 1897 1896 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02958 1897 1896 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02959 21 2945 1896 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02960 19 2945 1897 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02961 5182 1899 1898 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02962 1899 1898 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02963 22 2963 1898 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02964 20 2963 1899 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02965 5182 1901 1900 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02966 1901 1900 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02967 21 2963 1900 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02968 19 2963 1901 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02969 5182 1903 1902 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02970 1903 1902 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02971 22 2957 1902 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02972 20 2957 1903 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02973 5182 1905 1904 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02974 1905 1904 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02975 21 2957 1904 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02976 19 2957 1905 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02977 5182 1907 1906 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02978 1907 1906 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02979 22 2959 1906 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02980 20 2959 1907 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02981 5182 1909 1908 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02982 1909 1908 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02983 21 2959 1908 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02984 19 2959 1909 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02985 5182 1911 1910 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02986 1911 1910 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02987 22 2961 1910 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02988 20 2961 1911 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02989 5182 1913 1912 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02990 1913 1912 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02991 21 2961 1912 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02992 19 2961 1913 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02993 5182 1915 1914 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02994 1915 1914 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02995 22 2979 1914 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02996 20 2979 1915 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02997 5182 1917 1916 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02998 1917 1916 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02999 21 2979 1916 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03000 19 2979 1917 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03001 5182 1919 1918 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03002 1919 1918 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03003 22 2973 1918 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03004 20 2973 1919 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03005 5182 1921 1920 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03006 1921 1920 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03007 21 2973 1920 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03008 19 2973 1921 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03009 5182 1923 1922 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03010 1923 1922 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03011 22 2975 1922 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03012 20 2975 1923 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03013 5182 1925 1924 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03014 1925 1924 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03015 21 2975 1924 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03016 19 2975 1925 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03017 5182 1927 1926 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03018 1927 1926 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03019 22 2977 1926 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03020 20 2977 1927 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03021 5182 1929 1928 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03022 1929 1928 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03023 21 2977 1928 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03024 19 2977 1929 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03025 5182 1931 1930 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03026 1931 1930 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03027 22 2995 1930 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03028 20 2995 1931 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03029 5182 1933 1932 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03030 1933 1932 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03031 21 2995 1932 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03032 19 2995 1933 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03033 5182 1935 1934 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03034 1935 1934 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03035 22 2989 1934 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03036 20 2989 1935 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03037 5182 1937 1936 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03038 1937 1936 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03039 21 2989 1936 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03040 19 2989 1937 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03041 5182 1939 1938 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03042 1939 1938 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03043 22 2991 1938 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03044 20 2991 1939 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03045 5182 1941 1940 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03046 1941 1940 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03047 21 2991 1940 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03048 19 2991 1941 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03049 5182 1943 1942 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03050 1943 1942 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03051 22 2993 1942 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03052 20 2993 1943 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03053 5182 1945 1944 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03054 1945 1944 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03055 21 2993 1944 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03056 19 2993 1945 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03057 5182 1947 1946 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03058 1947 1946 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03059 22 3011 1946 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03060 20 3011 1947 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03061 5182 1949 1948 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03062 1949 1948 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03063 21 3011 1948 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03064 19 3011 1949 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03065 5182 1951 1950 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03066 1951 1950 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03067 22 3005 1950 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03068 20 3005 1951 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03069 5182 1953 1952 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03070 1953 1952 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03071 21 3005 1952 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03072 19 3005 1953 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03073 5182 1955 1954 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03074 1955 1954 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03075 22 3007 1954 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03076 20 3007 1955 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03077 5182 1957 1956 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03078 1957 1956 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03079 21 3007 1956 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03080 19 3007 1957 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03081 5182 1959 1958 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03082 1959 1958 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03083 22 3009 1958 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03084 20 3009 1959 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03085 5182 1961 1960 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03086 1961 1960 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03087 21 3009 1960 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03088 19 3009 1961 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03089 5182 1963 1962 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03090 1963 1962 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03091 22 3027 1962 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03092 20 3027 1963 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03093 5182 1965 1964 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03094 1965 1964 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03095 21 3027 1964 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03096 19 3027 1965 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03097 5182 1967 1966 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03098 1967 1966 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03099 22 3021 1966 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03100 20 3021 1967 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03101 5182 1969 1968 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03102 1969 1968 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03103 21 3021 1968 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03104 19 3021 1969 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03105 5182 1971 1970 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03106 1971 1970 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03107 22 3023 1970 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03108 20 3023 1971 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03109 5182 1973 1972 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03110 1973 1972 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03111 21 3023 1972 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03112 19 3023 1973 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03113 5182 1975 1974 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03114 1975 1974 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03115 22 3025 1974 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03116 20 3025 1975 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03117 5182 1977 1976 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03118 1977 1976 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03119 21 3025 1976 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03120 19 3025 1977 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03121 5182 1979 1978 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03122 1979 1978 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03123 22 3043 1978 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03124 20 3043 1979 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03125 5182 1981 1980 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03126 1981 1980 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03127 21 3043 1980 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03128 19 3043 1981 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03129 5182 1983 1982 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03130 1983 1982 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03131 22 3037 1982 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03132 20 3037 1983 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03133 5182 1985 1984 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03134 1985 1984 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03135 21 3037 1984 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03136 19 3037 1985 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03137 5182 1987 1986 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03138 1987 1986 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03139 22 3039 1986 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03140 20 3039 1987 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03141 5182 1989 1988 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03142 1989 1988 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03143 21 3039 1988 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03144 19 3039 1989 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03145 5182 1991 1990 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03146 1991 1990 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03147 22 3041 1990 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03148 20 3041 1991 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03149 5182 1993 1992 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03150 1993 1992 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03151 21 3041 1992 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03152 19 3041 1993 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03153 19 3045 26 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_03154 26 3046 20 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_03155 21 3045 27 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_03156 27 3046 22 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_03157 1997 3083 1995 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03158 2002 1997 23 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03159 23 3074 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03160 23 1995 1994 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03161 5182 3074 24 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03162 1996 27 24 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03163 24 26 1995 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03164 1997 27 25 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03165 25 3074 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03166 25 26 1998 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03167 5183 3083 27 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03168 27 3083 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03169 5183 3083 26 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03170 26 3083 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03171 1999 3077 27 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_03172 26 3077 2000 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_03173 27 3083 26 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_03174 5182 5190 1999 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_03175 2000 2001 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_03176 1999 5190 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_03177 5182 2001 2000 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_03178 5182 5190 2001 5182 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03179 5190 2003 5182 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03180 5182 2003 5190 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03181 5182 3077 2003 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03182 2003 2002 5182 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03183 2003 3074 2004 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03184 31 2529 29 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03185 31 2529 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03186 29 2529 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03187 30 2529 28 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03188 5183 2529 30 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03189 5183 2529 28 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03190 5182 2006 2005 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03191 2006 2005 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03192 31 2547 2005 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03193 29 2547 2006 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03194 5182 2008 2007 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03195 2008 2007 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03196 30 2547 2007 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03197 28 2547 2008 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03198 5182 2010 2009 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03199 2010 2009 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03200 31 2541 2009 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03201 29 2541 2010 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03202 5182 2012 2011 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03203 2012 2011 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03204 30 2541 2011 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03205 28 2541 2012 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03206 5182 2014 2013 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03207 2014 2013 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03208 31 2543 2013 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03209 29 2543 2014 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03210 5182 2016 2015 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03211 2016 2015 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03212 30 2543 2015 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03213 28 2543 2016 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03214 5182 2018 2017 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03215 2018 2017 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03216 31 2545 2017 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03217 29 2545 2018 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03218 5182 2020 2019 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03219 2020 2019 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03220 30 2545 2019 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03221 28 2545 2020 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03222 5182 2022 2021 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03223 2022 2021 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03224 31 2563 2021 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03225 29 2563 2022 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03226 5182 2024 2023 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03227 2024 2023 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03228 30 2563 2023 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03229 28 2563 2024 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03230 5182 2026 2025 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03231 2026 2025 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03232 31 2557 2025 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03233 29 2557 2026 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03234 5182 2028 2027 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03235 2028 2027 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03236 30 2557 2027 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03237 28 2557 2028 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03238 5182 2030 2029 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03239 2030 2029 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03240 31 2559 2029 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03241 29 2559 2030 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03242 5182 2032 2031 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03243 2032 2031 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03244 30 2559 2031 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03245 28 2559 2032 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03246 5182 2034 2033 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03247 2034 2033 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03248 31 2561 2033 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03249 29 2561 2034 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03250 5182 2036 2035 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03251 2036 2035 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03252 30 2561 2035 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03253 28 2561 2036 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03254 5182 2038 2037 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03255 2038 2037 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03256 31 2579 2037 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03257 29 2579 2038 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03258 5182 2040 2039 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03259 2040 2039 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03260 30 2579 2039 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03261 28 2579 2040 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03262 5182 2042 2041 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03263 2042 2041 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03264 31 2573 2041 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03265 29 2573 2042 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03266 5182 2044 2043 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03267 2044 2043 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03268 30 2573 2043 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03269 28 2573 2044 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03270 5182 2046 2045 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03271 2046 2045 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03272 31 2575 2045 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03273 29 2575 2046 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03274 5182 2048 2047 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03275 2048 2047 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03276 30 2575 2047 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03277 28 2575 2048 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03278 5182 2050 2049 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03279 2050 2049 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03280 31 2577 2049 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03281 29 2577 2050 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03282 5182 2052 2051 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03283 2052 2051 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03284 30 2577 2051 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03285 28 2577 2052 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03286 5182 2054 2053 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03287 2054 2053 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03288 31 2595 2053 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03289 29 2595 2054 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03290 5182 2056 2055 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03291 2056 2055 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03292 30 2595 2055 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03293 28 2595 2056 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03294 5182 2058 2057 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03295 2058 2057 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03296 31 2589 2057 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03297 29 2589 2058 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03298 5182 2060 2059 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03299 2060 2059 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03300 30 2589 2059 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03301 28 2589 2060 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03302 5182 2062 2061 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03303 2062 2061 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03304 31 2591 2061 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03305 29 2591 2062 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03306 5182 2064 2063 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03307 2064 2063 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03308 30 2591 2063 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03309 28 2591 2064 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03310 5182 2066 2065 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03311 2066 2065 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03312 31 2593 2065 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03313 29 2593 2066 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03314 5182 2068 2067 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03315 2068 2067 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03316 30 2593 2067 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03317 28 2593 2068 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03318 5182 2070 2069 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03319 2070 2069 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03320 31 2611 2069 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03321 29 2611 2070 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03322 5182 2072 2071 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03323 2072 2071 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03324 30 2611 2071 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03325 28 2611 2072 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03326 5182 2074 2073 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03327 2074 2073 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03328 31 2605 2073 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03329 29 2605 2074 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03330 5182 2076 2075 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03331 2076 2075 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03332 30 2605 2075 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03333 28 2605 2076 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03334 5182 2078 2077 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03335 2078 2077 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03336 31 2607 2077 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03337 29 2607 2078 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03338 5182 2080 2079 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03339 2080 2079 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03340 30 2607 2079 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03341 28 2607 2080 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03342 5182 2082 2081 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03343 2082 2081 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03344 31 2609 2081 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03345 29 2609 2082 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03346 5182 2084 2083 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03347 2084 2083 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03348 30 2609 2083 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03349 28 2609 2084 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03350 5182 2086 2085 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03351 2086 2085 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03352 31 2627 2085 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03353 29 2627 2086 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03354 5182 2088 2087 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03355 2088 2087 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03356 30 2627 2087 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03357 28 2627 2088 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03358 5182 2090 2089 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03359 2090 2089 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03360 31 2621 2089 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03361 29 2621 2090 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03362 5182 2092 2091 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03363 2092 2091 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03364 30 2621 2091 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03365 28 2621 2092 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03366 5182 2094 2093 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03367 2094 2093 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03368 31 2623 2093 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03369 29 2623 2094 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03370 5182 2096 2095 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03371 2096 2095 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03372 30 2623 2095 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03373 28 2623 2096 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03374 5182 2098 2097 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03375 2098 2097 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03376 31 2625 2097 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03377 29 2625 2098 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03378 5182 2100 2099 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03379 2100 2099 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03380 30 2625 2099 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03381 28 2625 2100 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03382 5182 2102 2101 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03383 2102 2101 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03384 31 2643 2101 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03385 29 2643 2102 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03386 5182 2104 2103 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03387 2104 2103 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03388 30 2643 2103 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03389 28 2643 2104 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03390 5182 2106 2105 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03391 2106 2105 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03392 31 2637 2105 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03393 29 2637 2106 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03394 5182 2108 2107 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03395 2108 2107 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03396 30 2637 2107 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03397 28 2637 2108 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03398 5182 2110 2109 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03399 2110 2109 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03400 31 2639 2109 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03401 29 2639 2110 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03402 5182 2112 2111 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03403 2112 2111 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03404 30 2639 2111 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03405 28 2639 2112 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03406 5182 2114 2113 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03407 2114 2113 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03408 31 2641 2113 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03409 29 2641 2114 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03410 5182 2116 2115 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03411 2116 2115 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03412 30 2641 2115 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03413 28 2641 2116 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03414 5182 2118 2117 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03415 2118 2117 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03416 31 2659 2117 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03417 29 2659 2118 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03418 5182 2120 2119 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03419 2120 2119 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03420 30 2659 2119 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03421 28 2659 2120 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03422 5182 2122 2121 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03423 2122 2121 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03424 31 2653 2121 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03425 29 2653 2122 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03426 5182 2124 2123 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03427 2124 2123 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03428 30 2653 2123 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03429 28 2653 2124 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03430 5182 2126 2125 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03431 2126 2125 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03432 31 2655 2125 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03433 29 2655 2126 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03434 5182 2128 2127 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03435 2128 2127 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03436 30 2655 2127 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03437 28 2655 2128 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03438 5182 2130 2129 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03439 2130 2129 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03440 31 2657 2129 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03441 29 2657 2130 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03442 5182 2132 2131 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03443 2132 2131 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03444 30 2657 2131 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03445 28 2657 2132 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03446 5182 2134 2133 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03447 2134 2133 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03448 31 2675 2133 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03449 29 2675 2134 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03450 5182 2136 2135 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03451 2136 2135 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03452 30 2675 2135 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03453 28 2675 2136 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03454 5182 2138 2137 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03455 2138 2137 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03456 31 2669 2137 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03457 29 2669 2138 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03458 5182 2140 2139 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03459 2140 2139 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03460 30 2669 2139 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03461 28 2669 2140 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03462 5182 2142 2141 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03463 2142 2141 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03464 31 2671 2141 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03465 29 2671 2142 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03466 5182 2144 2143 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03467 2144 2143 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03468 30 2671 2143 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03469 28 2671 2144 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03470 5182 2146 2145 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03471 2146 2145 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03472 31 2673 2145 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03473 29 2673 2146 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03474 5182 2148 2147 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03475 2148 2147 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03476 30 2673 2147 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03477 28 2673 2148 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03478 5182 2150 2149 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03479 2150 2149 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03480 31 2691 2149 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03481 29 2691 2150 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03482 5182 2152 2151 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03483 2152 2151 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03484 30 2691 2151 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03485 28 2691 2152 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03486 5182 2154 2153 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03487 2154 2153 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03488 31 2685 2153 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03489 29 2685 2154 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03490 5182 2156 2155 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03491 2156 2155 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03492 30 2685 2155 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03493 28 2685 2156 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03494 5182 2158 2157 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03495 2158 2157 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03496 31 2687 2157 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03497 29 2687 2158 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03498 5182 2160 2159 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03499 2160 2159 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03500 30 2687 2159 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03501 28 2687 2160 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03502 5182 2162 2161 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03503 2162 2161 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03504 31 2689 2161 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03505 29 2689 2162 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03506 5182 2164 2163 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03507 2164 2163 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03508 30 2689 2163 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03509 28 2689 2164 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03510 5182 2166 2165 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03511 2166 2165 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03512 31 2707 2165 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03513 29 2707 2166 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03514 5182 2168 2167 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03515 2168 2167 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03516 30 2707 2167 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03517 28 2707 2168 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03518 5182 2170 2169 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03519 2170 2169 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03520 31 2701 2169 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03521 29 2701 2170 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03522 5182 2172 2171 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03523 2172 2171 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03524 30 2701 2171 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03525 28 2701 2172 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03526 5182 2174 2173 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03527 2174 2173 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03528 31 2703 2173 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03529 29 2703 2174 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03530 5182 2176 2175 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03531 2176 2175 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03532 30 2703 2175 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03533 28 2703 2176 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03534 5182 2178 2177 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03535 2178 2177 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03536 31 2705 2177 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03537 29 2705 2178 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03538 5182 2180 2179 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03539 2180 2179 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03540 30 2705 2179 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03541 28 2705 2180 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03542 5182 2182 2181 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03543 2182 2181 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03544 31 2723 2181 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03545 29 2723 2182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03546 5182 2184 2183 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03547 2184 2183 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03548 30 2723 2183 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03549 28 2723 2184 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03550 5182 2186 2185 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03551 2186 2185 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03552 31 2717 2185 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03553 29 2717 2186 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03554 5182 2188 2187 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03555 2188 2187 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03556 30 2717 2187 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03557 28 2717 2188 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03558 5182 2190 2189 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03559 2190 2189 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03560 31 2719 2189 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03561 29 2719 2190 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03562 5182 2192 2191 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03563 2192 2191 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03564 30 2719 2191 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03565 28 2719 2192 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03566 5182 2194 2193 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03567 2194 2193 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03568 31 2721 2193 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03569 29 2721 2194 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03570 5182 2196 2195 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03571 2196 2195 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03572 30 2721 2195 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03573 28 2721 2196 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03574 5182 2198 2197 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03575 2198 2197 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03576 31 2739 2197 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03577 29 2739 2198 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03578 5182 2200 2199 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03579 2200 2199 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03580 30 2739 2199 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03581 28 2739 2200 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03582 5182 2202 2201 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03583 2202 2201 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03584 31 2733 2201 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03585 29 2733 2202 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03586 5182 2204 2203 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03587 2204 2203 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03588 30 2733 2203 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03589 28 2733 2204 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03590 5182 2206 2205 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03591 2206 2205 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03592 31 2735 2205 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03593 29 2735 2206 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03594 5182 2208 2207 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03595 2208 2207 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03596 30 2735 2207 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03597 28 2735 2208 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03598 5182 2210 2209 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03599 2210 2209 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03600 31 2737 2209 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03601 29 2737 2210 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03602 5182 2212 2211 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03603 2212 2211 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03604 30 2737 2211 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03605 28 2737 2212 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03606 5182 2214 2213 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03607 2214 2213 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03608 31 2755 2213 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03609 29 2755 2214 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03610 5182 2216 2215 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03611 2216 2215 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03612 30 2755 2215 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03613 28 2755 2216 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03614 5182 2218 2217 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03615 2218 2217 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03616 31 2749 2217 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03617 29 2749 2218 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03618 5182 2220 2219 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03619 2220 2219 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03620 30 2749 2219 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03621 28 2749 2220 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03622 5182 2222 2221 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03623 2222 2221 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03624 31 2751 2221 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03625 29 2751 2222 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03626 5182 2224 2223 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03627 2224 2223 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03628 30 2751 2223 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03629 28 2751 2224 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03630 5182 2226 2225 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03631 2226 2225 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03632 31 2753 2225 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03633 29 2753 2226 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03634 5182 2228 2227 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03635 2228 2227 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03636 30 2753 2227 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03637 28 2753 2228 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03638 5182 2230 2229 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03639 2230 2229 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03640 31 2771 2229 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03641 29 2771 2230 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03642 5182 2232 2231 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03643 2232 2231 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03644 30 2771 2231 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03645 28 2771 2232 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03646 5182 2234 2233 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03647 2234 2233 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03648 31 2765 2233 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03649 29 2765 2234 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03650 5182 2236 2235 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03651 2236 2235 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03652 30 2765 2235 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03653 28 2765 2236 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03654 5182 2238 2237 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03655 2238 2237 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03656 31 2767 2237 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03657 29 2767 2238 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03658 5182 2240 2239 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03659 2240 2239 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03660 30 2767 2239 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03661 28 2767 2240 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03662 5182 2242 2241 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03663 2242 2241 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03664 31 2769 2241 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03665 29 2769 2242 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03666 5182 2244 2243 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03667 2244 2243 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03668 30 2769 2243 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03669 28 2769 2244 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03670 5182 2246 2245 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03671 2246 2245 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03672 31 2787 2245 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03673 29 2787 2246 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03674 5182 2248 2247 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03675 2248 2247 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03676 30 2787 2247 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03677 28 2787 2248 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03678 5182 2250 2249 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03679 2250 2249 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03680 31 2781 2249 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03681 29 2781 2250 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03682 5182 2252 2251 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03683 2252 2251 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03684 30 2781 2251 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03685 28 2781 2252 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03686 5182 2254 2253 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03687 2254 2253 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03688 31 2783 2253 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03689 29 2783 2254 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03690 5182 2256 2255 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03691 2256 2255 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03692 30 2783 2255 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03693 28 2783 2256 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03694 5182 2258 2257 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03695 2258 2257 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03696 31 2785 2257 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03697 29 2785 2258 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03698 5182 2260 2259 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03699 2260 2259 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03700 30 2785 2259 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03701 28 2785 2260 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03702 5182 2262 2261 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03703 2262 2261 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03704 31 2803 2261 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03705 29 2803 2262 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03706 5182 2264 2263 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03707 2264 2263 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03708 30 2803 2263 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03709 28 2803 2264 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03710 5182 2266 2265 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03711 2266 2265 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03712 31 2797 2265 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03713 29 2797 2266 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03714 5182 2268 2267 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03715 2268 2267 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03716 30 2797 2267 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03717 28 2797 2268 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03718 5182 2270 2269 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03719 2270 2269 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03720 31 2799 2269 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03721 29 2799 2270 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03722 5182 2272 2271 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03723 2272 2271 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03724 30 2799 2271 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03725 28 2799 2272 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03726 5182 2274 2273 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03727 2274 2273 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03728 31 2801 2273 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03729 29 2801 2274 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03730 5182 2276 2275 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03731 2276 2275 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03732 30 2801 2275 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03733 28 2801 2276 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03734 5182 2278 2277 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03735 2278 2277 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03736 31 2819 2277 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03737 29 2819 2278 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03738 5182 2280 2279 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03739 2280 2279 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03740 30 2819 2279 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03741 28 2819 2280 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03742 5182 2282 2281 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03743 2282 2281 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03744 31 2813 2281 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03745 29 2813 2282 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03746 5182 2284 2283 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03747 2284 2283 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03748 30 2813 2283 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03749 28 2813 2284 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03750 5182 2286 2285 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03751 2286 2285 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03752 31 2815 2285 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03753 29 2815 2286 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03754 5182 2288 2287 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03755 2288 2287 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03756 30 2815 2287 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03757 28 2815 2288 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03758 5182 2290 2289 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03759 2290 2289 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03760 31 2817 2289 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03761 29 2817 2290 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03762 5182 2292 2291 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03763 2292 2291 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03764 30 2817 2291 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03765 28 2817 2292 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03766 5182 2294 2293 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03767 2294 2293 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03768 31 2835 2293 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03769 29 2835 2294 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03770 5182 2296 2295 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03771 2296 2295 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03772 30 2835 2295 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03773 28 2835 2296 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03774 5182 2298 2297 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03775 2298 2297 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03776 31 2829 2297 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03777 29 2829 2298 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03778 5182 2300 2299 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03779 2300 2299 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03780 30 2829 2299 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03781 28 2829 2300 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03782 5182 2302 2301 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03783 2302 2301 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03784 31 2831 2301 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03785 29 2831 2302 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03786 5182 2304 2303 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03787 2304 2303 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03788 30 2831 2303 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03789 28 2831 2304 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03790 5182 2306 2305 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03791 2306 2305 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03792 31 2833 2305 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03793 29 2833 2306 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03794 5182 2308 2307 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03795 2308 2307 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03796 30 2833 2307 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03797 28 2833 2308 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03798 5182 2310 2309 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03799 2310 2309 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03800 31 2851 2309 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03801 29 2851 2310 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03802 5182 2312 2311 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03803 2312 2311 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03804 30 2851 2311 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03805 28 2851 2312 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03806 5182 2314 2313 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03807 2314 2313 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03808 31 2845 2313 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03809 29 2845 2314 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03810 5182 2316 2315 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03811 2316 2315 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03812 30 2845 2315 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03813 28 2845 2316 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03814 5182 2318 2317 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03815 2318 2317 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03816 31 2847 2317 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03817 29 2847 2318 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03818 5182 2320 2319 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03819 2320 2319 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03820 30 2847 2319 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03821 28 2847 2320 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03822 5182 2322 2321 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03823 2322 2321 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03824 31 2849 2321 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03825 29 2849 2322 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03826 5182 2324 2323 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03827 2324 2323 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03828 30 2849 2323 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03829 28 2849 2324 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03830 5182 2326 2325 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03831 2326 2325 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03832 31 2867 2325 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03833 29 2867 2326 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03834 5182 2328 2327 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03835 2328 2327 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03836 30 2867 2327 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03837 28 2867 2328 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03838 5182 2330 2329 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03839 2330 2329 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03840 31 2861 2329 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03841 29 2861 2330 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03842 5182 2332 2331 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03843 2332 2331 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03844 30 2861 2331 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03845 28 2861 2332 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03846 5182 2334 2333 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03847 2334 2333 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03848 31 2863 2333 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03849 29 2863 2334 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03850 5182 2336 2335 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03851 2336 2335 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03852 30 2863 2335 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03853 28 2863 2336 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03854 5182 2338 2337 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03855 2338 2337 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03856 31 2865 2337 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03857 29 2865 2338 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03858 5182 2340 2339 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03859 2340 2339 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03860 30 2865 2339 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03861 28 2865 2340 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03862 5182 2342 2341 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03863 2342 2341 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03864 31 2883 2341 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03865 29 2883 2342 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03866 5182 2344 2343 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03867 2344 2343 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03868 30 2883 2343 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03869 28 2883 2344 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03870 5182 2346 2345 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03871 2346 2345 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03872 31 2877 2345 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03873 29 2877 2346 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03874 5182 2348 2347 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03875 2348 2347 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03876 30 2877 2347 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03877 28 2877 2348 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03878 5182 2350 2349 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03879 2350 2349 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03880 31 2879 2349 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03881 29 2879 2350 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03882 5182 2352 2351 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03883 2352 2351 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03884 30 2879 2351 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03885 28 2879 2352 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03886 5182 2354 2353 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03887 2354 2353 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03888 31 2881 2353 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03889 29 2881 2354 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03890 5182 2356 2355 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03891 2356 2355 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03892 30 2881 2355 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03893 28 2881 2356 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03894 5182 2358 2357 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03895 2358 2357 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03896 31 2899 2357 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03897 29 2899 2358 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03898 5182 2360 2359 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03899 2360 2359 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03900 30 2899 2359 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03901 28 2899 2360 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03902 5182 2362 2361 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03903 2362 2361 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03904 31 2893 2361 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03905 29 2893 2362 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03906 5182 2364 2363 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03907 2364 2363 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03908 30 2893 2363 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03909 28 2893 2364 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03910 5182 2366 2365 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03911 2366 2365 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03912 31 2895 2365 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03913 29 2895 2366 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03914 5182 2368 2367 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03915 2368 2367 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03916 30 2895 2367 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03917 28 2895 2368 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03918 5182 2370 2369 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03919 2370 2369 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03920 31 2897 2369 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03921 29 2897 2370 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03922 5182 2372 2371 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03923 2372 2371 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03924 30 2897 2371 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03925 28 2897 2372 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03926 5182 2374 2373 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03927 2374 2373 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03928 31 2915 2373 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03929 29 2915 2374 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03930 5182 2376 2375 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03931 2376 2375 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03932 30 2915 2375 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03933 28 2915 2376 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03934 5182 2378 2377 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03935 2378 2377 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03936 31 2909 2377 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03937 29 2909 2378 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03938 5182 2380 2379 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03939 2380 2379 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03940 30 2909 2379 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03941 28 2909 2380 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03942 5182 2382 2381 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03943 2382 2381 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03944 31 2911 2381 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03945 29 2911 2382 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03946 5182 2384 2383 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03947 2384 2383 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03948 30 2911 2383 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03949 28 2911 2384 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03950 5182 2386 2385 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03951 2386 2385 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03952 31 2913 2385 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03953 29 2913 2386 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03954 5182 2388 2387 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03955 2388 2387 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03956 30 2913 2387 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03957 28 2913 2388 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03958 5182 2390 2389 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03959 2390 2389 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03960 31 2931 2389 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03961 29 2931 2390 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03962 5182 2392 2391 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03963 2392 2391 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03964 30 2931 2391 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03965 28 2931 2392 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03966 5182 2394 2393 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03967 2394 2393 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03968 31 2925 2393 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03969 29 2925 2394 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03970 5182 2396 2395 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03971 2396 2395 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03972 30 2925 2395 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03973 28 2925 2396 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03974 5182 2398 2397 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03975 2398 2397 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03976 31 2927 2397 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03977 29 2927 2398 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03978 5182 2400 2399 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03979 2400 2399 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03980 30 2927 2399 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03981 28 2927 2400 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03982 5182 2402 2401 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03983 2402 2401 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03984 31 2929 2401 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03985 29 2929 2402 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03986 5182 2404 2403 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03987 2404 2403 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03988 30 2929 2403 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03989 28 2929 2404 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03990 5182 2406 2405 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03991 2406 2405 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03992 31 2947 2405 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03993 29 2947 2406 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03994 5182 2408 2407 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03995 2408 2407 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03996 30 2947 2407 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03997 28 2947 2408 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03998 5182 2410 2409 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03999 2410 2409 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04000 31 2941 2409 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04001 29 2941 2410 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04002 5182 2412 2411 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04003 2412 2411 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04004 30 2941 2411 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04005 28 2941 2412 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04006 5182 2414 2413 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04007 2414 2413 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04008 31 2943 2413 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04009 29 2943 2414 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04010 5182 2416 2415 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04011 2416 2415 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04012 30 2943 2415 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04013 28 2943 2416 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04014 5182 2418 2417 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04015 2418 2417 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04016 31 2945 2417 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04017 29 2945 2418 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04018 5182 2420 2419 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04019 2420 2419 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04020 30 2945 2419 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04021 28 2945 2420 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04022 5182 2422 2421 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04023 2422 2421 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04024 31 2963 2421 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04025 29 2963 2422 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04026 5182 2424 2423 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04027 2424 2423 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04028 30 2963 2423 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04029 28 2963 2424 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04030 5182 2426 2425 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04031 2426 2425 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04032 31 2957 2425 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04033 29 2957 2426 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04034 5182 2428 2427 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04035 2428 2427 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04036 30 2957 2427 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04037 28 2957 2428 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04038 5182 2430 2429 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04039 2430 2429 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04040 31 2959 2429 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04041 29 2959 2430 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04042 5182 2432 2431 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04043 2432 2431 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04044 30 2959 2431 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04045 28 2959 2432 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04046 5182 2434 2433 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04047 2434 2433 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04048 31 2961 2433 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04049 29 2961 2434 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04050 5182 2436 2435 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04051 2436 2435 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04052 30 2961 2435 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04053 28 2961 2436 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04054 5182 2438 2437 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04055 2438 2437 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04056 31 2979 2437 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04057 29 2979 2438 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04058 5182 2440 2439 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04059 2440 2439 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04060 30 2979 2439 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04061 28 2979 2440 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04062 5182 2442 2441 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04063 2442 2441 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04064 31 2973 2441 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04065 29 2973 2442 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04066 5182 2444 2443 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04067 2444 2443 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04068 30 2973 2443 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04069 28 2973 2444 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04070 5182 2446 2445 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04071 2446 2445 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04072 31 2975 2445 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04073 29 2975 2446 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04074 5182 2448 2447 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04075 2448 2447 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04076 30 2975 2447 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04077 28 2975 2448 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04078 5182 2450 2449 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04079 2450 2449 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04080 31 2977 2449 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04081 29 2977 2450 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04082 5182 2452 2451 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04083 2452 2451 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04084 30 2977 2451 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04085 28 2977 2452 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04086 5182 2454 2453 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04087 2454 2453 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04088 31 2995 2453 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04089 29 2995 2454 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04090 5182 2456 2455 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04091 2456 2455 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04092 30 2995 2455 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04093 28 2995 2456 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04094 5182 2458 2457 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04095 2458 2457 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04096 31 2989 2457 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04097 29 2989 2458 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04098 5182 2460 2459 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04099 2460 2459 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04100 30 2989 2459 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04101 28 2989 2460 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04102 5182 2462 2461 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04103 2462 2461 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04104 31 2991 2461 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04105 29 2991 2462 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04106 5182 2464 2463 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04107 2464 2463 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04108 30 2991 2463 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04109 28 2991 2464 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04110 5182 2466 2465 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04111 2466 2465 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04112 31 2993 2465 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04113 29 2993 2466 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04114 5182 2468 2467 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04115 2468 2467 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04116 30 2993 2467 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04117 28 2993 2468 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04118 5182 2470 2469 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04119 2470 2469 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04120 31 3011 2469 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04121 29 3011 2470 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04122 5182 2472 2471 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04123 2472 2471 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04124 30 3011 2471 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04125 28 3011 2472 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04126 5182 2474 2473 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04127 2474 2473 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04128 31 3005 2473 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04129 29 3005 2474 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04130 5182 2476 2475 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04131 2476 2475 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04132 30 3005 2475 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04133 28 3005 2476 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04134 5182 2478 2477 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04135 2478 2477 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04136 31 3007 2477 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04137 29 3007 2478 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04138 5182 2480 2479 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04139 2480 2479 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04140 30 3007 2479 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04141 28 3007 2480 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04142 5182 2482 2481 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04143 2482 2481 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04144 31 3009 2481 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04145 29 3009 2482 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04146 5182 2484 2483 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04147 2484 2483 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04148 30 3009 2483 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04149 28 3009 2484 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04150 5182 2486 2485 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04151 2486 2485 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04152 31 3027 2485 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04153 29 3027 2486 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04154 5182 2488 2487 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04155 2488 2487 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04156 30 3027 2487 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04157 28 3027 2488 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04158 5182 2490 2489 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04159 2490 2489 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04160 31 3021 2489 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04161 29 3021 2490 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04162 5182 2492 2491 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04163 2492 2491 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04164 30 3021 2491 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04165 28 3021 2492 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04166 5182 2494 2493 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04167 2494 2493 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04168 31 3023 2493 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04169 29 3023 2494 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04170 5182 2496 2495 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04171 2496 2495 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04172 30 3023 2495 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04173 28 3023 2496 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04174 5182 2498 2497 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04175 2498 2497 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04176 31 3025 2497 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04177 29 3025 2498 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04178 5182 2500 2499 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04179 2500 2499 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04180 30 3025 2499 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04181 28 3025 2500 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04182 5182 2502 2501 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04183 2502 2501 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04184 31 3043 2501 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04185 29 3043 2502 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04186 5182 2504 2503 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04187 2504 2503 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04188 30 3043 2503 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04189 28 3043 2504 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04190 5182 2506 2505 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04191 2506 2505 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04192 31 3037 2505 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04193 29 3037 2506 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04194 5182 2508 2507 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04195 2508 2507 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04196 30 3037 2507 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04197 28 3037 2508 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04198 5182 2510 2509 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04199 2510 2509 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04200 31 3039 2509 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04201 29 3039 2510 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04202 5182 2512 2511 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04203 2512 2511 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04204 30 3039 2511 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04205 28 3039 2512 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04206 5182 2514 2513 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04207 2514 2513 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04208 31 3041 2513 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04209 29 3041 2514 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04210 5182 2516 2515 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04211 2516 2515 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04212 30 3041 2515 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04213 28 3041 2516 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04214 28 3045 35 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04215 35 3046 29 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04216 30 3045 36 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04217 36 3046 31 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04218 2520 3083 2518 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04219 2525 2520 32 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_04220 32 3074 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_04221 32 2518 2517 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_04222 5182 3074 33 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_04223 2519 36 33 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_04224 33 35 2518 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_04225 2520 36 34 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_04226 34 3074 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_04227 34 35 2521 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_04228 5183 3083 36 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04229 36 3083 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04230 5183 3083 35 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04231 35 3083 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04232 2522 3077 36 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_04233 35 3077 2523 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_04234 36 3083 35 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_04235 5182 5189 2522 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_04236 2523 2524 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_04237 2522 5189 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_04238 5182 2524 2523 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_04239 5182 5189 2524 5182 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_04240 5189 2526 5182 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04241 5182 2526 5189 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04242 5182 3077 2526 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_04243 2526 2525 5182 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_04244 2526 3074 2527 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_04245 2528 2530 5182 5182 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_04246 5182 2530 2528 5182 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_04247 2528 2530 5182 5182 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_04248 5182 2530 2528 5182 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_04249 2529 2532 5182 5182 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_04250 5182 2532 2529 5182 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_04251 2529 2532 5182 5182 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_04252 5182 2532 2529 5182 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_04253 5182 3085 2531 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04254 37 2531 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04255 2530 3086 37 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04256 38 2531 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04257 2532 3086 38 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04258 39 3064 40 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04259 5182 2537 39 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04260 40 3085 2546 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04261 41 3085 2544 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04262 5182 2537 42 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04263 42 3068 41 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04264 43 2537 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04265 2542 3085 44 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04266 44 3067 43 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04267 45 2537 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04268 2548 3085 46 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04269 46 3071 45 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04270 2537 2540 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04271 5182 2539 2537 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04272 2536 2548 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04273 2534 2542 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04274 5182 2542 2534 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04275 2535 2544 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04276 5182 2544 2535 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04277 5182 2546 2533 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04278 2533 2546 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04279 5182 2548 2536 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04280 47 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04281 2539 3057 47 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04282 5182 3048 49 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04283 48 3054 2540 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04284 49 3051 48 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04285 2543 2544 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04286 5182 2544 2543 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04287 2545 2546 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04288 5182 2546 2545 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04289 2547 2548 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04290 5182 2548 2547 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04291 2541 2542 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04292 5182 2542 2541 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04293 50 3064 51 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04294 5182 2553 50 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04295 51 3085 2562 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04296 52 3085 2560 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04297 5182 2553 53 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04298 53 3068 52 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04299 54 2553 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04300 2558 3085 55 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04301 55 3067 54 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04302 56 2553 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04303 2564 3085 57 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04304 57 3071 56 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04305 2553 2556 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04306 5182 2555 2553 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04307 2552 2564 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04308 2550 2558 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04309 5182 2558 2550 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04310 2551 2560 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04311 5182 2560 2551 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04312 5182 2562 2549 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04313 2549 2562 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04314 5182 2564 2552 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04315 58 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04316 2555 3057 58 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04317 5182 3047 60 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04318 59 3054 2556 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04319 60 3051 59 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04320 2559 2560 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04321 5182 2560 2559 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04322 2561 2562 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04323 5182 2562 2561 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04324 2563 2564 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04325 5182 2564 2563 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04326 2557 2558 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04327 5182 2558 2557 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04328 61 3064 62 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04329 5182 2569 61 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04330 62 3085 2578 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04331 63 3085 2576 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04332 5182 2569 64 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04333 64 3068 63 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04334 65 2569 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04335 2574 3085 66 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04336 66 3067 65 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04337 67 2569 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04338 2580 3085 68 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04339 68 3071 67 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04340 2569 2572 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04341 5182 2571 2569 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04342 2568 2580 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04343 2566 2574 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04344 5182 2574 2566 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04345 2567 2576 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04346 5182 2576 2567 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04347 5182 2578 2565 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04348 2565 2578 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04349 5182 2580 2568 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04350 69 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04351 2571 3057 69 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04352 5182 3048 71 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04353 70 3054 2572 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04354 71 3050 70 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04355 2575 2576 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04356 5182 2576 2575 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04357 2577 2578 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04358 5182 2578 2577 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04359 2579 2580 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04360 5182 2580 2579 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04361 2573 2574 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04362 5182 2574 2573 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04363 72 3064 73 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04364 5182 2585 72 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04365 73 3085 2594 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04366 74 3085 2592 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04367 5182 2585 75 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04368 75 3068 74 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04369 76 2585 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04370 2590 3085 77 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04371 77 3067 76 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04372 78 2585 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04373 2596 3085 79 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04374 79 3071 78 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04375 2585 2588 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04376 5182 2587 2585 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04377 2584 2596 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04378 2582 2590 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04379 5182 2590 2582 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04380 2583 2592 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04381 5182 2592 2583 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04382 5182 2594 2581 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04383 2581 2594 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04384 5182 2596 2584 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04385 80 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04386 2587 3057 80 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04387 5182 3047 82 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04388 81 3054 2588 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04389 82 3050 81 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04390 2591 2592 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04391 5182 2592 2591 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04392 2593 2594 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04393 5182 2594 2593 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04394 2595 2596 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04395 5182 2596 2595 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04396 2589 2590 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04397 5182 2590 2589 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04398 83 3064 84 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04399 5182 2601 83 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04400 84 3085 2610 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04401 85 3085 2608 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04402 5182 2601 86 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04403 86 3068 85 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04404 87 2601 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04405 2606 3085 88 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04406 88 3067 87 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04407 89 2601 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04408 2612 3085 90 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04409 90 3071 89 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04410 2601 2604 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04411 5182 2603 2601 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04412 2600 2612 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04413 2598 2606 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04414 5182 2606 2598 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04415 2599 2608 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04416 5182 2608 2599 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04417 5182 2610 2597 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04418 2597 2610 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04419 5182 2612 2600 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04420 91 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04421 2603 3057 91 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04422 5182 3048 93 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04423 92 3053 2604 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04424 93 3051 92 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04425 2607 2608 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04426 5182 2608 2607 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04427 2609 2610 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04428 5182 2610 2609 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04429 2611 2612 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04430 5182 2612 2611 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04431 2605 2606 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04432 5182 2606 2605 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04433 94 3064 95 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04434 5182 2617 94 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04435 95 3085 2626 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04436 96 3085 2624 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04437 5182 2617 97 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04438 97 3068 96 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04439 98 2617 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04440 2622 3085 99 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04441 99 3067 98 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04442 100 2617 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04443 2628 3085 101 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04444 101 3071 100 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04445 2617 2620 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04446 5182 2619 2617 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04447 2616 2628 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04448 2614 2622 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04449 5182 2622 2614 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04450 2615 2624 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04451 5182 2624 2615 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04452 5182 2626 2613 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04453 2613 2626 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04454 5182 2628 2616 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04455 102 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04456 2619 3057 102 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04457 5182 3047 104 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04458 103 3053 2620 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04459 104 3051 103 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04460 2623 2624 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04461 5182 2624 2623 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04462 2625 2626 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04463 5182 2626 2625 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04464 2627 2628 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04465 5182 2628 2627 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04466 2621 2622 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04467 5182 2622 2621 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04468 105 3064 106 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04469 5182 2633 105 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04470 106 3085 2642 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04471 107 3085 2640 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04472 5182 2633 108 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04473 108 3068 107 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04474 109 2633 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04475 2638 3085 110 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04476 110 3067 109 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04477 111 2633 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04478 2644 3085 112 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04479 112 3071 111 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04480 2633 2636 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04481 5182 2635 2633 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04482 2632 2644 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04483 2630 2638 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04484 5182 2638 2630 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04485 2631 2640 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04486 5182 2640 2631 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04487 5182 2642 2629 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04488 2629 2642 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04489 5182 2644 2632 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04490 113 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04491 2635 3057 113 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04492 5182 3048 115 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04493 114 3053 2636 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04494 115 3050 114 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04495 2639 2640 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04496 5182 2640 2639 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04497 2641 2642 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04498 5182 2642 2641 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04499 2643 2644 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04500 5182 2644 2643 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04501 2637 2638 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04502 5182 2638 2637 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04503 116 3064 117 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04504 5182 2649 116 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04505 117 3085 2658 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04506 118 3085 2656 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04507 5182 2649 119 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04508 119 3068 118 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04509 120 2649 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04510 2654 3085 121 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04511 121 3067 120 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04512 122 2649 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04513 2660 3085 123 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04514 123 3071 122 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04515 2649 2652 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04516 5182 2651 2649 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04517 2648 2660 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04518 2646 2654 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04519 5182 2654 2646 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04520 2647 2656 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04521 5182 2656 2647 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04522 5182 2658 2645 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04523 2645 2658 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04524 5182 2660 2648 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04525 124 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04526 2651 3057 124 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04527 5182 3047 126 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04528 125 3053 2652 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04529 126 3050 125 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04530 2655 2656 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04531 5182 2656 2655 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04532 2657 2658 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04533 5182 2658 2657 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04534 2659 2660 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04535 5182 2660 2659 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04536 2653 2654 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04537 5182 2654 2653 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04538 127 3064 128 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04539 5182 2665 127 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04540 128 3085 2674 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04541 129 3085 2672 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04542 5182 2665 130 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04543 130 3068 129 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04544 131 2665 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04545 2670 3085 132 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04546 132 3067 131 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04547 133 2665 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04548 2676 3085 134 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04549 134 3071 133 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04550 2665 2668 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04551 5182 2667 2665 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04552 2664 2676 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04553 2662 2670 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04554 5182 2670 2662 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04555 2663 2672 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04556 5182 2672 2663 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04557 5182 2674 2661 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04558 2661 2674 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04559 5182 2676 2664 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04560 135 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04561 2667 3056 135 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04562 5182 3048 137 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04563 136 3054 2668 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04564 137 3051 136 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04565 2671 2672 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04566 5182 2672 2671 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04567 2673 2674 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04568 5182 2674 2673 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04569 2675 2676 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04570 5182 2676 2675 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04571 2669 2670 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04572 5182 2670 2669 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04573 138 3064 139 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04574 5182 2681 138 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04575 139 3085 2690 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04576 140 3085 2688 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04577 5182 2681 141 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04578 141 3068 140 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04579 142 2681 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04580 2686 3085 143 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04581 143 3067 142 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04582 144 2681 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04583 2692 3085 145 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04584 145 3071 144 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04585 2681 2684 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04586 5182 2683 2681 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04587 2680 2692 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04588 2678 2686 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04589 5182 2686 2678 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04590 2679 2688 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04591 5182 2688 2679 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04592 5182 2690 2677 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04593 2677 2690 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04594 5182 2692 2680 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04595 146 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04596 2683 3056 146 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04597 5182 3047 148 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04598 147 3054 2684 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04599 148 3051 147 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04600 2687 2688 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04601 5182 2688 2687 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04602 2689 2690 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04603 5182 2690 2689 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04604 2691 2692 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04605 5182 2692 2691 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04606 2685 2686 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04607 5182 2686 2685 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04608 149 3064 150 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04609 5182 2697 149 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04610 150 3085 2706 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04611 151 3085 2704 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04612 5182 2697 152 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04613 152 3068 151 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04614 153 2697 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04615 2702 3085 154 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04616 154 3067 153 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04617 155 2697 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04618 2708 3085 156 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04619 156 3071 155 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04620 2697 2700 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04621 5182 2699 2697 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04622 2696 2708 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04623 2694 2702 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04624 5182 2702 2694 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04625 2695 2704 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04626 5182 2704 2695 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04627 5182 2706 2693 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04628 2693 2706 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04629 5182 2708 2696 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04630 157 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04631 2699 3056 157 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04632 5182 3048 159 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04633 158 3054 2700 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04634 159 3050 158 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04635 2703 2704 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04636 5182 2704 2703 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04637 2705 2706 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04638 5182 2706 2705 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04639 2707 2708 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04640 5182 2708 2707 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04641 2701 2702 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04642 5182 2702 2701 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04643 160 3064 161 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04644 5182 2713 160 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04645 161 3085 2722 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04646 162 3085 2720 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04647 5182 2713 163 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04648 163 3068 162 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04649 164 2713 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04650 2718 3085 165 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04651 165 3067 164 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04652 166 2713 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04653 2724 3085 167 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04654 167 3071 166 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04655 2713 2716 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04656 5182 2715 2713 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04657 2712 2724 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04658 2710 2718 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04659 5182 2718 2710 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04660 2711 2720 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04661 5182 2720 2711 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04662 5182 2722 2709 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04663 2709 2722 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04664 5182 2724 2712 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04665 168 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04666 2715 3056 168 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04667 5182 3047 170 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04668 169 3054 2716 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04669 170 3050 169 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04670 2719 2720 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04671 5182 2720 2719 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04672 2721 2722 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04673 5182 2722 2721 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04674 2723 2724 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04675 5182 2724 2723 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04676 2717 2718 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04677 5182 2718 2717 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04678 171 3064 172 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04679 5182 2729 171 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04680 172 3085 2738 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04681 173 3085 2736 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04682 5182 2729 174 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04683 174 3068 173 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04684 175 2729 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04685 2734 3085 176 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04686 176 3067 175 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04687 177 2729 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04688 2740 3085 178 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04689 178 3071 177 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04690 2729 2732 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04691 5182 2731 2729 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04692 2728 2740 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04693 2726 2734 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04694 5182 2734 2726 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04695 2727 2736 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04696 5182 2736 2727 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04697 5182 2738 2725 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04698 2725 2738 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04699 5182 2740 2728 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04700 179 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04701 2731 3056 179 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04702 5182 3048 181 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04703 180 3053 2732 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04704 181 3051 180 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04705 2735 2736 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04706 5182 2736 2735 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04707 2737 2738 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04708 5182 2738 2737 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04709 2739 2740 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04710 5182 2740 2739 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04711 2733 2734 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04712 5182 2734 2733 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04713 182 3064 183 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04714 5182 2745 182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04715 183 3085 2754 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04716 184 3085 2752 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04717 5182 2745 185 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04718 185 3068 184 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04719 186 2745 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04720 2750 3085 187 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04721 187 3067 186 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04722 188 2745 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04723 2756 3085 189 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04724 189 3071 188 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04725 2745 2748 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04726 5182 2747 2745 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04727 2744 2756 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04728 2742 2750 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04729 5182 2750 2742 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04730 2743 2752 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04731 5182 2752 2743 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04732 5182 2754 2741 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04733 2741 2754 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04734 5182 2756 2744 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04735 190 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04736 2747 3056 190 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04737 5182 3047 192 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04738 191 3053 2748 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04739 192 3051 191 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04740 2751 2752 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04741 5182 2752 2751 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04742 2753 2754 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04743 5182 2754 2753 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04744 2755 2756 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04745 5182 2756 2755 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04746 2749 2750 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04747 5182 2750 2749 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04748 193 3064 194 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04749 5182 2761 193 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04750 194 3085 2770 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04751 195 3085 2768 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04752 5182 2761 196 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04753 196 3068 195 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04754 197 2761 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04755 2766 3085 198 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04756 198 3067 197 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04757 199 2761 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04758 2772 3085 200 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04759 200 3071 199 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04760 2761 2764 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04761 5182 2763 2761 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04762 2760 2772 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04763 2758 2766 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04764 5182 2766 2758 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04765 2759 2768 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04766 5182 2768 2759 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04767 5182 2770 2757 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04768 2757 2770 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04769 5182 2772 2760 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04770 201 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04771 2763 3056 201 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04772 5182 3048 203 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04773 202 3053 2764 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04774 203 3050 202 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04775 2767 2768 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04776 5182 2768 2767 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04777 2769 2770 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04778 5182 2770 2769 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04779 2771 2772 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04780 5182 2772 2771 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04781 2765 2766 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04782 5182 2766 2765 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04783 204 3064 205 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04784 5182 2777 204 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04785 205 3085 2786 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04786 206 3085 2784 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04787 5182 2777 207 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04788 207 3068 206 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04789 208 2777 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04790 2782 3085 209 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04791 209 3067 208 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04792 210 2777 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04793 2788 3085 211 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04794 211 3071 210 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04795 2777 2780 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04796 5182 2779 2777 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04797 2776 2788 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04798 2774 2782 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04799 5182 2782 2774 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04800 2775 2784 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04801 5182 2784 2775 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04802 5182 2786 2773 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04803 2773 2786 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04804 5182 2788 2776 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04805 212 3060 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04806 2779 3056 212 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04807 5182 3047 214 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04808 213 3053 2780 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04809 214 3050 213 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04810 2783 2784 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04811 5182 2784 2783 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04812 2785 2786 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04813 5182 2786 2785 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04814 2787 2788 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04815 5182 2788 2787 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04816 2781 2782 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04817 5182 2782 2781 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04818 215 3064 216 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04819 5182 2793 215 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04820 216 3085 2802 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04821 217 3085 2800 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04822 5182 2793 218 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04823 218 3068 217 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04824 219 2793 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04825 2798 3085 220 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04826 220 3067 219 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04827 221 2793 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04828 2804 3085 222 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04829 222 3071 221 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04830 2793 2796 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04831 5182 2795 2793 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04832 2792 2804 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04833 2790 2798 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04834 5182 2798 2790 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04835 2791 2800 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04836 5182 2800 2791 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04837 5182 2802 2789 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04838 2789 2802 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04839 5182 2804 2792 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04840 223 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04841 2795 3057 223 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04842 5182 3048 225 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04843 224 3054 2796 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04844 225 3051 224 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04845 2799 2800 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04846 5182 2800 2799 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04847 2801 2802 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04848 5182 2802 2801 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04849 2803 2804 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04850 5182 2804 2803 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04851 2797 2798 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04852 5182 2798 2797 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04853 226 3064 227 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04854 5182 2809 226 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04855 227 3085 2818 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04856 228 3085 2816 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04857 5182 2809 229 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04858 229 3068 228 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04859 230 2809 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04860 2814 3085 231 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04861 231 3067 230 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04862 232 2809 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04863 2820 3085 233 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04864 233 3071 232 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04865 2809 2812 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04866 5182 2811 2809 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04867 2808 2820 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04868 2806 2814 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04869 5182 2814 2806 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04870 2807 2816 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04871 5182 2816 2807 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04872 5182 2818 2805 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04873 2805 2818 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04874 5182 2820 2808 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04875 234 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04876 2811 3057 234 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04877 5182 3047 236 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04878 235 3054 2812 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04879 236 3051 235 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04880 2815 2816 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04881 5182 2816 2815 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04882 2817 2818 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04883 5182 2818 2817 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04884 2819 2820 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04885 5182 2820 2819 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04886 2813 2814 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04887 5182 2814 2813 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04888 237 3064 238 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04889 5182 2825 237 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04890 238 3085 2834 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04891 239 3085 2832 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04892 5182 2825 240 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04893 240 3068 239 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04894 241 2825 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04895 2830 3085 242 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04896 242 3067 241 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04897 243 2825 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04898 2836 3085 244 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04899 244 3071 243 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04900 2825 2828 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04901 5182 2827 2825 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04902 2824 2836 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04903 2822 2830 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04904 5182 2830 2822 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04905 2823 2832 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04906 5182 2832 2823 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04907 5182 2834 2821 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04908 2821 2834 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04909 5182 2836 2824 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04910 245 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04911 2827 3057 245 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04912 5182 3048 247 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04913 246 3054 2828 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04914 247 3050 246 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04915 2831 2832 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04916 5182 2832 2831 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04917 2833 2834 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04918 5182 2834 2833 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04919 2835 2836 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04920 5182 2836 2835 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04921 2829 2830 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04922 5182 2830 2829 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04923 248 3064 249 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04924 5182 2841 248 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04925 249 3085 2850 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04926 250 3085 2848 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04927 5182 2841 251 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04928 251 3068 250 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04929 252 2841 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04930 2846 3085 253 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04931 253 3067 252 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04932 254 2841 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04933 2852 3085 255 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04934 255 3071 254 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04935 2841 2844 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04936 5182 2843 2841 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04937 2840 2852 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04938 2838 2846 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04939 5182 2846 2838 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04940 2839 2848 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04941 5182 2848 2839 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04942 5182 2850 2837 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04943 2837 2850 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04944 5182 2852 2840 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04945 256 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04946 2843 3057 256 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04947 5182 3047 258 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04948 257 3054 2844 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04949 258 3050 257 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04950 2847 2848 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04951 5182 2848 2847 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04952 2849 2850 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04953 5182 2850 2849 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04954 2851 2852 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04955 5182 2852 2851 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04956 2845 2846 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04957 5182 2846 2845 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04958 259 3064 260 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04959 5182 2857 259 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04960 260 3085 2866 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04961 261 3085 2864 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04962 5182 2857 262 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04963 262 3068 261 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04964 263 2857 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04965 2862 3085 264 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04966 264 3067 263 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04967 265 2857 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04968 2868 3085 266 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04969 266 3071 265 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04970 2857 2860 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04971 5182 2859 2857 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04972 2856 2868 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04973 2854 2862 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04974 5182 2862 2854 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04975 2855 2864 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04976 5182 2864 2855 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04977 5182 2866 2853 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04978 2853 2866 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04979 5182 2868 2856 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04980 267 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04981 2859 3057 267 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04982 5182 3048 269 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04983 268 3053 2860 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04984 269 3051 268 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04985 2863 2864 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04986 5182 2864 2863 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04987 2865 2866 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04988 5182 2866 2865 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04989 2867 2868 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04990 5182 2868 2867 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04991 2861 2862 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04992 5182 2862 2861 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_04993 270 3064 271 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04994 5182 2873 270 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04995 271 3085 2882 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04996 272 3085 2880 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04997 5182 2873 273 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04998 273 3068 272 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_04999 274 2873 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05000 2878 3085 275 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05001 275 3067 274 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05002 276 2873 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05003 2884 3085 277 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05004 277 3071 276 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05005 2873 2876 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05006 5182 2875 2873 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05007 2872 2884 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05008 2870 2878 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05009 5182 2878 2870 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05010 2871 2880 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05011 5182 2880 2871 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05012 5182 2882 2869 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05013 2869 2882 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05014 5182 2884 2872 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05015 278 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05016 2875 3057 278 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05017 5182 3047 280 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05018 279 3053 2876 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05019 280 3051 279 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05020 2879 2880 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05021 5182 2880 2879 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05022 2881 2882 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05023 5182 2882 2881 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05024 2883 2884 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05025 5182 2884 2883 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05026 2877 2878 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05027 5182 2878 2877 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05028 281 3064 282 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05029 5182 2889 281 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05030 282 3085 2898 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05031 283 3085 2896 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05032 5182 2889 284 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05033 284 3068 283 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05034 285 2889 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05035 2894 3085 286 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05036 286 3067 285 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05037 287 2889 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05038 2900 3085 288 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05039 288 3071 287 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05040 2889 2892 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05041 5182 2891 2889 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05042 2888 2900 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05043 2886 2894 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05044 5182 2894 2886 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05045 2887 2896 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05046 5182 2896 2887 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05047 5182 2898 2885 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05048 2885 2898 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05049 5182 2900 2888 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05050 289 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05051 2891 3057 289 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05052 5182 3048 291 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05053 290 3053 2892 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05054 291 3050 290 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05055 2895 2896 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05056 5182 2896 2895 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05057 2897 2898 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05058 5182 2898 2897 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05059 2899 2900 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05060 5182 2900 2899 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05061 2893 2894 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05062 5182 2894 2893 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05063 292 3064 293 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05064 5182 2905 292 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05065 293 3085 2914 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05066 294 3085 2912 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05067 5182 2905 295 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05068 295 3068 294 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05069 296 2905 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05070 2910 3085 297 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05071 297 3067 296 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05072 298 2905 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05073 2916 3085 299 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05074 299 3071 298 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05075 2905 2908 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05076 5182 2907 2905 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05077 2904 2916 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05078 2902 2910 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05079 5182 2910 2902 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05080 2903 2912 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05081 5182 2912 2903 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05082 5182 2914 2901 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05083 2901 2914 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05084 5182 2916 2904 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05085 300 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05086 2907 3057 300 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05087 5182 3047 302 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05088 301 3053 2908 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05089 302 3050 301 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05090 2911 2912 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05091 5182 2912 2911 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05092 2913 2914 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05093 5182 2914 2913 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05094 2915 2916 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05095 5182 2916 2915 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05096 2909 2910 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05097 5182 2910 2909 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05098 303 3064 304 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05099 5182 2921 303 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05100 304 3085 2930 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05101 305 3085 2928 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05102 5182 2921 306 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05103 306 3068 305 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05104 307 2921 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05105 2926 3085 308 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05106 308 3067 307 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05107 309 2921 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05108 2932 3085 310 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05109 310 3071 309 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05110 2921 2924 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05111 5182 2923 2921 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05112 2920 2932 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05113 2918 2926 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05114 5182 2926 2918 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05115 2919 2928 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05116 5182 2928 2919 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05117 5182 2930 2917 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05118 2917 2930 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05119 5182 2932 2920 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05120 311 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05121 2923 3056 311 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05122 5182 3048 313 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05123 312 3054 2924 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05124 313 3051 312 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05125 2927 2928 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05126 5182 2928 2927 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05127 2929 2930 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05128 5182 2930 2929 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05129 2931 2932 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05130 5182 2932 2931 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05131 2925 2926 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05132 5182 2926 2925 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05133 314 3064 315 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05134 5182 2937 314 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05135 315 3085 2946 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05136 316 3085 2944 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05137 5182 2937 317 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05138 317 3068 316 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05139 318 2937 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05140 2942 3085 319 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05141 319 3067 318 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05142 320 2937 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05143 2948 3085 321 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05144 321 3071 320 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05145 2937 2940 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05146 5182 2939 2937 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05147 2936 2948 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05148 2934 2942 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05149 5182 2942 2934 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05150 2935 2944 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05151 5182 2944 2935 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05152 5182 2946 2933 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05153 2933 2946 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05154 5182 2948 2936 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05155 322 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05156 2939 3056 322 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05157 5182 3047 324 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05158 323 3054 2940 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05159 324 3051 323 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05160 2943 2944 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05161 5182 2944 2943 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05162 2945 2946 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05163 5182 2946 2945 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05164 2947 2948 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05165 5182 2948 2947 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05166 2941 2942 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05167 5182 2942 2941 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05168 325 3064 326 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05169 5182 2953 325 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05170 326 3085 2962 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05171 327 3085 2960 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05172 5182 2953 328 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05173 328 3068 327 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05174 329 2953 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05175 2958 3085 330 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05176 330 3067 329 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05177 331 2953 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05178 2964 3085 332 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05179 332 3071 331 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05180 2953 2956 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05181 5182 2955 2953 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05182 2952 2964 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05183 2950 2958 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05184 5182 2958 2950 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05185 2951 2960 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05186 5182 2960 2951 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05187 5182 2962 2949 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05188 2949 2962 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05189 5182 2964 2952 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05190 333 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05191 2955 3056 333 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05192 5182 3048 335 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05193 334 3054 2956 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05194 335 3050 334 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05195 2959 2960 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05196 5182 2960 2959 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05197 2961 2962 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05198 5182 2962 2961 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05199 2963 2964 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05200 5182 2964 2963 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05201 2957 2958 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05202 5182 2958 2957 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05203 336 3064 337 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05204 5182 2969 336 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05205 337 3085 2978 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05206 338 3085 2976 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05207 5182 2969 339 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05208 339 3068 338 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05209 340 2969 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05210 2974 3085 341 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05211 341 3067 340 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05212 342 2969 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05213 2980 3085 343 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05214 343 3071 342 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05215 2969 2972 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05216 5182 2971 2969 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05217 2968 2980 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05218 2966 2974 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05219 5182 2974 2966 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05220 2967 2976 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05221 5182 2976 2967 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05222 5182 2978 2965 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05223 2965 2978 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05224 5182 2980 2968 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05225 344 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05226 2971 3056 344 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05227 5182 3047 346 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05228 345 3054 2972 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05229 346 3050 345 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05230 2975 2976 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05231 5182 2976 2975 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05232 2977 2978 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05233 5182 2978 2977 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05234 2979 2980 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05235 5182 2980 2979 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05236 2973 2974 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05237 5182 2974 2973 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05238 347 3064 348 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05239 5182 2985 347 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05240 348 3085 2994 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05241 349 3085 2992 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05242 5182 2985 350 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05243 350 3068 349 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05244 351 2985 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05245 2990 3085 352 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05246 352 3067 351 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05247 353 2985 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05248 2996 3085 354 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05249 354 3071 353 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05250 2985 2988 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05251 5182 2987 2985 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05252 2984 2996 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05253 2982 2990 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05254 5182 2990 2982 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05255 2983 2992 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05256 5182 2992 2983 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05257 5182 2994 2981 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05258 2981 2994 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05259 5182 2996 2984 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05260 355 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05261 2987 3056 355 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05262 5182 3048 357 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05263 356 3053 2988 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05264 357 3051 356 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05265 2991 2992 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05266 5182 2992 2991 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05267 2993 2994 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05268 5182 2994 2993 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05269 2995 2996 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05270 5182 2996 2995 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05271 2989 2990 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05272 5182 2990 2989 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05273 358 3064 359 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05274 5182 3001 358 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05275 359 3085 3010 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05276 360 3085 3008 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05277 5182 3001 361 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05278 361 3068 360 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05279 362 3001 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05280 3006 3085 363 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05281 363 3067 362 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05282 364 3001 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05283 3012 3085 365 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05284 365 3071 364 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05285 3001 3004 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05286 5182 3003 3001 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05287 3000 3012 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05288 2998 3006 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05289 5182 3006 2998 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05290 2999 3008 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05291 5182 3008 2999 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05292 5182 3010 2997 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05293 2997 3010 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05294 5182 3012 3000 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05295 366 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05296 3003 3056 366 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05297 5182 3047 368 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05298 367 3053 3004 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05299 368 3051 367 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05300 3007 3008 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05301 5182 3008 3007 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05302 3009 3010 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05303 5182 3010 3009 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05304 3011 3012 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05305 5182 3012 3011 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05306 3005 3006 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05307 5182 3006 3005 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05308 369 3064 370 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05309 5182 3017 369 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05310 370 3085 3026 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05311 371 3085 3024 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05312 5182 3017 372 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05313 372 3068 371 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05314 373 3017 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05315 3022 3085 374 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05316 374 3067 373 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05317 375 3017 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05318 3028 3085 376 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05319 376 3071 375 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05320 3017 3020 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05321 5182 3019 3017 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05322 3016 3028 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05323 3014 3022 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05324 5182 3022 3014 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05325 3015 3024 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05326 5182 3024 3015 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05327 5182 3026 3013 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05328 3013 3026 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05329 5182 3028 3016 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05330 377 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05331 3019 3056 377 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05332 5182 3048 379 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05333 378 3053 3020 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05334 379 3050 378 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05335 3023 3024 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05336 5182 3024 3023 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05337 3025 3026 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05338 5182 3026 3025 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05339 3027 3028 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05340 5182 3028 3027 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05341 3021 3022 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05342 5182 3022 3021 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05343 380 3064 381 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05344 5182 3033 380 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05345 381 3085 3042 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05346 382 3085 3040 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05347 5182 3033 383 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05348 383 3068 382 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05349 384 3033 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05350 3038 3085 385 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05351 385 3067 384 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05352 386 3033 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05353 3044 3085 387 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05354 387 3071 386 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05355 3033 3036 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05356 5182 3035 3033 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05357 3032 3044 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05358 3030 3038 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05359 5182 3038 3030 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05360 3031 3040 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05361 5182 3040 3031 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05362 5182 3042 3029 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05363 3029 3042 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05364 5182 3044 3032 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05365 388 3059 5182 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05366 3035 3056 388 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05367 5182 3047 390 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05368 389 3053 3036 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05369 390 3050 389 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05370 3039 3040 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05371 5182 3040 3039 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05372 3041 3042 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05373 5182 3042 3041 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05374 3043 3044 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05375 5182 3044 3043 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05376 3037 3038 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05377 5182 3038 3037 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05378 3046 3073 5182 5182 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_05379 5182 3072 3045 5182 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_05380 5182 3049 3048 5182 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_05381 3047 5198 5182 5182 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_05382 5182 5198 3049 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05383 5182 3052 3051 5182 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_05384 3050 5197 5182 5182 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_05385 5182 5197 3052 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05386 5182 3055 3054 5182 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_05387 3053 5196 5182 5182 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_05388 5182 5196 3055 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05389 5182 3058 3057 5182 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_05390 3056 5195 5182 5182 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_05391 5182 5195 3058 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05392 5182 3061 3060 5182 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_05393 3059 5194 5182 5182 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_05394 5182 5194 3061 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_05395 5182 5200 3062 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05396 5182 5199 3063 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05397 5182 5200 391 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_05398 391 3063 3069 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_05399 3070 5200 392 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_05400 392 5199 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_05401 5182 3062 393 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_05402 393 3063 3065 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_05403 3066 3062 394 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_05404 394 5199 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_05405 5182 3065 3064 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05406 3067 3066 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05407 5182 3069 3068 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05408 3071 3070 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05409 3072 3073 5182 5182 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_05410 5182 5201 3073 5182 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_05411 3074 3075 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05412 5182 3075 3074 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05413 3075 3078 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05414 5176 3076 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05415 5182 3076 5176 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05416 3076 3079 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05417 3077 3078 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05418 5182 3078 3077 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05419 395 3085 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05420 3078 5181 395 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05421 5179 3079 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05422 5182 3079 5179 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05423 396 3085 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05424 3079 5181 396 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05425 3080 3084 397 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05426 397 3086 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05427 5182 3080 3081 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05428 3081 3080 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05429 3082 3084 398 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05430 398 3086 5182 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05431 5182 3082 3083 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05432 3083 3082 5182 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_05433 5182 3085 3084 5182 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_05434 3085 3086 5182 5182 tn L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_05435 5182 3086 3085 5182 tn L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_05436 399 5193 3086 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05437 5182 5184 399 5182 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_05438 403 2528 401 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05439 403 2528 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_05440 401 2528 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_05441 402 2528 400 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05442 5183 2528 402 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_05443 5183 2528 400 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_05444 5182 3088 3087 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05445 3088 3087 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05446 403 2536 3087 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05447 401 2536 3088 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05448 5182 3090 3089 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05449 3090 3089 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05450 402 2536 3089 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05451 400 2536 3090 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05452 5182 3092 3091 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05453 3092 3091 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05454 403 2534 3091 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05455 401 2534 3092 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05456 5182 3094 3093 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05457 3094 3093 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05458 402 2534 3093 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05459 400 2534 3094 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05460 5182 3096 3095 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05461 3096 3095 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05462 403 2535 3095 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05463 401 2535 3096 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05464 5182 3098 3097 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05465 3098 3097 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05466 402 2535 3097 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05467 400 2535 3098 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05468 5182 3100 3099 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05469 3100 3099 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05470 403 2533 3099 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05471 401 2533 3100 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05472 5182 3102 3101 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05473 3102 3101 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05474 402 2533 3101 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05475 400 2533 3102 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05476 5182 3104 3103 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05477 3104 3103 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05478 403 2552 3103 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05479 401 2552 3104 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05480 5182 3106 3105 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05481 3106 3105 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05482 402 2552 3105 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05483 400 2552 3106 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05484 5182 3108 3107 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05485 3108 3107 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05486 403 2550 3107 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05487 401 2550 3108 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05488 5182 3110 3109 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05489 3110 3109 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05490 402 2550 3109 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05491 400 2550 3110 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05492 5182 3112 3111 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05493 3112 3111 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05494 403 2551 3111 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05495 401 2551 3112 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05496 5182 3114 3113 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05497 3114 3113 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05498 402 2551 3113 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05499 400 2551 3114 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05500 5182 3116 3115 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05501 3116 3115 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05502 403 2549 3115 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05503 401 2549 3116 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05504 5182 3118 3117 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05505 3118 3117 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05506 402 2549 3117 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05507 400 2549 3118 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05508 5182 3120 3119 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05509 3120 3119 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05510 403 2568 3119 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05511 401 2568 3120 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05512 5182 3122 3121 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05513 3122 3121 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05514 402 2568 3121 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05515 400 2568 3122 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05516 5182 3124 3123 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05517 3124 3123 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05518 403 2566 3123 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05519 401 2566 3124 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05520 5182 3126 3125 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05521 3126 3125 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05522 402 2566 3125 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05523 400 2566 3126 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05524 5182 3128 3127 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05525 3128 3127 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05526 403 2567 3127 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05527 401 2567 3128 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05528 5182 3130 3129 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05529 3130 3129 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05530 402 2567 3129 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05531 400 2567 3130 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05532 5182 3132 3131 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05533 3132 3131 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05534 403 2565 3131 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05535 401 2565 3132 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05536 5182 3134 3133 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05537 3134 3133 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05538 402 2565 3133 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05539 400 2565 3134 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05540 5182 3136 3135 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05541 3136 3135 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05542 403 2584 3135 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05543 401 2584 3136 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05544 5182 3138 3137 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05545 3138 3137 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05546 402 2584 3137 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05547 400 2584 3138 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05548 5182 3140 3139 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05549 3140 3139 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05550 403 2582 3139 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05551 401 2582 3140 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05552 5182 3142 3141 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05553 3142 3141 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05554 402 2582 3141 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05555 400 2582 3142 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05556 5182 3144 3143 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05557 3144 3143 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05558 403 2583 3143 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05559 401 2583 3144 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05560 5182 3146 3145 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05561 3146 3145 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05562 402 2583 3145 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05563 400 2583 3146 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05564 5182 3148 3147 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05565 3148 3147 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05566 403 2581 3147 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05567 401 2581 3148 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05568 5182 3150 3149 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05569 3150 3149 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05570 402 2581 3149 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05571 400 2581 3150 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05572 5182 3152 3151 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05573 3152 3151 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05574 403 2600 3151 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05575 401 2600 3152 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05576 5182 3154 3153 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05577 3154 3153 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05578 402 2600 3153 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05579 400 2600 3154 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05580 5182 3156 3155 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05581 3156 3155 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05582 403 2598 3155 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05583 401 2598 3156 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05584 5182 3158 3157 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05585 3158 3157 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05586 402 2598 3157 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05587 400 2598 3158 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05588 5182 3160 3159 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05589 3160 3159 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05590 403 2599 3159 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05591 401 2599 3160 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05592 5182 3162 3161 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05593 3162 3161 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05594 402 2599 3161 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05595 400 2599 3162 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05596 5182 3164 3163 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05597 3164 3163 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05598 403 2597 3163 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05599 401 2597 3164 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05600 5182 3166 3165 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05601 3166 3165 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05602 402 2597 3165 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05603 400 2597 3166 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05604 5182 3168 3167 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05605 3168 3167 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05606 403 2616 3167 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05607 401 2616 3168 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05608 5182 3170 3169 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05609 3170 3169 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05610 402 2616 3169 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05611 400 2616 3170 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05612 5182 3172 3171 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05613 3172 3171 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05614 403 2614 3171 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05615 401 2614 3172 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05616 5182 3174 3173 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05617 3174 3173 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05618 402 2614 3173 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05619 400 2614 3174 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05620 5182 3176 3175 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05621 3176 3175 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05622 403 2615 3175 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05623 401 2615 3176 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05624 5182 3178 3177 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05625 3178 3177 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05626 402 2615 3177 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05627 400 2615 3178 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05628 5182 3180 3179 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05629 3180 3179 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05630 403 2613 3179 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05631 401 2613 3180 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05632 5182 3182 3181 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05633 3182 3181 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05634 402 2613 3181 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05635 400 2613 3182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05636 5182 3184 3183 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05637 3184 3183 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05638 403 2632 3183 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05639 401 2632 3184 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05640 5182 3186 3185 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05641 3186 3185 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05642 402 2632 3185 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05643 400 2632 3186 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05644 5182 3188 3187 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05645 3188 3187 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05646 403 2630 3187 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05647 401 2630 3188 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05648 5182 3190 3189 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05649 3190 3189 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05650 402 2630 3189 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05651 400 2630 3190 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05652 5182 3192 3191 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05653 3192 3191 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05654 403 2631 3191 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05655 401 2631 3192 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05656 5182 3194 3193 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05657 3194 3193 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05658 402 2631 3193 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05659 400 2631 3194 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05660 5182 3196 3195 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05661 3196 3195 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05662 403 2629 3195 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05663 401 2629 3196 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05664 5182 3198 3197 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05665 3198 3197 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05666 402 2629 3197 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05667 400 2629 3198 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05668 5182 3200 3199 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05669 3200 3199 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05670 403 2648 3199 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05671 401 2648 3200 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05672 5182 3202 3201 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05673 3202 3201 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05674 402 2648 3201 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05675 400 2648 3202 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05676 5182 3204 3203 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05677 3204 3203 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05678 403 2646 3203 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05679 401 2646 3204 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05680 5182 3206 3205 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05681 3206 3205 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05682 402 2646 3205 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05683 400 2646 3206 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05684 5182 3208 3207 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05685 3208 3207 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05686 403 2647 3207 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05687 401 2647 3208 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05688 5182 3210 3209 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05689 3210 3209 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05690 402 2647 3209 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05691 400 2647 3210 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05692 5182 3212 3211 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05693 3212 3211 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05694 403 2645 3211 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05695 401 2645 3212 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05696 5182 3214 3213 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05697 3214 3213 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05698 402 2645 3213 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05699 400 2645 3214 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05700 5182 3216 3215 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05701 3216 3215 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05702 403 2664 3215 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05703 401 2664 3216 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05704 5182 3218 3217 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05705 3218 3217 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05706 402 2664 3217 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05707 400 2664 3218 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05708 5182 3220 3219 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05709 3220 3219 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05710 403 2662 3219 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05711 401 2662 3220 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05712 5182 3222 3221 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05713 3222 3221 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05714 402 2662 3221 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05715 400 2662 3222 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05716 5182 3224 3223 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05717 3224 3223 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05718 403 2663 3223 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05719 401 2663 3224 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05720 5182 3226 3225 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05721 3226 3225 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05722 402 2663 3225 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05723 400 2663 3226 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05724 5182 3228 3227 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05725 3228 3227 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05726 403 2661 3227 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05727 401 2661 3228 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05728 5182 3230 3229 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05729 3230 3229 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05730 402 2661 3229 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05731 400 2661 3230 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05732 5182 3232 3231 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05733 3232 3231 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05734 403 2680 3231 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05735 401 2680 3232 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05736 5182 3234 3233 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05737 3234 3233 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05738 402 2680 3233 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05739 400 2680 3234 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05740 5182 3236 3235 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05741 3236 3235 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05742 403 2678 3235 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05743 401 2678 3236 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05744 5182 3238 3237 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05745 3238 3237 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05746 402 2678 3237 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05747 400 2678 3238 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05748 5182 3240 3239 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05749 3240 3239 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05750 403 2679 3239 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05751 401 2679 3240 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05752 5182 3242 3241 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05753 3242 3241 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05754 402 2679 3241 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05755 400 2679 3242 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05756 5182 3244 3243 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05757 3244 3243 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05758 403 2677 3243 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05759 401 2677 3244 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05760 5182 3246 3245 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05761 3246 3245 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05762 402 2677 3245 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05763 400 2677 3246 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05764 5182 3248 3247 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05765 3248 3247 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05766 403 2696 3247 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05767 401 2696 3248 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05768 5182 3250 3249 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05769 3250 3249 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05770 402 2696 3249 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05771 400 2696 3250 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05772 5182 3252 3251 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05773 3252 3251 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05774 403 2694 3251 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05775 401 2694 3252 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05776 5182 3254 3253 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05777 3254 3253 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05778 402 2694 3253 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05779 400 2694 3254 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05780 5182 3256 3255 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05781 3256 3255 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05782 403 2695 3255 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05783 401 2695 3256 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05784 5182 3258 3257 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05785 3258 3257 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05786 402 2695 3257 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05787 400 2695 3258 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05788 5182 3260 3259 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05789 3260 3259 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05790 403 2693 3259 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05791 401 2693 3260 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05792 5182 3262 3261 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05793 3262 3261 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05794 402 2693 3261 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05795 400 2693 3262 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05796 5182 3264 3263 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05797 3264 3263 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05798 403 2712 3263 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05799 401 2712 3264 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05800 5182 3266 3265 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05801 3266 3265 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05802 402 2712 3265 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05803 400 2712 3266 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05804 5182 3268 3267 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05805 3268 3267 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05806 403 2710 3267 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05807 401 2710 3268 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05808 5182 3270 3269 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05809 3270 3269 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05810 402 2710 3269 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05811 400 2710 3270 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05812 5182 3272 3271 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05813 3272 3271 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05814 403 2711 3271 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05815 401 2711 3272 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05816 5182 3274 3273 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05817 3274 3273 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05818 402 2711 3273 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05819 400 2711 3274 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05820 5182 3276 3275 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05821 3276 3275 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05822 403 2709 3275 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05823 401 2709 3276 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05824 5182 3278 3277 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05825 3278 3277 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05826 402 2709 3277 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05827 400 2709 3278 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05828 5182 3280 3279 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05829 3280 3279 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05830 403 2728 3279 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05831 401 2728 3280 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05832 5182 3282 3281 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05833 3282 3281 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05834 402 2728 3281 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05835 400 2728 3282 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05836 5182 3284 3283 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05837 3284 3283 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05838 403 2726 3283 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05839 401 2726 3284 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05840 5182 3286 3285 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05841 3286 3285 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05842 402 2726 3285 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05843 400 2726 3286 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05844 5182 3288 3287 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05845 3288 3287 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05846 403 2727 3287 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05847 401 2727 3288 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05848 5182 3290 3289 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05849 3290 3289 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05850 402 2727 3289 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05851 400 2727 3290 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05852 5182 3292 3291 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05853 3292 3291 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05854 403 2725 3291 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05855 401 2725 3292 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05856 5182 3294 3293 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05857 3294 3293 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05858 402 2725 3293 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05859 400 2725 3294 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05860 5182 3296 3295 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05861 3296 3295 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05862 403 2744 3295 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05863 401 2744 3296 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05864 5182 3298 3297 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05865 3298 3297 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05866 402 2744 3297 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05867 400 2744 3298 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05868 5182 3300 3299 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05869 3300 3299 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05870 403 2742 3299 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05871 401 2742 3300 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05872 5182 3302 3301 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05873 3302 3301 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05874 402 2742 3301 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05875 400 2742 3302 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05876 5182 3304 3303 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05877 3304 3303 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05878 403 2743 3303 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05879 401 2743 3304 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05880 5182 3306 3305 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05881 3306 3305 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05882 402 2743 3305 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05883 400 2743 3306 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05884 5182 3308 3307 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05885 3308 3307 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05886 403 2741 3307 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05887 401 2741 3308 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05888 5182 3310 3309 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05889 3310 3309 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05890 402 2741 3309 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05891 400 2741 3310 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05892 5182 3312 3311 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05893 3312 3311 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05894 403 2760 3311 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05895 401 2760 3312 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05896 5182 3314 3313 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05897 3314 3313 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05898 402 2760 3313 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05899 400 2760 3314 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05900 5182 3316 3315 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05901 3316 3315 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05902 403 2758 3315 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05903 401 2758 3316 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05904 5182 3318 3317 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05905 3318 3317 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05906 402 2758 3317 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05907 400 2758 3318 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05908 5182 3320 3319 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05909 3320 3319 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05910 403 2759 3319 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05911 401 2759 3320 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05912 5182 3322 3321 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05913 3322 3321 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05914 402 2759 3321 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05915 400 2759 3322 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05916 5182 3324 3323 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05917 3324 3323 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05918 403 2757 3323 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05919 401 2757 3324 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05920 5182 3326 3325 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05921 3326 3325 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05922 402 2757 3325 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05923 400 2757 3326 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05924 5182 3328 3327 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05925 3328 3327 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05926 403 2776 3327 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05927 401 2776 3328 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05928 5182 3330 3329 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05929 3330 3329 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05930 402 2776 3329 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05931 400 2776 3330 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05932 5182 3332 3331 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05933 3332 3331 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05934 403 2774 3331 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05935 401 2774 3332 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05936 5182 3334 3333 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05937 3334 3333 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05938 402 2774 3333 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05939 400 2774 3334 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05940 5182 3336 3335 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05941 3336 3335 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05942 403 2775 3335 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05943 401 2775 3336 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05944 5182 3338 3337 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05945 3338 3337 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05946 402 2775 3337 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05947 400 2775 3338 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05948 5182 3340 3339 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05949 3340 3339 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05950 403 2773 3339 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05951 401 2773 3340 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05952 5182 3342 3341 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05953 3342 3341 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05954 402 2773 3341 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05955 400 2773 3342 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05956 5182 3344 3343 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05957 3344 3343 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05958 403 2792 3343 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05959 401 2792 3344 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05960 5182 3346 3345 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05961 3346 3345 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05962 402 2792 3345 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05963 400 2792 3346 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05964 5182 3348 3347 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05965 3348 3347 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05966 403 2790 3347 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05967 401 2790 3348 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05968 5182 3350 3349 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05969 3350 3349 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05970 402 2790 3349 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05971 400 2790 3350 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05972 5182 3352 3351 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05973 3352 3351 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05974 403 2791 3351 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05975 401 2791 3352 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05976 5182 3354 3353 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05977 3354 3353 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05978 402 2791 3353 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05979 400 2791 3354 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05980 5182 3356 3355 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05981 3356 3355 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05982 403 2789 3355 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05983 401 2789 3356 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05984 5182 3358 3357 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05985 3358 3357 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05986 402 2789 3357 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05987 400 2789 3358 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05988 5182 3360 3359 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05989 3360 3359 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05990 403 2808 3359 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05991 401 2808 3360 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05992 5182 3362 3361 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05993 3362 3361 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05994 402 2808 3361 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05995 400 2808 3362 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05996 5182 3364 3363 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05997 3364 3363 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05998 403 2806 3363 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_05999 401 2806 3364 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06000 5182 3366 3365 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06001 3366 3365 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06002 402 2806 3365 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06003 400 2806 3366 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06004 5182 3368 3367 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06005 3368 3367 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06006 403 2807 3367 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06007 401 2807 3368 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06008 5182 3370 3369 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06009 3370 3369 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06010 402 2807 3369 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06011 400 2807 3370 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06012 5182 3372 3371 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06013 3372 3371 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06014 403 2805 3371 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06015 401 2805 3372 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06016 5182 3374 3373 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06017 3374 3373 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06018 402 2805 3373 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06019 400 2805 3374 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06020 5182 3376 3375 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06021 3376 3375 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06022 403 2824 3375 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06023 401 2824 3376 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06024 5182 3378 3377 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06025 3378 3377 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06026 402 2824 3377 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06027 400 2824 3378 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06028 5182 3380 3379 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06029 3380 3379 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06030 403 2822 3379 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06031 401 2822 3380 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06032 5182 3382 3381 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06033 3382 3381 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06034 402 2822 3381 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06035 400 2822 3382 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06036 5182 3384 3383 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06037 3384 3383 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06038 403 2823 3383 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06039 401 2823 3384 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06040 5182 3386 3385 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06041 3386 3385 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06042 402 2823 3385 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06043 400 2823 3386 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06044 5182 3388 3387 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06045 3388 3387 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06046 403 2821 3387 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06047 401 2821 3388 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06048 5182 3390 3389 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06049 3390 3389 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06050 402 2821 3389 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06051 400 2821 3390 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06052 5182 3392 3391 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06053 3392 3391 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06054 403 2840 3391 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06055 401 2840 3392 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06056 5182 3394 3393 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06057 3394 3393 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06058 402 2840 3393 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06059 400 2840 3394 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06060 5182 3396 3395 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06061 3396 3395 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06062 403 2838 3395 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06063 401 2838 3396 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06064 5182 3398 3397 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06065 3398 3397 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06066 402 2838 3397 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06067 400 2838 3398 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06068 5182 3400 3399 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06069 3400 3399 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06070 403 2839 3399 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06071 401 2839 3400 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06072 5182 3402 3401 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06073 3402 3401 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06074 402 2839 3401 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06075 400 2839 3402 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06076 5182 3404 3403 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06077 3404 3403 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06078 403 2837 3403 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06079 401 2837 3404 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06080 5182 3406 3405 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06081 3406 3405 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06082 402 2837 3405 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06083 400 2837 3406 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06084 5182 3408 3407 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06085 3408 3407 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06086 403 2856 3407 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06087 401 2856 3408 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06088 5182 3410 3409 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06089 3410 3409 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06090 402 2856 3409 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06091 400 2856 3410 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06092 5182 3412 3411 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06093 3412 3411 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06094 403 2854 3411 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06095 401 2854 3412 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06096 5182 3414 3413 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06097 3414 3413 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06098 402 2854 3413 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06099 400 2854 3414 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06100 5182 3416 3415 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06101 3416 3415 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06102 403 2855 3415 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06103 401 2855 3416 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06104 5182 3418 3417 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06105 3418 3417 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06106 402 2855 3417 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06107 400 2855 3418 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06108 5182 3420 3419 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06109 3420 3419 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06110 403 2853 3419 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06111 401 2853 3420 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06112 5182 3422 3421 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06113 3422 3421 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06114 402 2853 3421 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06115 400 2853 3422 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06116 5182 3424 3423 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06117 3424 3423 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06118 403 2872 3423 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06119 401 2872 3424 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06120 5182 3426 3425 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06121 3426 3425 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06122 402 2872 3425 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06123 400 2872 3426 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06124 5182 3428 3427 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06125 3428 3427 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06126 403 2870 3427 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06127 401 2870 3428 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06128 5182 3430 3429 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06129 3430 3429 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06130 402 2870 3429 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06131 400 2870 3430 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06132 5182 3432 3431 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06133 3432 3431 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06134 403 2871 3431 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06135 401 2871 3432 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06136 5182 3434 3433 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06137 3434 3433 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06138 402 2871 3433 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06139 400 2871 3434 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06140 5182 3436 3435 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06141 3436 3435 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06142 403 2869 3435 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06143 401 2869 3436 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06144 5182 3438 3437 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06145 3438 3437 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06146 402 2869 3437 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06147 400 2869 3438 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06148 5182 3440 3439 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06149 3440 3439 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06150 403 2888 3439 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06151 401 2888 3440 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06152 5182 3442 3441 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06153 3442 3441 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06154 402 2888 3441 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06155 400 2888 3442 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06156 5182 3444 3443 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06157 3444 3443 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06158 403 2886 3443 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06159 401 2886 3444 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06160 5182 3446 3445 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06161 3446 3445 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06162 402 2886 3445 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06163 400 2886 3446 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06164 5182 3448 3447 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06165 3448 3447 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06166 403 2887 3447 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06167 401 2887 3448 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06168 5182 3450 3449 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06169 3450 3449 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06170 402 2887 3449 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06171 400 2887 3450 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06172 5182 3452 3451 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06173 3452 3451 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06174 403 2885 3451 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06175 401 2885 3452 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06176 5182 3454 3453 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06177 3454 3453 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06178 402 2885 3453 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06179 400 2885 3454 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06180 5182 3456 3455 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06181 3456 3455 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06182 403 2904 3455 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06183 401 2904 3456 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06184 5182 3458 3457 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06185 3458 3457 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06186 402 2904 3457 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06187 400 2904 3458 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06188 5182 3460 3459 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06189 3460 3459 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06190 403 2902 3459 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06191 401 2902 3460 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06192 5182 3462 3461 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06193 3462 3461 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06194 402 2902 3461 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06195 400 2902 3462 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06196 5182 3464 3463 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06197 3464 3463 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06198 403 2903 3463 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06199 401 2903 3464 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06200 5182 3466 3465 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06201 3466 3465 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06202 402 2903 3465 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06203 400 2903 3466 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06204 5182 3468 3467 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06205 3468 3467 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06206 403 2901 3467 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06207 401 2901 3468 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06208 5182 3470 3469 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06209 3470 3469 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06210 402 2901 3469 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06211 400 2901 3470 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06212 5182 3472 3471 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06213 3472 3471 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06214 403 2920 3471 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06215 401 2920 3472 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06216 5182 3474 3473 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06217 3474 3473 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06218 402 2920 3473 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06219 400 2920 3474 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06220 5182 3476 3475 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06221 3476 3475 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06222 403 2918 3475 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06223 401 2918 3476 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06224 5182 3478 3477 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06225 3478 3477 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06226 402 2918 3477 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06227 400 2918 3478 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06228 5182 3480 3479 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06229 3480 3479 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06230 403 2919 3479 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06231 401 2919 3480 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06232 5182 3482 3481 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06233 3482 3481 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06234 402 2919 3481 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06235 400 2919 3482 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06236 5182 3484 3483 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06237 3484 3483 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06238 403 2917 3483 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06239 401 2917 3484 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06240 5182 3486 3485 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06241 3486 3485 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06242 402 2917 3485 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06243 400 2917 3486 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06244 5182 3488 3487 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06245 3488 3487 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06246 403 2936 3487 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06247 401 2936 3488 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06248 5182 3490 3489 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06249 3490 3489 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06250 402 2936 3489 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06251 400 2936 3490 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06252 5182 3492 3491 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06253 3492 3491 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06254 403 2934 3491 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06255 401 2934 3492 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06256 5182 3494 3493 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06257 3494 3493 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06258 402 2934 3493 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06259 400 2934 3494 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06260 5182 3496 3495 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06261 3496 3495 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06262 403 2935 3495 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06263 401 2935 3496 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06264 5182 3498 3497 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06265 3498 3497 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06266 402 2935 3497 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06267 400 2935 3498 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06268 5182 3500 3499 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06269 3500 3499 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06270 403 2933 3499 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06271 401 2933 3500 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06272 5182 3502 3501 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06273 3502 3501 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06274 402 2933 3501 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06275 400 2933 3502 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06276 5182 3504 3503 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06277 3504 3503 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06278 403 2952 3503 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06279 401 2952 3504 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06280 5182 3506 3505 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06281 3506 3505 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06282 402 2952 3505 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06283 400 2952 3506 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06284 5182 3508 3507 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06285 3508 3507 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06286 403 2950 3507 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06287 401 2950 3508 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06288 5182 3510 3509 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06289 3510 3509 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06290 402 2950 3509 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06291 400 2950 3510 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06292 5182 3512 3511 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06293 3512 3511 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06294 403 2951 3511 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06295 401 2951 3512 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06296 5182 3514 3513 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06297 3514 3513 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06298 402 2951 3513 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06299 400 2951 3514 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06300 5182 3516 3515 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06301 3516 3515 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06302 403 2949 3515 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06303 401 2949 3516 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06304 5182 3518 3517 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06305 3518 3517 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06306 402 2949 3517 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06307 400 2949 3518 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06308 5182 3520 3519 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06309 3520 3519 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06310 403 2968 3519 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06311 401 2968 3520 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06312 5182 3522 3521 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06313 3522 3521 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06314 402 2968 3521 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06315 400 2968 3522 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06316 5182 3524 3523 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06317 3524 3523 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06318 403 2966 3523 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06319 401 2966 3524 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06320 5182 3526 3525 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06321 3526 3525 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06322 402 2966 3525 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06323 400 2966 3526 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06324 5182 3528 3527 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06325 3528 3527 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06326 403 2967 3527 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06327 401 2967 3528 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06328 5182 3530 3529 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06329 3530 3529 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06330 402 2967 3529 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06331 400 2967 3530 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06332 5182 3532 3531 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06333 3532 3531 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06334 403 2965 3531 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06335 401 2965 3532 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06336 5182 3534 3533 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06337 3534 3533 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06338 402 2965 3533 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06339 400 2965 3534 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06340 5182 3536 3535 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06341 3536 3535 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06342 403 2984 3535 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06343 401 2984 3536 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06344 5182 3538 3537 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06345 3538 3537 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06346 402 2984 3537 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06347 400 2984 3538 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06348 5182 3540 3539 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06349 3540 3539 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06350 403 2982 3539 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06351 401 2982 3540 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06352 5182 3542 3541 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06353 3542 3541 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06354 402 2982 3541 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06355 400 2982 3542 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06356 5182 3544 3543 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06357 3544 3543 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06358 403 2983 3543 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06359 401 2983 3544 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06360 5182 3546 3545 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06361 3546 3545 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06362 402 2983 3545 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06363 400 2983 3546 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06364 5182 3548 3547 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06365 3548 3547 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06366 403 2981 3547 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06367 401 2981 3548 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06368 5182 3550 3549 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06369 3550 3549 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06370 402 2981 3549 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06371 400 2981 3550 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06372 5182 3552 3551 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06373 3552 3551 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06374 403 3000 3551 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06375 401 3000 3552 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06376 5182 3554 3553 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06377 3554 3553 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06378 402 3000 3553 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06379 400 3000 3554 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06380 5182 3556 3555 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06381 3556 3555 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06382 403 2998 3555 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06383 401 2998 3556 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06384 5182 3558 3557 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06385 3558 3557 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06386 402 2998 3557 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06387 400 2998 3558 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06388 5182 3560 3559 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06389 3560 3559 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06390 403 2999 3559 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06391 401 2999 3560 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06392 5182 3562 3561 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06393 3562 3561 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06394 402 2999 3561 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06395 400 2999 3562 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06396 5182 3564 3563 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06397 3564 3563 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06398 403 2997 3563 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06399 401 2997 3564 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06400 5182 3566 3565 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06401 3566 3565 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06402 402 2997 3565 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06403 400 2997 3566 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06404 5182 3568 3567 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06405 3568 3567 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06406 403 3016 3567 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06407 401 3016 3568 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06408 5182 3570 3569 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06409 3570 3569 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06410 402 3016 3569 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06411 400 3016 3570 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06412 5182 3572 3571 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06413 3572 3571 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06414 403 3014 3571 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06415 401 3014 3572 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06416 5182 3574 3573 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06417 3574 3573 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06418 402 3014 3573 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06419 400 3014 3574 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06420 5182 3576 3575 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06421 3576 3575 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06422 403 3015 3575 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06423 401 3015 3576 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06424 5182 3578 3577 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06425 3578 3577 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06426 402 3015 3577 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06427 400 3015 3578 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06428 5182 3580 3579 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06429 3580 3579 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06430 403 3013 3579 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06431 401 3013 3580 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06432 5182 3582 3581 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06433 3582 3581 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06434 402 3013 3581 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06435 400 3013 3582 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06436 5182 3584 3583 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06437 3584 3583 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06438 403 3032 3583 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06439 401 3032 3584 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06440 5182 3586 3585 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06441 3586 3585 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06442 402 3032 3585 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06443 400 3032 3586 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06444 5182 3588 3587 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06445 3588 3587 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06446 403 3030 3587 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06447 401 3030 3588 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06448 5182 3590 3589 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06449 3590 3589 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06450 402 3030 3589 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06451 400 3030 3590 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06452 5182 3592 3591 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06453 3592 3591 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06454 403 3031 3591 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06455 401 3031 3592 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06456 5182 3594 3593 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06457 3594 3593 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06458 402 3031 3593 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06459 400 3031 3594 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06460 5182 3596 3595 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06461 3596 3595 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06462 403 3029 3595 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06463 401 3029 3596 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06464 5182 3598 3597 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06465 3598 3597 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06466 402 3029 3597 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06467 400 3029 3598 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06468 400 3045 407 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_06469 407 3046 401 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_06470 402 3045 408 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_06471 408 3046 403 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_06472 3602 3081 3600 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_06473 3607 3602 404 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_06474 404 5176 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_06475 404 3600 3599 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_06476 5182 5176 405 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_06477 3601 408 405 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_06478 405 407 3600 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_06479 3602 408 406 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_06480 406 5176 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_06481 406 407 3603 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_06482 5183 3081 408 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_06483 408 3081 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_06484 5183 3081 407 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_06485 407 3081 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_06486 3604 5179 408 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_06487 407 5179 3605 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_06488 408 3081 407 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_06489 5182 5188 3604 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_06490 3605 3606 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_06491 3604 5188 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_06492 5182 3606 3605 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_06493 5182 5188 3606 5182 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_06494 5188 3608 5182 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_06495 5182 3608 5188 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_06496 5182 5179 3608 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_06497 3608 3607 5182 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_06498 3608 5176 3609 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_06499 412 2528 410 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06500 412 2528 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_06501 410 2528 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_06502 411 2528 409 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06503 5183 2528 411 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_06504 5183 2528 409 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_06505 5182 3611 3610 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06506 3611 3610 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06507 412 2536 3610 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06508 410 2536 3611 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06509 5182 3613 3612 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06510 3613 3612 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06511 411 2536 3612 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06512 409 2536 3613 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06513 5182 3615 3614 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06514 3615 3614 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06515 412 2534 3614 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06516 410 2534 3615 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06517 5182 3617 3616 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06518 3617 3616 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06519 411 2534 3616 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06520 409 2534 3617 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06521 5182 3619 3618 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06522 3619 3618 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06523 412 2535 3618 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06524 410 2535 3619 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06525 5182 3621 3620 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06526 3621 3620 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06527 411 2535 3620 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06528 409 2535 3621 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06529 5182 3623 3622 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06530 3623 3622 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06531 412 2533 3622 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06532 410 2533 3623 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06533 5182 3625 3624 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06534 3625 3624 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06535 411 2533 3624 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06536 409 2533 3625 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06537 5182 3627 3626 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06538 3627 3626 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06539 412 2552 3626 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06540 410 2552 3627 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06541 5182 3629 3628 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06542 3629 3628 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06543 411 2552 3628 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06544 409 2552 3629 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06545 5182 3631 3630 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06546 3631 3630 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06547 412 2550 3630 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06548 410 2550 3631 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06549 5182 3633 3632 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06550 3633 3632 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06551 411 2550 3632 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06552 409 2550 3633 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06553 5182 3635 3634 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06554 3635 3634 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06555 412 2551 3634 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06556 410 2551 3635 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06557 5182 3637 3636 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06558 3637 3636 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06559 411 2551 3636 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06560 409 2551 3637 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06561 5182 3639 3638 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06562 3639 3638 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06563 412 2549 3638 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06564 410 2549 3639 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06565 5182 3641 3640 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06566 3641 3640 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06567 411 2549 3640 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06568 409 2549 3641 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06569 5182 3643 3642 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06570 3643 3642 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06571 412 2568 3642 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06572 410 2568 3643 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06573 5182 3645 3644 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06574 3645 3644 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06575 411 2568 3644 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06576 409 2568 3645 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06577 5182 3647 3646 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06578 3647 3646 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06579 412 2566 3646 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06580 410 2566 3647 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06581 5182 3649 3648 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06582 3649 3648 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06583 411 2566 3648 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06584 409 2566 3649 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06585 5182 3651 3650 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06586 3651 3650 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06587 412 2567 3650 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06588 410 2567 3651 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06589 5182 3653 3652 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06590 3653 3652 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06591 411 2567 3652 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06592 409 2567 3653 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06593 5182 3655 3654 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06594 3655 3654 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06595 412 2565 3654 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06596 410 2565 3655 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06597 5182 3657 3656 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06598 3657 3656 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06599 411 2565 3656 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06600 409 2565 3657 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06601 5182 3659 3658 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06602 3659 3658 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06603 412 2584 3658 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06604 410 2584 3659 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06605 5182 3661 3660 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06606 3661 3660 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06607 411 2584 3660 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06608 409 2584 3661 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06609 5182 3663 3662 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06610 3663 3662 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06611 412 2582 3662 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06612 410 2582 3663 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06613 5182 3665 3664 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06614 3665 3664 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06615 411 2582 3664 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06616 409 2582 3665 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06617 5182 3667 3666 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06618 3667 3666 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06619 412 2583 3666 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06620 410 2583 3667 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06621 5182 3669 3668 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06622 3669 3668 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06623 411 2583 3668 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06624 409 2583 3669 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06625 5182 3671 3670 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06626 3671 3670 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06627 412 2581 3670 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06628 410 2581 3671 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06629 5182 3673 3672 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06630 3673 3672 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06631 411 2581 3672 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06632 409 2581 3673 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06633 5182 3675 3674 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06634 3675 3674 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06635 412 2600 3674 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06636 410 2600 3675 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06637 5182 3677 3676 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06638 3677 3676 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06639 411 2600 3676 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06640 409 2600 3677 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06641 5182 3679 3678 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06642 3679 3678 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06643 412 2598 3678 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06644 410 2598 3679 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06645 5182 3681 3680 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06646 3681 3680 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06647 411 2598 3680 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06648 409 2598 3681 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06649 5182 3683 3682 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06650 3683 3682 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06651 412 2599 3682 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06652 410 2599 3683 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06653 5182 3685 3684 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06654 3685 3684 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06655 411 2599 3684 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06656 409 2599 3685 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06657 5182 3687 3686 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06658 3687 3686 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06659 412 2597 3686 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06660 410 2597 3687 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06661 5182 3689 3688 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06662 3689 3688 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06663 411 2597 3688 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06664 409 2597 3689 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06665 5182 3691 3690 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06666 3691 3690 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06667 412 2616 3690 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06668 410 2616 3691 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06669 5182 3693 3692 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06670 3693 3692 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06671 411 2616 3692 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06672 409 2616 3693 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06673 5182 3695 3694 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06674 3695 3694 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06675 412 2614 3694 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06676 410 2614 3695 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06677 5182 3697 3696 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06678 3697 3696 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06679 411 2614 3696 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06680 409 2614 3697 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06681 5182 3699 3698 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06682 3699 3698 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06683 412 2615 3698 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06684 410 2615 3699 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06685 5182 3701 3700 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06686 3701 3700 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06687 411 2615 3700 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06688 409 2615 3701 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06689 5182 3703 3702 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06690 3703 3702 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06691 412 2613 3702 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06692 410 2613 3703 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06693 5182 3705 3704 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06694 3705 3704 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06695 411 2613 3704 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06696 409 2613 3705 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06697 5182 3707 3706 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06698 3707 3706 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06699 412 2632 3706 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06700 410 2632 3707 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06701 5182 3709 3708 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06702 3709 3708 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06703 411 2632 3708 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06704 409 2632 3709 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06705 5182 3711 3710 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06706 3711 3710 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06707 412 2630 3710 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06708 410 2630 3711 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06709 5182 3713 3712 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06710 3713 3712 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06711 411 2630 3712 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06712 409 2630 3713 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06713 5182 3715 3714 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06714 3715 3714 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06715 412 2631 3714 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06716 410 2631 3715 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06717 5182 3717 3716 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06718 3717 3716 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06719 411 2631 3716 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06720 409 2631 3717 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06721 5182 3719 3718 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06722 3719 3718 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06723 412 2629 3718 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06724 410 2629 3719 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06725 5182 3721 3720 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06726 3721 3720 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06727 411 2629 3720 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06728 409 2629 3721 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06729 5182 3723 3722 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06730 3723 3722 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06731 412 2648 3722 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06732 410 2648 3723 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06733 5182 3725 3724 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06734 3725 3724 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06735 411 2648 3724 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06736 409 2648 3725 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06737 5182 3727 3726 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06738 3727 3726 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06739 412 2646 3726 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06740 410 2646 3727 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06741 5182 3729 3728 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06742 3729 3728 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06743 411 2646 3728 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06744 409 2646 3729 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06745 5182 3731 3730 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06746 3731 3730 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06747 412 2647 3730 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06748 410 2647 3731 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06749 5182 3733 3732 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06750 3733 3732 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06751 411 2647 3732 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06752 409 2647 3733 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06753 5182 3735 3734 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06754 3735 3734 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06755 412 2645 3734 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06756 410 2645 3735 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06757 5182 3737 3736 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06758 3737 3736 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06759 411 2645 3736 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06760 409 2645 3737 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06761 5182 3739 3738 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06762 3739 3738 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06763 412 2664 3738 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06764 410 2664 3739 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06765 5182 3741 3740 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06766 3741 3740 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06767 411 2664 3740 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06768 409 2664 3741 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06769 5182 3743 3742 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06770 3743 3742 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06771 412 2662 3742 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06772 410 2662 3743 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06773 5182 3745 3744 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06774 3745 3744 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06775 411 2662 3744 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06776 409 2662 3745 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06777 5182 3747 3746 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06778 3747 3746 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06779 412 2663 3746 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06780 410 2663 3747 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06781 5182 3749 3748 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06782 3749 3748 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06783 411 2663 3748 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06784 409 2663 3749 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06785 5182 3751 3750 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06786 3751 3750 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06787 412 2661 3750 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06788 410 2661 3751 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06789 5182 3753 3752 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06790 3753 3752 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06791 411 2661 3752 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06792 409 2661 3753 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06793 5182 3755 3754 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06794 3755 3754 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06795 412 2680 3754 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06796 410 2680 3755 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06797 5182 3757 3756 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06798 3757 3756 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06799 411 2680 3756 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06800 409 2680 3757 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06801 5182 3759 3758 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06802 3759 3758 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06803 412 2678 3758 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06804 410 2678 3759 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06805 5182 3761 3760 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06806 3761 3760 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06807 411 2678 3760 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06808 409 2678 3761 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06809 5182 3763 3762 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06810 3763 3762 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06811 412 2679 3762 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06812 410 2679 3763 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06813 5182 3765 3764 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06814 3765 3764 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06815 411 2679 3764 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06816 409 2679 3765 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06817 5182 3767 3766 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06818 3767 3766 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06819 412 2677 3766 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06820 410 2677 3767 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06821 5182 3769 3768 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06822 3769 3768 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06823 411 2677 3768 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06824 409 2677 3769 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06825 5182 3771 3770 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06826 3771 3770 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06827 412 2696 3770 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06828 410 2696 3771 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06829 5182 3773 3772 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06830 3773 3772 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06831 411 2696 3772 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06832 409 2696 3773 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06833 5182 3775 3774 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06834 3775 3774 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06835 412 2694 3774 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06836 410 2694 3775 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06837 5182 3777 3776 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06838 3777 3776 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06839 411 2694 3776 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06840 409 2694 3777 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06841 5182 3779 3778 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06842 3779 3778 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06843 412 2695 3778 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06844 410 2695 3779 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06845 5182 3781 3780 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06846 3781 3780 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06847 411 2695 3780 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06848 409 2695 3781 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06849 5182 3783 3782 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06850 3783 3782 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06851 412 2693 3782 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06852 410 2693 3783 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06853 5182 3785 3784 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06854 3785 3784 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06855 411 2693 3784 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06856 409 2693 3785 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06857 5182 3787 3786 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06858 3787 3786 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06859 412 2712 3786 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06860 410 2712 3787 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06861 5182 3789 3788 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06862 3789 3788 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06863 411 2712 3788 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06864 409 2712 3789 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06865 5182 3791 3790 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06866 3791 3790 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06867 412 2710 3790 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06868 410 2710 3791 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06869 5182 3793 3792 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06870 3793 3792 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06871 411 2710 3792 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06872 409 2710 3793 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06873 5182 3795 3794 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06874 3795 3794 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06875 412 2711 3794 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06876 410 2711 3795 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06877 5182 3797 3796 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06878 3797 3796 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06879 411 2711 3796 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06880 409 2711 3797 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06881 5182 3799 3798 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06882 3799 3798 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06883 412 2709 3798 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06884 410 2709 3799 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06885 5182 3801 3800 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06886 3801 3800 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06887 411 2709 3800 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06888 409 2709 3801 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06889 5182 3803 3802 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06890 3803 3802 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06891 412 2728 3802 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06892 410 2728 3803 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06893 5182 3805 3804 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06894 3805 3804 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06895 411 2728 3804 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06896 409 2728 3805 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06897 5182 3807 3806 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06898 3807 3806 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06899 412 2726 3806 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06900 410 2726 3807 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06901 5182 3809 3808 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06902 3809 3808 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06903 411 2726 3808 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06904 409 2726 3809 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06905 5182 3811 3810 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06906 3811 3810 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06907 412 2727 3810 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06908 410 2727 3811 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06909 5182 3813 3812 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06910 3813 3812 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06911 411 2727 3812 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06912 409 2727 3813 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06913 5182 3815 3814 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06914 3815 3814 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06915 412 2725 3814 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06916 410 2725 3815 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06917 5182 3817 3816 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06918 3817 3816 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06919 411 2725 3816 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06920 409 2725 3817 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06921 5182 3819 3818 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06922 3819 3818 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06923 412 2744 3818 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06924 410 2744 3819 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06925 5182 3821 3820 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06926 3821 3820 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06927 411 2744 3820 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06928 409 2744 3821 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06929 5182 3823 3822 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06930 3823 3822 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06931 412 2742 3822 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06932 410 2742 3823 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06933 5182 3825 3824 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06934 3825 3824 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06935 411 2742 3824 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06936 409 2742 3825 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06937 5182 3827 3826 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06938 3827 3826 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06939 412 2743 3826 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06940 410 2743 3827 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06941 5182 3829 3828 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06942 3829 3828 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06943 411 2743 3828 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06944 409 2743 3829 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06945 5182 3831 3830 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06946 3831 3830 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06947 412 2741 3830 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06948 410 2741 3831 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06949 5182 3833 3832 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06950 3833 3832 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06951 411 2741 3832 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06952 409 2741 3833 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06953 5182 3835 3834 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06954 3835 3834 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06955 412 2760 3834 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06956 410 2760 3835 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06957 5182 3837 3836 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06958 3837 3836 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06959 411 2760 3836 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06960 409 2760 3837 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06961 5182 3839 3838 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06962 3839 3838 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06963 412 2758 3838 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06964 410 2758 3839 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06965 5182 3841 3840 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06966 3841 3840 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06967 411 2758 3840 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06968 409 2758 3841 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06969 5182 3843 3842 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06970 3843 3842 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06971 412 2759 3842 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06972 410 2759 3843 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06973 5182 3845 3844 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06974 3845 3844 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06975 411 2759 3844 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06976 409 2759 3845 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06977 5182 3847 3846 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06978 3847 3846 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06979 412 2757 3846 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06980 410 2757 3847 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06981 5182 3849 3848 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06982 3849 3848 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06983 411 2757 3848 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06984 409 2757 3849 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06985 5182 3851 3850 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06986 3851 3850 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06987 412 2776 3850 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06988 410 2776 3851 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06989 5182 3853 3852 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06990 3853 3852 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06991 411 2776 3852 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06992 409 2776 3853 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06993 5182 3855 3854 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06994 3855 3854 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06995 412 2774 3854 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06996 410 2774 3855 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06997 5182 3857 3856 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06998 3857 3856 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_06999 411 2774 3856 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07000 409 2774 3857 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07001 5182 3859 3858 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07002 3859 3858 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07003 412 2775 3858 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07004 410 2775 3859 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07005 5182 3861 3860 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07006 3861 3860 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07007 411 2775 3860 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07008 409 2775 3861 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07009 5182 3863 3862 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07010 3863 3862 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07011 412 2773 3862 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07012 410 2773 3863 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07013 5182 3865 3864 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07014 3865 3864 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07015 411 2773 3864 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07016 409 2773 3865 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07017 5182 3867 3866 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07018 3867 3866 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07019 412 2792 3866 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07020 410 2792 3867 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07021 5182 3869 3868 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07022 3869 3868 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07023 411 2792 3868 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07024 409 2792 3869 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07025 5182 3871 3870 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07026 3871 3870 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07027 412 2790 3870 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07028 410 2790 3871 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07029 5182 3873 3872 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07030 3873 3872 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07031 411 2790 3872 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07032 409 2790 3873 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07033 5182 3875 3874 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07034 3875 3874 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07035 412 2791 3874 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07036 410 2791 3875 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07037 5182 3877 3876 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07038 3877 3876 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07039 411 2791 3876 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07040 409 2791 3877 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07041 5182 3879 3878 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07042 3879 3878 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07043 412 2789 3878 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07044 410 2789 3879 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07045 5182 3881 3880 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07046 3881 3880 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07047 411 2789 3880 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07048 409 2789 3881 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07049 5182 3883 3882 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07050 3883 3882 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07051 412 2808 3882 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07052 410 2808 3883 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07053 5182 3885 3884 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07054 3885 3884 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07055 411 2808 3884 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07056 409 2808 3885 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07057 5182 3887 3886 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07058 3887 3886 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07059 412 2806 3886 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07060 410 2806 3887 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07061 5182 3889 3888 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07062 3889 3888 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07063 411 2806 3888 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07064 409 2806 3889 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07065 5182 3891 3890 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07066 3891 3890 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07067 412 2807 3890 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07068 410 2807 3891 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07069 5182 3893 3892 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07070 3893 3892 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07071 411 2807 3892 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07072 409 2807 3893 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07073 5182 3895 3894 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07074 3895 3894 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07075 412 2805 3894 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07076 410 2805 3895 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07077 5182 3897 3896 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07078 3897 3896 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07079 411 2805 3896 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07080 409 2805 3897 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07081 5182 3899 3898 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07082 3899 3898 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07083 412 2824 3898 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07084 410 2824 3899 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07085 5182 3901 3900 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07086 3901 3900 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07087 411 2824 3900 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07088 409 2824 3901 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07089 5182 3903 3902 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07090 3903 3902 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07091 412 2822 3902 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07092 410 2822 3903 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07093 5182 3905 3904 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07094 3905 3904 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07095 411 2822 3904 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07096 409 2822 3905 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07097 5182 3907 3906 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07098 3907 3906 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07099 412 2823 3906 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07100 410 2823 3907 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07101 5182 3909 3908 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07102 3909 3908 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07103 411 2823 3908 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07104 409 2823 3909 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07105 5182 3911 3910 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07106 3911 3910 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07107 412 2821 3910 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07108 410 2821 3911 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07109 5182 3913 3912 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07110 3913 3912 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07111 411 2821 3912 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07112 409 2821 3913 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07113 5182 3915 3914 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07114 3915 3914 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07115 412 2840 3914 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07116 410 2840 3915 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07117 5182 3917 3916 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07118 3917 3916 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07119 411 2840 3916 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07120 409 2840 3917 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07121 5182 3919 3918 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07122 3919 3918 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07123 412 2838 3918 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07124 410 2838 3919 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07125 5182 3921 3920 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07126 3921 3920 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07127 411 2838 3920 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07128 409 2838 3921 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07129 5182 3923 3922 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07130 3923 3922 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07131 412 2839 3922 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07132 410 2839 3923 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07133 5182 3925 3924 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07134 3925 3924 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07135 411 2839 3924 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07136 409 2839 3925 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07137 5182 3927 3926 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07138 3927 3926 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07139 412 2837 3926 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07140 410 2837 3927 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07141 5182 3929 3928 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07142 3929 3928 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07143 411 2837 3928 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07144 409 2837 3929 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07145 5182 3931 3930 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07146 3931 3930 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07147 412 2856 3930 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07148 410 2856 3931 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07149 5182 3933 3932 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07150 3933 3932 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07151 411 2856 3932 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07152 409 2856 3933 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07153 5182 3935 3934 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07154 3935 3934 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07155 412 2854 3934 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07156 410 2854 3935 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07157 5182 3937 3936 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07158 3937 3936 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07159 411 2854 3936 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07160 409 2854 3937 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07161 5182 3939 3938 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07162 3939 3938 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07163 412 2855 3938 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07164 410 2855 3939 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07165 5182 3941 3940 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07166 3941 3940 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07167 411 2855 3940 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07168 409 2855 3941 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07169 5182 3943 3942 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07170 3943 3942 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07171 412 2853 3942 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07172 410 2853 3943 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07173 5182 3945 3944 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07174 3945 3944 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07175 411 2853 3944 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07176 409 2853 3945 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07177 5182 3947 3946 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07178 3947 3946 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07179 412 2872 3946 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07180 410 2872 3947 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07181 5182 3949 3948 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07182 3949 3948 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07183 411 2872 3948 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07184 409 2872 3949 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07185 5182 3951 3950 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07186 3951 3950 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07187 412 2870 3950 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07188 410 2870 3951 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07189 5182 3953 3952 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07190 3953 3952 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07191 411 2870 3952 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07192 409 2870 3953 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07193 5182 3955 3954 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07194 3955 3954 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07195 412 2871 3954 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07196 410 2871 3955 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07197 5182 3957 3956 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07198 3957 3956 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07199 411 2871 3956 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07200 409 2871 3957 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07201 5182 3959 3958 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07202 3959 3958 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07203 412 2869 3958 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07204 410 2869 3959 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07205 5182 3961 3960 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07206 3961 3960 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07207 411 2869 3960 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07208 409 2869 3961 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07209 5182 3963 3962 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07210 3963 3962 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07211 412 2888 3962 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07212 410 2888 3963 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07213 5182 3965 3964 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07214 3965 3964 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07215 411 2888 3964 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07216 409 2888 3965 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07217 5182 3967 3966 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07218 3967 3966 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07219 412 2886 3966 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07220 410 2886 3967 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07221 5182 3969 3968 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07222 3969 3968 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07223 411 2886 3968 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07224 409 2886 3969 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07225 5182 3971 3970 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07226 3971 3970 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07227 412 2887 3970 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07228 410 2887 3971 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07229 5182 3973 3972 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07230 3973 3972 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07231 411 2887 3972 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07232 409 2887 3973 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07233 5182 3975 3974 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07234 3975 3974 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07235 412 2885 3974 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07236 410 2885 3975 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07237 5182 3977 3976 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07238 3977 3976 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07239 411 2885 3976 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07240 409 2885 3977 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07241 5182 3979 3978 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07242 3979 3978 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07243 412 2904 3978 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07244 410 2904 3979 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07245 5182 3981 3980 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07246 3981 3980 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07247 411 2904 3980 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07248 409 2904 3981 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07249 5182 3983 3982 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07250 3983 3982 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07251 412 2902 3982 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07252 410 2902 3983 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07253 5182 3985 3984 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07254 3985 3984 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07255 411 2902 3984 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07256 409 2902 3985 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07257 5182 3987 3986 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07258 3987 3986 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07259 412 2903 3986 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07260 410 2903 3987 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07261 5182 3989 3988 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07262 3989 3988 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07263 411 2903 3988 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07264 409 2903 3989 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07265 5182 3991 3990 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07266 3991 3990 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07267 412 2901 3990 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07268 410 2901 3991 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07269 5182 3993 3992 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07270 3993 3992 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07271 411 2901 3992 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07272 409 2901 3993 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07273 5182 3995 3994 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07274 3995 3994 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07275 412 2920 3994 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07276 410 2920 3995 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07277 5182 3997 3996 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07278 3997 3996 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07279 411 2920 3996 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07280 409 2920 3997 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07281 5182 3999 3998 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07282 3999 3998 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07283 412 2918 3998 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07284 410 2918 3999 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07285 5182 4001 4000 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07286 4001 4000 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07287 411 2918 4000 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07288 409 2918 4001 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07289 5182 4003 4002 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07290 4003 4002 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07291 412 2919 4002 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07292 410 2919 4003 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07293 5182 4005 4004 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07294 4005 4004 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07295 411 2919 4004 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07296 409 2919 4005 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07297 5182 4007 4006 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07298 4007 4006 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07299 412 2917 4006 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07300 410 2917 4007 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07301 5182 4009 4008 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07302 4009 4008 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07303 411 2917 4008 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07304 409 2917 4009 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07305 5182 4011 4010 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07306 4011 4010 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07307 412 2936 4010 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07308 410 2936 4011 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07309 5182 4013 4012 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07310 4013 4012 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07311 411 2936 4012 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07312 409 2936 4013 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07313 5182 4015 4014 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07314 4015 4014 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07315 412 2934 4014 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07316 410 2934 4015 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07317 5182 4017 4016 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07318 4017 4016 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07319 411 2934 4016 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07320 409 2934 4017 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07321 5182 4019 4018 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07322 4019 4018 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07323 412 2935 4018 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07324 410 2935 4019 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07325 5182 4021 4020 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07326 4021 4020 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07327 411 2935 4020 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07328 409 2935 4021 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07329 5182 4023 4022 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07330 4023 4022 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07331 412 2933 4022 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07332 410 2933 4023 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07333 5182 4025 4024 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07334 4025 4024 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07335 411 2933 4024 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07336 409 2933 4025 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07337 5182 4027 4026 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07338 4027 4026 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07339 412 2952 4026 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07340 410 2952 4027 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07341 5182 4029 4028 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07342 4029 4028 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07343 411 2952 4028 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07344 409 2952 4029 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07345 5182 4031 4030 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07346 4031 4030 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07347 412 2950 4030 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07348 410 2950 4031 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07349 5182 4033 4032 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07350 4033 4032 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07351 411 2950 4032 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07352 409 2950 4033 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07353 5182 4035 4034 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07354 4035 4034 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07355 412 2951 4034 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07356 410 2951 4035 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07357 5182 4037 4036 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07358 4037 4036 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07359 411 2951 4036 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07360 409 2951 4037 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07361 5182 4039 4038 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07362 4039 4038 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07363 412 2949 4038 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07364 410 2949 4039 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07365 5182 4041 4040 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07366 4041 4040 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07367 411 2949 4040 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07368 409 2949 4041 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07369 5182 4043 4042 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07370 4043 4042 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07371 412 2968 4042 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07372 410 2968 4043 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07373 5182 4045 4044 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07374 4045 4044 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07375 411 2968 4044 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07376 409 2968 4045 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07377 5182 4047 4046 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07378 4047 4046 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07379 412 2966 4046 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07380 410 2966 4047 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07381 5182 4049 4048 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07382 4049 4048 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07383 411 2966 4048 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07384 409 2966 4049 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07385 5182 4051 4050 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07386 4051 4050 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07387 412 2967 4050 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07388 410 2967 4051 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07389 5182 4053 4052 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07390 4053 4052 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07391 411 2967 4052 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07392 409 2967 4053 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07393 5182 4055 4054 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07394 4055 4054 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07395 412 2965 4054 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07396 410 2965 4055 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07397 5182 4057 4056 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07398 4057 4056 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07399 411 2965 4056 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07400 409 2965 4057 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07401 5182 4059 4058 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07402 4059 4058 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07403 412 2984 4058 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07404 410 2984 4059 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07405 5182 4061 4060 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07406 4061 4060 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07407 411 2984 4060 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07408 409 2984 4061 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07409 5182 4063 4062 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07410 4063 4062 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07411 412 2982 4062 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07412 410 2982 4063 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07413 5182 4065 4064 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07414 4065 4064 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07415 411 2982 4064 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07416 409 2982 4065 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07417 5182 4067 4066 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07418 4067 4066 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07419 412 2983 4066 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07420 410 2983 4067 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07421 5182 4069 4068 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07422 4069 4068 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07423 411 2983 4068 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07424 409 2983 4069 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07425 5182 4071 4070 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07426 4071 4070 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07427 412 2981 4070 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07428 410 2981 4071 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07429 5182 4073 4072 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07430 4073 4072 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07431 411 2981 4072 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07432 409 2981 4073 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07433 5182 4075 4074 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07434 4075 4074 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07435 412 3000 4074 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07436 410 3000 4075 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07437 5182 4077 4076 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07438 4077 4076 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07439 411 3000 4076 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07440 409 3000 4077 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07441 5182 4079 4078 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07442 4079 4078 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07443 412 2998 4078 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07444 410 2998 4079 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07445 5182 4081 4080 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07446 4081 4080 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07447 411 2998 4080 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07448 409 2998 4081 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07449 5182 4083 4082 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07450 4083 4082 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07451 412 2999 4082 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07452 410 2999 4083 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07453 5182 4085 4084 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07454 4085 4084 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07455 411 2999 4084 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07456 409 2999 4085 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07457 5182 4087 4086 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07458 4087 4086 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07459 412 2997 4086 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07460 410 2997 4087 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07461 5182 4089 4088 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07462 4089 4088 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07463 411 2997 4088 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07464 409 2997 4089 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07465 5182 4091 4090 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07466 4091 4090 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07467 412 3016 4090 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07468 410 3016 4091 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07469 5182 4093 4092 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07470 4093 4092 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07471 411 3016 4092 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07472 409 3016 4093 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07473 5182 4095 4094 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07474 4095 4094 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07475 412 3014 4094 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07476 410 3014 4095 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07477 5182 4097 4096 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07478 4097 4096 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07479 411 3014 4096 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07480 409 3014 4097 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07481 5182 4099 4098 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07482 4099 4098 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07483 412 3015 4098 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07484 410 3015 4099 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07485 5182 4101 4100 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07486 4101 4100 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07487 411 3015 4100 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07488 409 3015 4101 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07489 5182 4103 4102 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07490 4103 4102 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07491 412 3013 4102 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07492 410 3013 4103 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07493 5182 4105 4104 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07494 4105 4104 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07495 411 3013 4104 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07496 409 3013 4105 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07497 5182 4107 4106 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07498 4107 4106 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07499 412 3032 4106 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07500 410 3032 4107 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07501 5182 4109 4108 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07502 4109 4108 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07503 411 3032 4108 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07504 409 3032 4109 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07505 5182 4111 4110 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07506 4111 4110 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07507 412 3030 4110 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07508 410 3030 4111 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07509 5182 4113 4112 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07510 4113 4112 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07511 411 3030 4112 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07512 409 3030 4113 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07513 5182 4115 4114 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07514 4115 4114 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07515 412 3031 4114 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07516 410 3031 4115 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07517 5182 4117 4116 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07518 4117 4116 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07519 411 3031 4116 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07520 409 3031 4117 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07521 5182 4119 4118 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07522 4119 4118 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07523 412 3029 4118 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07524 410 3029 4119 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07525 5182 4121 4120 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07526 4121 4120 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07527 411 3029 4120 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07528 409 3029 4121 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07529 409 3045 416 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_07530 416 3046 410 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_07531 411 3045 417 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_07532 417 3046 412 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_07533 4125 3081 4123 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_07534 4130 4125 413 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_07535 413 5176 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_07536 413 4123 4122 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_07537 5182 5176 414 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_07538 4124 417 414 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_07539 414 416 4123 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_07540 4125 417 415 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_07541 415 5176 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_07542 415 416 4126 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_07543 5183 3081 417 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_07544 417 3081 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_07545 5183 3081 416 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_07546 416 3081 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_07547 4127 5179 417 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_07548 416 5179 4128 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_07549 417 3081 416 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_07550 5182 5187 4127 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_07551 4128 4129 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_07552 4127 5187 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_07553 5182 4129 4128 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_07554 5182 5187 4129 5182 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_07555 5187 4131 5182 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_07556 5182 4131 5187 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_07557 5182 5179 4131 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_07558 4131 4130 5182 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_07559 4131 5176 4132 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_07560 421 2528 419 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07561 421 2528 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_07562 419 2528 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_07563 420 2528 418 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07564 5183 2528 420 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_07565 5183 2528 418 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_07566 5182 4134 4133 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07567 4134 4133 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07568 421 2536 4133 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07569 419 2536 4134 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07570 5182 4136 4135 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07571 4136 4135 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07572 420 2536 4135 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07573 418 2536 4136 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07574 5182 4138 4137 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07575 4138 4137 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07576 421 2534 4137 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07577 419 2534 4138 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07578 5182 4140 4139 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07579 4140 4139 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07580 420 2534 4139 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07581 418 2534 4140 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07582 5182 4142 4141 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07583 4142 4141 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07584 421 2535 4141 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07585 419 2535 4142 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07586 5182 4144 4143 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07587 4144 4143 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07588 420 2535 4143 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07589 418 2535 4144 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07590 5182 4146 4145 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07591 4146 4145 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07592 421 2533 4145 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07593 419 2533 4146 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07594 5182 4148 4147 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07595 4148 4147 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07596 420 2533 4147 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07597 418 2533 4148 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07598 5182 4150 4149 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07599 4150 4149 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07600 421 2552 4149 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07601 419 2552 4150 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07602 5182 4152 4151 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07603 4152 4151 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07604 420 2552 4151 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07605 418 2552 4152 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07606 5182 4154 4153 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07607 4154 4153 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07608 421 2550 4153 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07609 419 2550 4154 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07610 5182 4156 4155 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07611 4156 4155 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07612 420 2550 4155 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07613 418 2550 4156 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07614 5182 4158 4157 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07615 4158 4157 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07616 421 2551 4157 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07617 419 2551 4158 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07618 5182 4160 4159 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07619 4160 4159 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07620 420 2551 4159 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07621 418 2551 4160 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07622 5182 4162 4161 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07623 4162 4161 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07624 421 2549 4161 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07625 419 2549 4162 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07626 5182 4164 4163 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07627 4164 4163 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07628 420 2549 4163 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07629 418 2549 4164 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07630 5182 4166 4165 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07631 4166 4165 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07632 421 2568 4165 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07633 419 2568 4166 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07634 5182 4168 4167 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07635 4168 4167 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07636 420 2568 4167 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07637 418 2568 4168 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07638 5182 4170 4169 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07639 4170 4169 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07640 421 2566 4169 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07641 419 2566 4170 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07642 5182 4172 4171 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07643 4172 4171 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07644 420 2566 4171 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07645 418 2566 4172 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07646 5182 4174 4173 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07647 4174 4173 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07648 421 2567 4173 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07649 419 2567 4174 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07650 5182 4176 4175 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07651 4176 4175 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07652 420 2567 4175 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07653 418 2567 4176 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07654 5182 4178 4177 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07655 4178 4177 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07656 421 2565 4177 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07657 419 2565 4178 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07658 5182 4180 4179 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07659 4180 4179 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07660 420 2565 4179 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07661 418 2565 4180 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07662 5182 4182 4181 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07663 4182 4181 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07664 421 2584 4181 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07665 419 2584 4182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07666 5182 4184 4183 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07667 4184 4183 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07668 420 2584 4183 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07669 418 2584 4184 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07670 5182 4186 4185 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07671 4186 4185 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07672 421 2582 4185 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07673 419 2582 4186 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07674 5182 4188 4187 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07675 4188 4187 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07676 420 2582 4187 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07677 418 2582 4188 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07678 5182 4190 4189 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07679 4190 4189 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07680 421 2583 4189 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07681 419 2583 4190 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07682 5182 4192 4191 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07683 4192 4191 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07684 420 2583 4191 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07685 418 2583 4192 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07686 5182 4194 4193 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07687 4194 4193 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07688 421 2581 4193 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07689 419 2581 4194 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07690 5182 4196 4195 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07691 4196 4195 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07692 420 2581 4195 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07693 418 2581 4196 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07694 5182 4198 4197 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07695 4198 4197 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07696 421 2600 4197 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07697 419 2600 4198 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07698 5182 4200 4199 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07699 4200 4199 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07700 420 2600 4199 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07701 418 2600 4200 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07702 5182 4202 4201 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07703 4202 4201 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07704 421 2598 4201 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07705 419 2598 4202 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07706 5182 4204 4203 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07707 4204 4203 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07708 420 2598 4203 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07709 418 2598 4204 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07710 5182 4206 4205 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07711 4206 4205 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07712 421 2599 4205 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07713 419 2599 4206 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07714 5182 4208 4207 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07715 4208 4207 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07716 420 2599 4207 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07717 418 2599 4208 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07718 5182 4210 4209 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07719 4210 4209 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07720 421 2597 4209 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07721 419 2597 4210 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07722 5182 4212 4211 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07723 4212 4211 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07724 420 2597 4211 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07725 418 2597 4212 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07726 5182 4214 4213 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07727 4214 4213 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07728 421 2616 4213 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07729 419 2616 4214 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07730 5182 4216 4215 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07731 4216 4215 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07732 420 2616 4215 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07733 418 2616 4216 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07734 5182 4218 4217 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07735 4218 4217 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07736 421 2614 4217 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07737 419 2614 4218 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07738 5182 4220 4219 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07739 4220 4219 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07740 420 2614 4219 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07741 418 2614 4220 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07742 5182 4222 4221 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07743 4222 4221 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07744 421 2615 4221 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07745 419 2615 4222 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07746 5182 4224 4223 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07747 4224 4223 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07748 420 2615 4223 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07749 418 2615 4224 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07750 5182 4226 4225 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07751 4226 4225 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07752 421 2613 4225 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07753 419 2613 4226 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07754 5182 4228 4227 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07755 4228 4227 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07756 420 2613 4227 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07757 418 2613 4228 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07758 5182 4230 4229 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07759 4230 4229 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07760 421 2632 4229 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07761 419 2632 4230 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07762 5182 4232 4231 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07763 4232 4231 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07764 420 2632 4231 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07765 418 2632 4232 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07766 5182 4234 4233 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07767 4234 4233 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07768 421 2630 4233 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07769 419 2630 4234 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07770 5182 4236 4235 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07771 4236 4235 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07772 420 2630 4235 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07773 418 2630 4236 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07774 5182 4238 4237 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07775 4238 4237 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07776 421 2631 4237 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07777 419 2631 4238 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07778 5182 4240 4239 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07779 4240 4239 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07780 420 2631 4239 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07781 418 2631 4240 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07782 5182 4242 4241 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07783 4242 4241 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07784 421 2629 4241 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07785 419 2629 4242 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07786 5182 4244 4243 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07787 4244 4243 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07788 420 2629 4243 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07789 418 2629 4244 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07790 5182 4246 4245 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07791 4246 4245 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07792 421 2648 4245 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07793 419 2648 4246 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07794 5182 4248 4247 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07795 4248 4247 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07796 420 2648 4247 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07797 418 2648 4248 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07798 5182 4250 4249 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07799 4250 4249 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07800 421 2646 4249 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07801 419 2646 4250 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07802 5182 4252 4251 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07803 4252 4251 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07804 420 2646 4251 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07805 418 2646 4252 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07806 5182 4254 4253 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07807 4254 4253 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07808 421 2647 4253 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07809 419 2647 4254 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07810 5182 4256 4255 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07811 4256 4255 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07812 420 2647 4255 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07813 418 2647 4256 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07814 5182 4258 4257 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07815 4258 4257 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07816 421 2645 4257 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07817 419 2645 4258 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07818 5182 4260 4259 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07819 4260 4259 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07820 420 2645 4259 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07821 418 2645 4260 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07822 5182 4262 4261 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07823 4262 4261 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07824 421 2664 4261 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07825 419 2664 4262 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07826 5182 4264 4263 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07827 4264 4263 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07828 420 2664 4263 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07829 418 2664 4264 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07830 5182 4266 4265 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07831 4266 4265 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07832 421 2662 4265 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07833 419 2662 4266 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07834 5182 4268 4267 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07835 4268 4267 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07836 420 2662 4267 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07837 418 2662 4268 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07838 5182 4270 4269 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07839 4270 4269 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07840 421 2663 4269 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07841 419 2663 4270 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07842 5182 4272 4271 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07843 4272 4271 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07844 420 2663 4271 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07845 418 2663 4272 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07846 5182 4274 4273 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07847 4274 4273 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07848 421 2661 4273 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07849 419 2661 4274 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07850 5182 4276 4275 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07851 4276 4275 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07852 420 2661 4275 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07853 418 2661 4276 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07854 5182 4278 4277 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07855 4278 4277 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07856 421 2680 4277 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07857 419 2680 4278 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07858 5182 4280 4279 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07859 4280 4279 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07860 420 2680 4279 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07861 418 2680 4280 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07862 5182 4282 4281 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07863 4282 4281 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07864 421 2678 4281 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07865 419 2678 4282 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07866 5182 4284 4283 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07867 4284 4283 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07868 420 2678 4283 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07869 418 2678 4284 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07870 5182 4286 4285 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07871 4286 4285 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07872 421 2679 4285 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07873 419 2679 4286 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07874 5182 4288 4287 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07875 4288 4287 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07876 420 2679 4287 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07877 418 2679 4288 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07878 5182 4290 4289 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07879 4290 4289 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07880 421 2677 4289 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07881 419 2677 4290 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07882 5182 4292 4291 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07883 4292 4291 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07884 420 2677 4291 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07885 418 2677 4292 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07886 5182 4294 4293 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07887 4294 4293 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07888 421 2696 4293 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07889 419 2696 4294 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07890 5182 4296 4295 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07891 4296 4295 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07892 420 2696 4295 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07893 418 2696 4296 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07894 5182 4298 4297 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07895 4298 4297 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07896 421 2694 4297 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07897 419 2694 4298 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07898 5182 4300 4299 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07899 4300 4299 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07900 420 2694 4299 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07901 418 2694 4300 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07902 5182 4302 4301 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07903 4302 4301 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07904 421 2695 4301 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07905 419 2695 4302 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07906 5182 4304 4303 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07907 4304 4303 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07908 420 2695 4303 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07909 418 2695 4304 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07910 5182 4306 4305 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07911 4306 4305 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07912 421 2693 4305 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07913 419 2693 4306 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07914 5182 4308 4307 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07915 4308 4307 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07916 420 2693 4307 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07917 418 2693 4308 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07918 5182 4310 4309 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07919 4310 4309 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07920 421 2712 4309 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07921 419 2712 4310 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07922 5182 4312 4311 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07923 4312 4311 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07924 420 2712 4311 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07925 418 2712 4312 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07926 5182 4314 4313 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07927 4314 4313 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07928 421 2710 4313 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07929 419 2710 4314 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07930 5182 4316 4315 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07931 4316 4315 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07932 420 2710 4315 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07933 418 2710 4316 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07934 5182 4318 4317 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07935 4318 4317 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07936 421 2711 4317 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07937 419 2711 4318 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07938 5182 4320 4319 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07939 4320 4319 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07940 420 2711 4319 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07941 418 2711 4320 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07942 5182 4322 4321 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07943 4322 4321 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07944 421 2709 4321 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07945 419 2709 4322 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07946 5182 4324 4323 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07947 4324 4323 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07948 420 2709 4323 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07949 418 2709 4324 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07950 5182 4326 4325 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07951 4326 4325 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07952 421 2728 4325 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07953 419 2728 4326 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07954 5182 4328 4327 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07955 4328 4327 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07956 420 2728 4327 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07957 418 2728 4328 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07958 5182 4330 4329 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07959 4330 4329 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07960 421 2726 4329 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07961 419 2726 4330 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07962 5182 4332 4331 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07963 4332 4331 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07964 420 2726 4331 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07965 418 2726 4332 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07966 5182 4334 4333 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07967 4334 4333 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07968 421 2727 4333 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07969 419 2727 4334 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07970 5182 4336 4335 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07971 4336 4335 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07972 420 2727 4335 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07973 418 2727 4336 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07974 5182 4338 4337 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07975 4338 4337 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07976 421 2725 4337 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07977 419 2725 4338 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07978 5182 4340 4339 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07979 4340 4339 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07980 420 2725 4339 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07981 418 2725 4340 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07982 5182 4342 4341 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07983 4342 4341 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07984 421 2744 4341 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07985 419 2744 4342 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07986 5182 4344 4343 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07987 4344 4343 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07988 420 2744 4343 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07989 418 2744 4344 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07990 5182 4346 4345 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07991 4346 4345 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07992 421 2742 4345 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07993 419 2742 4346 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07994 5182 4348 4347 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07995 4348 4347 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07996 420 2742 4347 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07997 418 2742 4348 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07998 5182 4350 4349 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_07999 4350 4349 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08000 421 2743 4349 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08001 419 2743 4350 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08002 5182 4352 4351 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08003 4352 4351 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08004 420 2743 4351 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08005 418 2743 4352 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08006 5182 4354 4353 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08007 4354 4353 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08008 421 2741 4353 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08009 419 2741 4354 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08010 5182 4356 4355 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08011 4356 4355 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08012 420 2741 4355 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08013 418 2741 4356 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08014 5182 4358 4357 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08015 4358 4357 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08016 421 2760 4357 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08017 419 2760 4358 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08018 5182 4360 4359 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08019 4360 4359 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08020 420 2760 4359 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08021 418 2760 4360 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08022 5182 4362 4361 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08023 4362 4361 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08024 421 2758 4361 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08025 419 2758 4362 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08026 5182 4364 4363 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08027 4364 4363 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08028 420 2758 4363 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08029 418 2758 4364 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08030 5182 4366 4365 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08031 4366 4365 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08032 421 2759 4365 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08033 419 2759 4366 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08034 5182 4368 4367 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08035 4368 4367 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08036 420 2759 4367 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08037 418 2759 4368 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08038 5182 4370 4369 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08039 4370 4369 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08040 421 2757 4369 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08041 419 2757 4370 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08042 5182 4372 4371 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08043 4372 4371 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08044 420 2757 4371 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08045 418 2757 4372 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08046 5182 4374 4373 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08047 4374 4373 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08048 421 2776 4373 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08049 419 2776 4374 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08050 5182 4376 4375 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08051 4376 4375 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08052 420 2776 4375 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08053 418 2776 4376 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08054 5182 4378 4377 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08055 4378 4377 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08056 421 2774 4377 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08057 419 2774 4378 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08058 5182 4380 4379 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08059 4380 4379 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08060 420 2774 4379 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08061 418 2774 4380 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08062 5182 4382 4381 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08063 4382 4381 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08064 421 2775 4381 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08065 419 2775 4382 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08066 5182 4384 4383 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08067 4384 4383 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08068 420 2775 4383 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08069 418 2775 4384 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08070 5182 4386 4385 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08071 4386 4385 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08072 421 2773 4385 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08073 419 2773 4386 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08074 5182 4388 4387 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08075 4388 4387 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08076 420 2773 4387 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08077 418 2773 4388 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08078 5182 4390 4389 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08079 4390 4389 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08080 421 2792 4389 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08081 419 2792 4390 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08082 5182 4392 4391 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08083 4392 4391 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08084 420 2792 4391 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08085 418 2792 4392 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08086 5182 4394 4393 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08087 4394 4393 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08088 421 2790 4393 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08089 419 2790 4394 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08090 5182 4396 4395 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08091 4396 4395 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08092 420 2790 4395 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08093 418 2790 4396 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08094 5182 4398 4397 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08095 4398 4397 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08096 421 2791 4397 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08097 419 2791 4398 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08098 5182 4400 4399 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08099 4400 4399 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08100 420 2791 4399 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08101 418 2791 4400 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08102 5182 4402 4401 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08103 4402 4401 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08104 421 2789 4401 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08105 419 2789 4402 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08106 5182 4404 4403 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08107 4404 4403 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08108 420 2789 4403 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08109 418 2789 4404 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08110 5182 4406 4405 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08111 4406 4405 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08112 421 2808 4405 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08113 419 2808 4406 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08114 5182 4408 4407 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08115 4408 4407 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08116 420 2808 4407 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08117 418 2808 4408 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08118 5182 4410 4409 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08119 4410 4409 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08120 421 2806 4409 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08121 419 2806 4410 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08122 5182 4412 4411 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08123 4412 4411 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08124 420 2806 4411 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08125 418 2806 4412 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08126 5182 4414 4413 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08127 4414 4413 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08128 421 2807 4413 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08129 419 2807 4414 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08130 5182 4416 4415 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08131 4416 4415 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08132 420 2807 4415 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08133 418 2807 4416 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08134 5182 4418 4417 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08135 4418 4417 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08136 421 2805 4417 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08137 419 2805 4418 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08138 5182 4420 4419 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08139 4420 4419 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08140 420 2805 4419 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08141 418 2805 4420 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08142 5182 4422 4421 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08143 4422 4421 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08144 421 2824 4421 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08145 419 2824 4422 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08146 5182 4424 4423 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08147 4424 4423 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08148 420 2824 4423 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08149 418 2824 4424 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08150 5182 4426 4425 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08151 4426 4425 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08152 421 2822 4425 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08153 419 2822 4426 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08154 5182 4428 4427 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08155 4428 4427 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08156 420 2822 4427 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08157 418 2822 4428 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08158 5182 4430 4429 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08159 4430 4429 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08160 421 2823 4429 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08161 419 2823 4430 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08162 5182 4432 4431 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08163 4432 4431 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08164 420 2823 4431 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08165 418 2823 4432 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08166 5182 4434 4433 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08167 4434 4433 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08168 421 2821 4433 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08169 419 2821 4434 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08170 5182 4436 4435 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08171 4436 4435 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08172 420 2821 4435 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08173 418 2821 4436 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08174 5182 4438 4437 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08175 4438 4437 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08176 421 2840 4437 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08177 419 2840 4438 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08178 5182 4440 4439 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08179 4440 4439 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08180 420 2840 4439 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08181 418 2840 4440 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08182 5182 4442 4441 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08183 4442 4441 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08184 421 2838 4441 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08185 419 2838 4442 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08186 5182 4444 4443 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08187 4444 4443 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08188 420 2838 4443 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08189 418 2838 4444 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08190 5182 4446 4445 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08191 4446 4445 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08192 421 2839 4445 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08193 419 2839 4446 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08194 5182 4448 4447 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08195 4448 4447 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08196 420 2839 4447 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08197 418 2839 4448 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08198 5182 4450 4449 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08199 4450 4449 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08200 421 2837 4449 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08201 419 2837 4450 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08202 5182 4452 4451 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08203 4452 4451 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08204 420 2837 4451 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08205 418 2837 4452 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08206 5182 4454 4453 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08207 4454 4453 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08208 421 2856 4453 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08209 419 2856 4454 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08210 5182 4456 4455 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08211 4456 4455 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08212 420 2856 4455 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08213 418 2856 4456 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08214 5182 4458 4457 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08215 4458 4457 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08216 421 2854 4457 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08217 419 2854 4458 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08218 5182 4460 4459 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08219 4460 4459 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08220 420 2854 4459 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08221 418 2854 4460 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08222 5182 4462 4461 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08223 4462 4461 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08224 421 2855 4461 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08225 419 2855 4462 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08226 5182 4464 4463 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08227 4464 4463 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08228 420 2855 4463 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08229 418 2855 4464 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08230 5182 4466 4465 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08231 4466 4465 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08232 421 2853 4465 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08233 419 2853 4466 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08234 5182 4468 4467 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08235 4468 4467 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08236 420 2853 4467 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08237 418 2853 4468 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08238 5182 4470 4469 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08239 4470 4469 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08240 421 2872 4469 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08241 419 2872 4470 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08242 5182 4472 4471 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08243 4472 4471 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08244 420 2872 4471 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08245 418 2872 4472 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08246 5182 4474 4473 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08247 4474 4473 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08248 421 2870 4473 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08249 419 2870 4474 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08250 5182 4476 4475 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08251 4476 4475 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08252 420 2870 4475 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08253 418 2870 4476 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08254 5182 4478 4477 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08255 4478 4477 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08256 421 2871 4477 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08257 419 2871 4478 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08258 5182 4480 4479 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08259 4480 4479 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08260 420 2871 4479 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08261 418 2871 4480 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08262 5182 4482 4481 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08263 4482 4481 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08264 421 2869 4481 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08265 419 2869 4482 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08266 5182 4484 4483 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08267 4484 4483 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08268 420 2869 4483 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08269 418 2869 4484 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08270 5182 4486 4485 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08271 4486 4485 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08272 421 2888 4485 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08273 419 2888 4486 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08274 5182 4488 4487 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08275 4488 4487 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08276 420 2888 4487 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08277 418 2888 4488 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08278 5182 4490 4489 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08279 4490 4489 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08280 421 2886 4489 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08281 419 2886 4490 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08282 5182 4492 4491 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08283 4492 4491 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08284 420 2886 4491 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08285 418 2886 4492 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08286 5182 4494 4493 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08287 4494 4493 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08288 421 2887 4493 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08289 419 2887 4494 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08290 5182 4496 4495 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08291 4496 4495 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08292 420 2887 4495 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08293 418 2887 4496 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08294 5182 4498 4497 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08295 4498 4497 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08296 421 2885 4497 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08297 419 2885 4498 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08298 5182 4500 4499 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08299 4500 4499 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08300 420 2885 4499 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08301 418 2885 4500 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08302 5182 4502 4501 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08303 4502 4501 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08304 421 2904 4501 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08305 419 2904 4502 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08306 5182 4504 4503 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08307 4504 4503 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08308 420 2904 4503 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08309 418 2904 4504 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08310 5182 4506 4505 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08311 4506 4505 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08312 421 2902 4505 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08313 419 2902 4506 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08314 5182 4508 4507 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08315 4508 4507 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08316 420 2902 4507 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08317 418 2902 4508 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08318 5182 4510 4509 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08319 4510 4509 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08320 421 2903 4509 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08321 419 2903 4510 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08322 5182 4512 4511 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08323 4512 4511 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08324 420 2903 4511 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08325 418 2903 4512 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08326 5182 4514 4513 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08327 4514 4513 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08328 421 2901 4513 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08329 419 2901 4514 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08330 5182 4516 4515 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08331 4516 4515 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08332 420 2901 4515 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08333 418 2901 4516 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08334 5182 4518 4517 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08335 4518 4517 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08336 421 2920 4517 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08337 419 2920 4518 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08338 5182 4520 4519 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08339 4520 4519 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08340 420 2920 4519 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08341 418 2920 4520 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08342 5182 4522 4521 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08343 4522 4521 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08344 421 2918 4521 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08345 419 2918 4522 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08346 5182 4524 4523 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08347 4524 4523 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08348 420 2918 4523 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08349 418 2918 4524 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08350 5182 4526 4525 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08351 4526 4525 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08352 421 2919 4525 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08353 419 2919 4526 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08354 5182 4528 4527 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08355 4528 4527 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08356 420 2919 4527 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08357 418 2919 4528 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08358 5182 4530 4529 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08359 4530 4529 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08360 421 2917 4529 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08361 419 2917 4530 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08362 5182 4532 4531 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08363 4532 4531 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08364 420 2917 4531 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08365 418 2917 4532 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08366 5182 4534 4533 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08367 4534 4533 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08368 421 2936 4533 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08369 419 2936 4534 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08370 5182 4536 4535 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08371 4536 4535 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08372 420 2936 4535 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08373 418 2936 4536 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08374 5182 4538 4537 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08375 4538 4537 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08376 421 2934 4537 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08377 419 2934 4538 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08378 5182 4540 4539 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08379 4540 4539 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08380 420 2934 4539 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08381 418 2934 4540 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08382 5182 4542 4541 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08383 4542 4541 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08384 421 2935 4541 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08385 419 2935 4542 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08386 5182 4544 4543 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08387 4544 4543 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08388 420 2935 4543 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08389 418 2935 4544 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08390 5182 4546 4545 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08391 4546 4545 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08392 421 2933 4545 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08393 419 2933 4546 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08394 5182 4548 4547 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08395 4548 4547 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08396 420 2933 4547 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08397 418 2933 4548 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08398 5182 4550 4549 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08399 4550 4549 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08400 421 2952 4549 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08401 419 2952 4550 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08402 5182 4552 4551 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08403 4552 4551 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08404 420 2952 4551 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08405 418 2952 4552 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08406 5182 4554 4553 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08407 4554 4553 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08408 421 2950 4553 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08409 419 2950 4554 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08410 5182 4556 4555 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08411 4556 4555 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08412 420 2950 4555 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08413 418 2950 4556 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08414 5182 4558 4557 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08415 4558 4557 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08416 421 2951 4557 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08417 419 2951 4558 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08418 5182 4560 4559 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08419 4560 4559 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08420 420 2951 4559 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08421 418 2951 4560 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08422 5182 4562 4561 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08423 4562 4561 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08424 421 2949 4561 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08425 419 2949 4562 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08426 5182 4564 4563 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08427 4564 4563 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08428 420 2949 4563 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08429 418 2949 4564 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08430 5182 4566 4565 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08431 4566 4565 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08432 421 2968 4565 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08433 419 2968 4566 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08434 5182 4568 4567 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08435 4568 4567 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08436 420 2968 4567 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08437 418 2968 4568 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08438 5182 4570 4569 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08439 4570 4569 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08440 421 2966 4569 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08441 419 2966 4570 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08442 5182 4572 4571 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08443 4572 4571 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08444 420 2966 4571 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08445 418 2966 4572 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08446 5182 4574 4573 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08447 4574 4573 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08448 421 2967 4573 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08449 419 2967 4574 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08450 5182 4576 4575 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08451 4576 4575 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08452 420 2967 4575 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08453 418 2967 4576 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08454 5182 4578 4577 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08455 4578 4577 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08456 421 2965 4577 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08457 419 2965 4578 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08458 5182 4580 4579 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08459 4580 4579 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08460 420 2965 4579 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08461 418 2965 4580 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08462 5182 4582 4581 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08463 4582 4581 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08464 421 2984 4581 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08465 419 2984 4582 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08466 5182 4584 4583 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08467 4584 4583 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08468 420 2984 4583 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08469 418 2984 4584 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08470 5182 4586 4585 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08471 4586 4585 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08472 421 2982 4585 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08473 419 2982 4586 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08474 5182 4588 4587 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08475 4588 4587 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08476 420 2982 4587 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08477 418 2982 4588 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08478 5182 4590 4589 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08479 4590 4589 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08480 421 2983 4589 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08481 419 2983 4590 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08482 5182 4592 4591 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08483 4592 4591 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08484 420 2983 4591 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08485 418 2983 4592 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08486 5182 4594 4593 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08487 4594 4593 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08488 421 2981 4593 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08489 419 2981 4594 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08490 5182 4596 4595 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08491 4596 4595 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08492 420 2981 4595 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08493 418 2981 4596 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08494 5182 4598 4597 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08495 4598 4597 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08496 421 3000 4597 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08497 419 3000 4598 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08498 5182 4600 4599 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08499 4600 4599 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08500 420 3000 4599 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08501 418 3000 4600 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08502 5182 4602 4601 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08503 4602 4601 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08504 421 2998 4601 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08505 419 2998 4602 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08506 5182 4604 4603 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08507 4604 4603 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08508 420 2998 4603 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08509 418 2998 4604 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08510 5182 4606 4605 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08511 4606 4605 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08512 421 2999 4605 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08513 419 2999 4606 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08514 5182 4608 4607 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08515 4608 4607 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08516 420 2999 4607 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08517 418 2999 4608 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08518 5182 4610 4609 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08519 4610 4609 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08520 421 2997 4609 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08521 419 2997 4610 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08522 5182 4612 4611 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08523 4612 4611 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08524 420 2997 4611 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08525 418 2997 4612 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08526 5182 4614 4613 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08527 4614 4613 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08528 421 3016 4613 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08529 419 3016 4614 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08530 5182 4616 4615 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08531 4616 4615 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08532 420 3016 4615 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08533 418 3016 4616 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08534 5182 4618 4617 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08535 4618 4617 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08536 421 3014 4617 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08537 419 3014 4618 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08538 5182 4620 4619 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08539 4620 4619 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08540 420 3014 4619 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08541 418 3014 4620 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08542 5182 4622 4621 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08543 4622 4621 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08544 421 3015 4621 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08545 419 3015 4622 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08546 5182 4624 4623 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08547 4624 4623 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08548 420 3015 4623 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08549 418 3015 4624 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08550 5182 4626 4625 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08551 4626 4625 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08552 421 3013 4625 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08553 419 3013 4626 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08554 5182 4628 4627 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08555 4628 4627 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08556 420 3013 4627 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08557 418 3013 4628 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08558 5182 4630 4629 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08559 4630 4629 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08560 421 3032 4629 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08561 419 3032 4630 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08562 5182 4632 4631 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08563 4632 4631 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08564 420 3032 4631 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08565 418 3032 4632 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08566 5182 4634 4633 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08567 4634 4633 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08568 421 3030 4633 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08569 419 3030 4634 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08570 5182 4636 4635 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08571 4636 4635 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08572 420 3030 4635 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08573 418 3030 4636 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08574 5182 4638 4637 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08575 4638 4637 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08576 421 3031 4637 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08577 419 3031 4638 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08578 5182 4640 4639 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08579 4640 4639 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08580 420 3031 4639 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08581 418 3031 4640 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08582 5182 4642 4641 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08583 4642 4641 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08584 421 3029 4641 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08585 419 3029 4642 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08586 5182 4644 4643 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08587 4644 4643 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08588 420 3029 4643 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08589 418 3029 4644 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08590 418 3045 425 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_08591 425 3046 419 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_08592 420 3045 426 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_08593 426 3046 421 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_08594 4648 3081 4646 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_08595 4653 4648 422 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_08596 422 5176 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_08597 422 4646 4645 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_08598 5182 5176 423 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_08599 4647 426 423 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_08600 423 425 4646 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_08601 4648 426 424 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_08602 424 5176 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_08603 424 425 4649 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_08604 5183 3081 426 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_08605 426 3081 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_08606 5183 3081 425 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_08607 425 3081 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_08608 4650 5179 426 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_08609 425 5179 4651 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_08610 426 3081 425 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_08611 5182 5186 4650 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_08612 4651 4652 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_08613 4650 5186 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_08614 5182 4652 4651 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_08615 5182 5186 4652 5182 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_08616 5186 4654 5182 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_08617 5182 4654 5186 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_08618 5182 5179 4654 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_08619 4654 4653 5182 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_08620 4654 5176 4655 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_08621 430 2528 428 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08622 430 2528 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_08623 428 2528 5183 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_08624 429 2528 427 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08625 5183 2528 429 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_08626 5183 2528 427 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_08627 5182 4657 4656 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08628 4657 4656 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08629 430 2536 4656 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08630 428 2536 4657 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08631 5182 4659 4658 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08632 4659 4658 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08633 429 2536 4658 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08634 427 2536 4659 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08635 5182 4661 4660 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08636 4661 4660 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08637 430 2534 4660 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08638 428 2534 4661 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08639 5182 4663 4662 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08640 4663 4662 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08641 429 2534 4662 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08642 427 2534 4663 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08643 5182 4665 4664 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08644 4665 4664 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08645 430 2535 4664 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08646 428 2535 4665 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08647 5182 4667 4666 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08648 4667 4666 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08649 429 2535 4666 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08650 427 2535 4667 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08651 5182 4669 4668 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08652 4669 4668 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08653 430 2533 4668 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08654 428 2533 4669 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08655 5182 4671 4670 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08656 4671 4670 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08657 429 2533 4670 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08658 427 2533 4671 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08659 5182 4673 4672 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08660 4673 4672 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08661 430 2552 4672 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08662 428 2552 4673 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08663 5182 4675 4674 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08664 4675 4674 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08665 429 2552 4674 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08666 427 2552 4675 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08667 5182 4677 4676 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08668 4677 4676 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08669 430 2550 4676 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08670 428 2550 4677 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08671 5182 4679 4678 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08672 4679 4678 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08673 429 2550 4678 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08674 427 2550 4679 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08675 5182 4681 4680 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08676 4681 4680 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08677 430 2551 4680 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08678 428 2551 4681 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08679 5182 4683 4682 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08680 4683 4682 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08681 429 2551 4682 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08682 427 2551 4683 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08683 5182 4685 4684 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08684 4685 4684 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08685 430 2549 4684 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08686 428 2549 4685 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08687 5182 4687 4686 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08688 4687 4686 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08689 429 2549 4686 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08690 427 2549 4687 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08691 5182 4689 4688 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08692 4689 4688 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08693 430 2568 4688 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08694 428 2568 4689 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08695 5182 4691 4690 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08696 4691 4690 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08697 429 2568 4690 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08698 427 2568 4691 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08699 5182 4693 4692 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08700 4693 4692 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08701 430 2566 4692 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08702 428 2566 4693 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08703 5182 4695 4694 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08704 4695 4694 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08705 429 2566 4694 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08706 427 2566 4695 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08707 5182 4697 4696 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08708 4697 4696 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08709 430 2567 4696 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08710 428 2567 4697 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08711 5182 4699 4698 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08712 4699 4698 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08713 429 2567 4698 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08714 427 2567 4699 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08715 5182 4701 4700 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08716 4701 4700 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08717 430 2565 4700 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08718 428 2565 4701 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08719 5182 4703 4702 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08720 4703 4702 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08721 429 2565 4702 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08722 427 2565 4703 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08723 5182 4705 4704 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08724 4705 4704 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08725 430 2584 4704 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08726 428 2584 4705 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08727 5182 4707 4706 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08728 4707 4706 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08729 429 2584 4706 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08730 427 2584 4707 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08731 5182 4709 4708 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08732 4709 4708 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08733 430 2582 4708 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08734 428 2582 4709 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08735 5182 4711 4710 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08736 4711 4710 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08737 429 2582 4710 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08738 427 2582 4711 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08739 5182 4713 4712 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08740 4713 4712 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08741 430 2583 4712 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08742 428 2583 4713 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08743 5182 4715 4714 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08744 4715 4714 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08745 429 2583 4714 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08746 427 2583 4715 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08747 5182 4717 4716 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08748 4717 4716 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08749 430 2581 4716 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08750 428 2581 4717 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08751 5182 4719 4718 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08752 4719 4718 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08753 429 2581 4718 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08754 427 2581 4719 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08755 5182 4721 4720 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08756 4721 4720 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08757 430 2600 4720 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08758 428 2600 4721 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08759 5182 4723 4722 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08760 4723 4722 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08761 429 2600 4722 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08762 427 2600 4723 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08763 5182 4725 4724 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08764 4725 4724 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08765 430 2598 4724 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08766 428 2598 4725 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08767 5182 4727 4726 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08768 4727 4726 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08769 429 2598 4726 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08770 427 2598 4727 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08771 5182 4729 4728 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08772 4729 4728 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08773 430 2599 4728 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08774 428 2599 4729 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08775 5182 4731 4730 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08776 4731 4730 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08777 429 2599 4730 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08778 427 2599 4731 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08779 5182 4733 4732 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08780 4733 4732 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08781 430 2597 4732 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08782 428 2597 4733 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08783 5182 4735 4734 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08784 4735 4734 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08785 429 2597 4734 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08786 427 2597 4735 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08787 5182 4737 4736 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08788 4737 4736 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08789 430 2616 4736 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08790 428 2616 4737 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08791 5182 4739 4738 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08792 4739 4738 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08793 429 2616 4738 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08794 427 2616 4739 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08795 5182 4741 4740 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08796 4741 4740 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08797 430 2614 4740 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08798 428 2614 4741 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08799 5182 4743 4742 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08800 4743 4742 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08801 429 2614 4742 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08802 427 2614 4743 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08803 5182 4745 4744 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08804 4745 4744 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08805 430 2615 4744 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08806 428 2615 4745 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08807 5182 4747 4746 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08808 4747 4746 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08809 429 2615 4746 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08810 427 2615 4747 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08811 5182 4749 4748 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08812 4749 4748 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08813 430 2613 4748 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08814 428 2613 4749 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08815 5182 4751 4750 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08816 4751 4750 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08817 429 2613 4750 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08818 427 2613 4751 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08819 5182 4753 4752 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08820 4753 4752 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08821 430 2632 4752 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08822 428 2632 4753 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08823 5182 4755 4754 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08824 4755 4754 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08825 429 2632 4754 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08826 427 2632 4755 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08827 5182 4757 4756 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08828 4757 4756 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08829 430 2630 4756 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08830 428 2630 4757 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08831 5182 4759 4758 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08832 4759 4758 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08833 429 2630 4758 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08834 427 2630 4759 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08835 5182 4761 4760 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08836 4761 4760 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08837 430 2631 4760 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08838 428 2631 4761 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08839 5182 4763 4762 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08840 4763 4762 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08841 429 2631 4762 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08842 427 2631 4763 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08843 5182 4765 4764 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08844 4765 4764 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08845 430 2629 4764 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08846 428 2629 4765 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08847 5182 4767 4766 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08848 4767 4766 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08849 429 2629 4766 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08850 427 2629 4767 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08851 5182 4769 4768 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08852 4769 4768 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08853 430 2648 4768 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08854 428 2648 4769 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08855 5182 4771 4770 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08856 4771 4770 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08857 429 2648 4770 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08858 427 2648 4771 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08859 5182 4773 4772 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08860 4773 4772 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08861 430 2646 4772 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08862 428 2646 4773 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08863 5182 4775 4774 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08864 4775 4774 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08865 429 2646 4774 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08866 427 2646 4775 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08867 5182 4777 4776 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08868 4777 4776 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08869 430 2647 4776 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08870 428 2647 4777 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08871 5182 4779 4778 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08872 4779 4778 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08873 429 2647 4778 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08874 427 2647 4779 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08875 5182 4781 4780 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08876 4781 4780 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08877 430 2645 4780 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08878 428 2645 4781 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08879 5182 4783 4782 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08880 4783 4782 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08881 429 2645 4782 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08882 427 2645 4783 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08883 5182 4785 4784 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08884 4785 4784 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08885 430 2664 4784 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08886 428 2664 4785 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08887 5182 4787 4786 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08888 4787 4786 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08889 429 2664 4786 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08890 427 2664 4787 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08891 5182 4789 4788 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08892 4789 4788 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08893 430 2662 4788 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08894 428 2662 4789 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08895 5182 4791 4790 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08896 4791 4790 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08897 429 2662 4790 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08898 427 2662 4791 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08899 5182 4793 4792 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08900 4793 4792 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08901 430 2663 4792 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08902 428 2663 4793 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08903 5182 4795 4794 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08904 4795 4794 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08905 429 2663 4794 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08906 427 2663 4795 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08907 5182 4797 4796 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08908 4797 4796 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08909 430 2661 4796 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08910 428 2661 4797 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08911 5182 4799 4798 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08912 4799 4798 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08913 429 2661 4798 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08914 427 2661 4799 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08915 5182 4801 4800 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08916 4801 4800 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08917 430 2680 4800 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08918 428 2680 4801 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08919 5182 4803 4802 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08920 4803 4802 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08921 429 2680 4802 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08922 427 2680 4803 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08923 5182 4805 4804 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08924 4805 4804 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08925 430 2678 4804 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08926 428 2678 4805 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08927 5182 4807 4806 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08928 4807 4806 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08929 429 2678 4806 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08930 427 2678 4807 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08931 5182 4809 4808 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08932 4809 4808 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08933 430 2679 4808 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08934 428 2679 4809 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08935 5182 4811 4810 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08936 4811 4810 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08937 429 2679 4810 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08938 427 2679 4811 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08939 5182 4813 4812 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08940 4813 4812 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08941 430 2677 4812 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08942 428 2677 4813 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08943 5182 4815 4814 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08944 4815 4814 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08945 429 2677 4814 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08946 427 2677 4815 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08947 5182 4817 4816 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08948 4817 4816 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08949 430 2696 4816 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08950 428 2696 4817 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08951 5182 4819 4818 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08952 4819 4818 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08953 429 2696 4818 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08954 427 2696 4819 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08955 5182 4821 4820 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08956 4821 4820 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08957 430 2694 4820 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08958 428 2694 4821 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08959 5182 4823 4822 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08960 4823 4822 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08961 429 2694 4822 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08962 427 2694 4823 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08963 5182 4825 4824 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08964 4825 4824 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08965 430 2695 4824 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08966 428 2695 4825 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08967 5182 4827 4826 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08968 4827 4826 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08969 429 2695 4826 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08970 427 2695 4827 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08971 5182 4829 4828 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08972 4829 4828 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08973 430 2693 4828 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08974 428 2693 4829 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08975 5182 4831 4830 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08976 4831 4830 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08977 429 2693 4830 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08978 427 2693 4831 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08979 5182 4833 4832 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08980 4833 4832 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08981 430 2712 4832 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08982 428 2712 4833 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08983 5182 4835 4834 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08984 4835 4834 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08985 429 2712 4834 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08986 427 2712 4835 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08987 5182 4837 4836 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08988 4837 4836 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08989 430 2710 4836 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08990 428 2710 4837 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08991 5182 4839 4838 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08992 4839 4838 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08993 429 2710 4838 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08994 427 2710 4839 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08995 5182 4841 4840 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08996 4841 4840 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08997 430 2711 4840 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08998 428 2711 4841 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_08999 5182 4843 4842 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09000 4843 4842 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09001 429 2711 4842 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09002 427 2711 4843 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09003 5182 4845 4844 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09004 4845 4844 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09005 430 2709 4844 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09006 428 2709 4845 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09007 5182 4847 4846 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09008 4847 4846 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09009 429 2709 4846 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09010 427 2709 4847 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09011 5182 4849 4848 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09012 4849 4848 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09013 430 2728 4848 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09014 428 2728 4849 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09015 5182 4851 4850 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09016 4851 4850 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09017 429 2728 4850 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09018 427 2728 4851 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09019 5182 4853 4852 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09020 4853 4852 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09021 430 2726 4852 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09022 428 2726 4853 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09023 5182 4855 4854 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09024 4855 4854 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09025 429 2726 4854 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09026 427 2726 4855 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09027 5182 4857 4856 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09028 4857 4856 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09029 430 2727 4856 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09030 428 2727 4857 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09031 5182 4859 4858 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09032 4859 4858 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09033 429 2727 4858 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09034 427 2727 4859 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09035 5182 4861 4860 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09036 4861 4860 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09037 430 2725 4860 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09038 428 2725 4861 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09039 5182 4863 4862 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09040 4863 4862 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09041 429 2725 4862 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09042 427 2725 4863 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09043 5182 4865 4864 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09044 4865 4864 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09045 430 2744 4864 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09046 428 2744 4865 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09047 5182 4867 4866 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09048 4867 4866 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09049 429 2744 4866 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09050 427 2744 4867 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09051 5182 4869 4868 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09052 4869 4868 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09053 430 2742 4868 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09054 428 2742 4869 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09055 5182 4871 4870 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09056 4871 4870 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09057 429 2742 4870 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09058 427 2742 4871 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09059 5182 4873 4872 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09060 4873 4872 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09061 430 2743 4872 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09062 428 2743 4873 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09063 5182 4875 4874 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09064 4875 4874 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09065 429 2743 4874 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09066 427 2743 4875 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09067 5182 4877 4876 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09068 4877 4876 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09069 430 2741 4876 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09070 428 2741 4877 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09071 5182 4879 4878 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09072 4879 4878 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09073 429 2741 4878 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09074 427 2741 4879 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09075 5182 4881 4880 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09076 4881 4880 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09077 430 2760 4880 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09078 428 2760 4881 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09079 5182 4883 4882 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09080 4883 4882 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09081 429 2760 4882 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09082 427 2760 4883 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09083 5182 4885 4884 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09084 4885 4884 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09085 430 2758 4884 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09086 428 2758 4885 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09087 5182 4887 4886 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09088 4887 4886 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09089 429 2758 4886 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09090 427 2758 4887 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09091 5182 4889 4888 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09092 4889 4888 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09093 430 2759 4888 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09094 428 2759 4889 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09095 5182 4891 4890 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09096 4891 4890 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09097 429 2759 4890 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09098 427 2759 4891 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09099 5182 4893 4892 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09100 4893 4892 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09101 430 2757 4892 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09102 428 2757 4893 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09103 5182 4895 4894 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09104 4895 4894 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09105 429 2757 4894 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09106 427 2757 4895 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09107 5182 4897 4896 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09108 4897 4896 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09109 430 2776 4896 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09110 428 2776 4897 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09111 5182 4899 4898 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09112 4899 4898 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09113 429 2776 4898 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09114 427 2776 4899 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09115 5182 4901 4900 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09116 4901 4900 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09117 430 2774 4900 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09118 428 2774 4901 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09119 5182 4903 4902 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09120 4903 4902 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09121 429 2774 4902 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09122 427 2774 4903 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09123 5182 4905 4904 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09124 4905 4904 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09125 430 2775 4904 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09126 428 2775 4905 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09127 5182 4907 4906 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09128 4907 4906 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09129 429 2775 4906 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09130 427 2775 4907 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09131 5182 4909 4908 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09132 4909 4908 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09133 430 2773 4908 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09134 428 2773 4909 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09135 5182 4911 4910 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09136 4911 4910 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09137 429 2773 4910 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09138 427 2773 4911 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09139 5182 4913 4912 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09140 4913 4912 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09141 430 2792 4912 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09142 428 2792 4913 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09143 5182 4915 4914 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09144 4915 4914 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09145 429 2792 4914 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09146 427 2792 4915 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09147 5182 4917 4916 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09148 4917 4916 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09149 430 2790 4916 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09150 428 2790 4917 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09151 5182 4919 4918 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09152 4919 4918 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09153 429 2790 4918 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09154 427 2790 4919 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09155 5182 4921 4920 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09156 4921 4920 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09157 430 2791 4920 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09158 428 2791 4921 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09159 5182 4923 4922 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09160 4923 4922 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09161 429 2791 4922 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09162 427 2791 4923 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09163 5182 4925 4924 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09164 4925 4924 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09165 430 2789 4924 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09166 428 2789 4925 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09167 5182 4927 4926 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09168 4927 4926 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09169 429 2789 4926 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09170 427 2789 4927 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09171 5182 4929 4928 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09172 4929 4928 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09173 430 2808 4928 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09174 428 2808 4929 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09175 5182 4931 4930 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09176 4931 4930 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09177 429 2808 4930 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09178 427 2808 4931 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09179 5182 4933 4932 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09180 4933 4932 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09181 430 2806 4932 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09182 428 2806 4933 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09183 5182 4935 4934 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09184 4935 4934 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09185 429 2806 4934 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09186 427 2806 4935 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09187 5182 4937 4936 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09188 4937 4936 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09189 430 2807 4936 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09190 428 2807 4937 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09191 5182 4939 4938 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09192 4939 4938 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09193 429 2807 4938 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09194 427 2807 4939 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09195 5182 4941 4940 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09196 4941 4940 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09197 430 2805 4940 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09198 428 2805 4941 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09199 5182 4943 4942 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09200 4943 4942 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09201 429 2805 4942 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09202 427 2805 4943 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09203 5182 4945 4944 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09204 4945 4944 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09205 430 2824 4944 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09206 428 2824 4945 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09207 5182 4947 4946 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09208 4947 4946 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09209 429 2824 4946 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09210 427 2824 4947 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09211 5182 4949 4948 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09212 4949 4948 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09213 430 2822 4948 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09214 428 2822 4949 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09215 5182 4951 4950 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09216 4951 4950 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09217 429 2822 4950 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09218 427 2822 4951 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09219 5182 4953 4952 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09220 4953 4952 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09221 430 2823 4952 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09222 428 2823 4953 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09223 5182 4955 4954 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09224 4955 4954 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09225 429 2823 4954 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09226 427 2823 4955 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09227 5182 4957 4956 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09228 4957 4956 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09229 430 2821 4956 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09230 428 2821 4957 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09231 5182 4959 4958 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09232 4959 4958 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09233 429 2821 4958 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09234 427 2821 4959 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09235 5182 4961 4960 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09236 4961 4960 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09237 430 2840 4960 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09238 428 2840 4961 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09239 5182 4963 4962 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09240 4963 4962 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09241 429 2840 4962 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09242 427 2840 4963 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09243 5182 4965 4964 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09244 4965 4964 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09245 430 2838 4964 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09246 428 2838 4965 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09247 5182 4967 4966 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09248 4967 4966 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09249 429 2838 4966 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09250 427 2838 4967 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09251 5182 4969 4968 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09252 4969 4968 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09253 430 2839 4968 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09254 428 2839 4969 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09255 5182 4971 4970 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09256 4971 4970 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09257 429 2839 4970 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09258 427 2839 4971 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09259 5182 4973 4972 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09260 4973 4972 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09261 430 2837 4972 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09262 428 2837 4973 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09263 5182 4975 4974 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09264 4975 4974 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09265 429 2837 4974 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09266 427 2837 4975 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09267 5182 4977 4976 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09268 4977 4976 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09269 430 2856 4976 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09270 428 2856 4977 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09271 5182 4979 4978 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09272 4979 4978 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09273 429 2856 4978 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09274 427 2856 4979 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09275 5182 4981 4980 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09276 4981 4980 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09277 430 2854 4980 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09278 428 2854 4981 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09279 5182 4983 4982 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09280 4983 4982 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09281 429 2854 4982 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09282 427 2854 4983 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09283 5182 4985 4984 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09284 4985 4984 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09285 430 2855 4984 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09286 428 2855 4985 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09287 5182 4987 4986 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09288 4987 4986 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09289 429 2855 4986 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09290 427 2855 4987 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09291 5182 4989 4988 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09292 4989 4988 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09293 430 2853 4988 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09294 428 2853 4989 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09295 5182 4991 4990 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09296 4991 4990 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09297 429 2853 4990 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09298 427 2853 4991 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09299 5182 4993 4992 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09300 4993 4992 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09301 430 2872 4992 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09302 428 2872 4993 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09303 5182 4995 4994 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09304 4995 4994 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09305 429 2872 4994 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09306 427 2872 4995 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09307 5182 4997 4996 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09308 4997 4996 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09309 430 2870 4996 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09310 428 2870 4997 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09311 5182 4999 4998 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09312 4999 4998 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09313 429 2870 4998 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09314 427 2870 4999 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09315 5182 5001 5000 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09316 5001 5000 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09317 430 2871 5000 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09318 428 2871 5001 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09319 5182 5003 5002 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09320 5003 5002 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09321 429 2871 5002 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09322 427 2871 5003 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09323 5182 5005 5004 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09324 5005 5004 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09325 430 2869 5004 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09326 428 2869 5005 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09327 5182 5007 5006 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09328 5007 5006 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09329 429 2869 5006 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09330 427 2869 5007 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09331 5182 5009 5008 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09332 5009 5008 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09333 430 2888 5008 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09334 428 2888 5009 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09335 5182 5011 5010 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09336 5011 5010 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09337 429 2888 5010 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09338 427 2888 5011 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09339 5182 5013 5012 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09340 5013 5012 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09341 430 2886 5012 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09342 428 2886 5013 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09343 5182 5015 5014 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09344 5015 5014 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09345 429 2886 5014 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09346 427 2886 5015 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09347 5182 5017 5016 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09348 5017 5016 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09349 430 2887 5016 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09350 428 2887 5017 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09351 5182 5019 5018 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09352 5019 5018 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09353 429 2887 5018 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09354 427 2887 5019 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09355 5182 5021 5020 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09356 5021 5020 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09357 430 2885 5020 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09358 428 2885 5021 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09359 5182 5023 5022 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09360 5023 5022 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09361 429 2885 5022 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09362 427 2885 5023 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09363 5182 5025 5024 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09364 5025 5024 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09365 430 2904 5024 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09366 428 2904 5025 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09367 5182 5027 5026 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09368 5027 5026 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09369 429 2904 5026 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09370 427 2904 5027 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09371 5182 5029 5028 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09372 5029 5028 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09373 430 2902 5028 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09374 428 2902 5029 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09375 5182 5031 5030 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09376 5031 5030 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09377 429 2902 5030 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09378 427 2902 5031 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09379 5182 5033 5032 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09380 5033 5032 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09381 430 2903 5032 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09382 428 2903 5033 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09383 5182 5035 5034 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09384 5035 5034 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09385 429 2903 5034 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09386 427 2903 5035 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09387 5182 5037 5036 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09388 5037 5036 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09389 430 2901 5036 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09390 428 2901 5037 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09391 5182 5039 5038 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09392 5039 5038 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09393 429 2901 5038 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09394 427 2901 5039 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09395 5182 5041 5040 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09396 5041 5040 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09397 430 2920 5040 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09398 428 2920 5041 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09399 5182 5043 5042 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09400 5043 5042 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09401 429 2920 5042 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09402 427 2920 5043 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09403 5182 5045 5044 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09404 5045 5044 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09405 430 2918 5044 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09406 428 2918 5045 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09407 5182 5047 5046 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09408 5047 5046 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09409 429 2918 5046 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09410 427 2918 5047 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09411 5182 5049 5048 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09412 5049 5048 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09413 430 2919 5048 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09414 428 2919 5049 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09415 5182 5051 5050 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09416 5051 5050 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09417 429 2919 5050 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09418 427 2919 5051 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09419 5182 5053 5052 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09420 5053 5052 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09421 430 2917 5052 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09422 428 2917 5053 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09423 5182 5055 5054 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09424 5055 5054 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09425 429 2917 5054 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09426 427 2917 5055 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09427 5182 5057 5056 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09428 5057 5056 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09429 430 2936 5056 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09430 428 2936 5057 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09431 5182 5059 5058 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09432 5059 5058 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09433 429 2936 5058 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09434 427 2936 5059 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09435 5182 5061 5060 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09436 5061 5060 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09437 430 2934 5060 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09438 428 2934 5061 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09439 5182 5063 5062 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09440 5063 5062 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09441 429 2934 5062 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09442 427 2934 5063 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09443 5182 5065 5064 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09444 5065 5064 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09445 430 2935 5064 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09446 428 2935 5065 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09447 5182 5067 5066 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09448 5067 5066 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09449 429 2935 5066 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09450 427 2935 5067 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09451 5182 5069 5068 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09452 5069 5068 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09453 430 2933 5068 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09454 428 2933 5069 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09455 5182 5071 5070 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09456 5071 5070 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09457 429 2933 5070 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09458 427 2933 5071 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09459 5182 5073 5072 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09460 5073 5072 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09461 430 2952 5072 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09462 428 2952 5073 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09463 5182 5075 5074 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09464 5075 5074 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09465 429 2952 5074 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09466 427 2952 5075 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09467 5182 5077 5076 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09468 5077 5076 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09469 430 2950 5076 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09470 428 2950 5077 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09471 5182 5079 5078 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09472 5079 5078 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09473 429 2950 5078 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09474 427 2950 5079 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09475 5182 5081 5080 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09476 5081 5080 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09477 430 2951 5080 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09478 428 2951 5081 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09479 5182 5083 5082 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09480 5083 5082 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09481 429 2951 5082 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09482 427 2951 5083 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09483 5182 5085 5084 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09484 5085 5084 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09485 430 2949 5084 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09486 428 2949 5085 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09487 5182 5087 5086 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09488 5087 5086 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09489 429 2949 5086 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09490 427 2949 5087 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09491 5182 5089 5088 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09492 5089 5088 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09493 430 2968 5088 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09494 428 2968 5089 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09495 5182 5091 5090 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09496 5091 5090 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09497 429 2968 5090 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09498 427 2968 5091 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09499 5182 5093 5092 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09500 5093 5092 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09501 430 2966 5092 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09502 428 2966 5093 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09503 5182 5095 5094 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09504 5095 5094 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09505 429 2966 5094 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09506 427 2966 5095 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09507 5182 5097 5096 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09508 5097 5096 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09509 430 2967 5096 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09510 428 2967 5097 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09511 5182 5099 5098 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09512 5099 5098 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09513 429 2967 5098 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09514 427 2967 5099 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09515 5182 5101 5100 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09516 5101 5100 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09517 430 2965 5100 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09518 428 2965 5101 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09519 5182 5103 5102 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09520 5103 5102 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09521 429 2965 5102 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09522 427 2965 5103 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09523 5182 5105 5104 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09524 5105 5104 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09525 430 2984 5104 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09526 428 2984 5105 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09527 5182 5107 5106 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09528 5107 5106 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09529 429 2984 5106 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09530 427 2984 5107 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09531 5182 5109 5108 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09532 5109 5108 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09533 430 2982 5108 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09534 428 2982 5109 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09535 5182 5111 5110 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09536 5111 5110 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09537 429 2982 5110 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09538 427 2982 5111 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09539 5182 5113 5112 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09540 5113 5112 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09541 430 2983 5112 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09542 428 2983 5113 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09543 5182 5115 5114 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09544 5115 5114 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09545 429 2983 5114 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09546 427 2983 5115 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09547 5182 5117 5116 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09548 5117 5116 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09549 430 2981 5116 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09550 428 2981 5117 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09551 5182 5119 5118 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09552 5119 5118 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09553 429 2981 5118 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09554 427 2981 5119 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09555 5182 5121 5120 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09556 5121 5120 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09557 430 3000 5120 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09558 428 3000 5121 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09559 5182 5123 5122 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09560 5123 5122 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09561 429 3000 5122 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09562 427 3000 5123 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09563 5182 5125 5124 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09564 5125 5124 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09565 430 2998 5124 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09566 428 2998 5125 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09567 5182 5127 5126 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09568 5127 5126 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09569 429 2998 5126 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09570 427 2998 5127 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09571 5182 5129 5128 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09572 5129 5128 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09573 430 2999 5128 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09574 428 2999 5129 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09575 5182 5131 5130 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09576 5131 5130 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09577 429 2999 5130 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09578 427 2999 5131 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09579 5182 5133 5132 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09580 5133 5132 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09581 430 2997 5132 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09582 428 2997 5133 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09583 5182 5135 5134 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09584 5135 5134 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09585 429 2997 5134 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09586 427 2997 5135 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09587 5182 5137 5136 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09588 5137 5136 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09589 430 3016 5136 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09590 428 3016 5137 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09591 5182 5139 5138 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09592 5139 5138 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09593 429 3016 5138 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09594 427 3016 5139 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09595 5182 5141 5140 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09596 5141 5140 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09597 430 3014 5140 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09598 428 3014 5141 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09599 5182 5143 5142 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09600 5143 5142 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09601 429 3014 5142 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09602 427 3014 5143 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09603 5182 5145 5144 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09604 5145 5144 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09605 430 3015 5144 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09606 428 3015 5145 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09607 5182 5147 5146 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09608 5147 5146 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09609 429 3015 5146 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09610 427 3015 5147 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09611 5182 5149 5148 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09612 5149 5148 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09613 430 3013 5148 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09614 428 3013 5149 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09615 5182 5151 5150 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09616 5151 5150 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09617 429 3013 5150 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09618 427 3013 5151 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09619 5182 5153 5152 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09620 5153 5152 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09621 430 3032 5152 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09622 428 3032 5153 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09623 5182 5155 5154 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09624 5155 5154 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09625 429 3032 5154 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09626 427 3032 5155 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09627 5182 5157 5156 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09628 5157 5156 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09629 430 3030 5156 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09630 428 3030 5157 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09631 5182 5159 5158 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09632 5159 5158 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09633 429 3030 5158 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09634 427 3030 5159 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09635 5182 5161 5160 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09636 5161 5160 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09637 430 3031 5160 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09638 428 3031 5161 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09639 5182 5163 5162 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09640 5163 5162 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09641 429 3031 5162 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09642 427 3031 5163 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09643 5182 5165 5164 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09644 5165 5164 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09645 430 3029 5164 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09646 428 3029 5165 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09647 5182 5167 5166 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09648 5167 5166 5182 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09649 429 3029 5166 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09650 427 3029 5167 5182 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09651 427 3045 434 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_09652 434 3046 428 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_09653 429 3045 435 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_09654 435 3046 430 5182 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_09655 5171 3081 5169 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_09656 5177 5171 431 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_09657 431 5176 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_09658 431 5169 5168 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_09659 5182 5176 432 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_09660 5170 435 432 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_09661 432 434 5169 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_09662 5171 435 433 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_09663 433 5176 5182 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_09664 433 434 5172 5182 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_09665 5183 3081 435 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_09666 435 3081 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_09667 5183 3081 434 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_09668 434 3081 5183 5182 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_09669 5173 5179 435 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_09670 434 5179 5174 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_09671 435 3081 434 5182 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_09672 5182 5185 5173 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_09673 5174 5175 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_09674 5173 5185 5182 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_09675 5182 5175 5174 5182 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_09676 5182 5185 5175 5182 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_09677 5185 5178 5182 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_09678 5182 5178 5185 5182 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_09679 5182 5179 5178 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_09680 5178 5177 5182 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_09681 5178 5176 5180 5182 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_09682 437 436 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09683 5183 437 436 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09684 439 438 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09685 5183 439 438 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09686 441 440 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09687 5183 441 440 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09688 443 442 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09689 5183 443 442 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09690 445 444 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09691 5183 445 444 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09692 447 446 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09693 5183 447 446 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09694 449 448 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09695 5183 449 448 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09696 451 450 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09697 5183 451 450 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09698 453 452 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09699 5183 453 452 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09700 455 454 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09701 5183 455 454 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09702 457 456 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09703 5183 457 456 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09704 459 458 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09705 5183 459 458 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09706 461 460 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09707 5183 461 460 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09708 463 462 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09709 5183 463 462 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09710 465 464 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09711 5183 465 464 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09712 467 466 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09713 5183 467 466 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09714 469 468 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09715 5183 469 468 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09716 471 470 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09717 5183 471 470 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09718 473 472 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09719 5183 473 472 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09720 475 474 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09721 5183 475 474 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09722 477 476 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09723 5183 477 476 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09724 479 478 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09725 5183 479 478 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09726 481 480 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09727 5183 481 480 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09728 483 482 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09729 5183 483 482 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09730 485 484 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09731 5183 485 484 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09732 487 486 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09733 5183 487 486 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09734 489 488 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09735 5183 489 488 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09736 491 490 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09737 5183 491 490 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09738 493 492 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09739 5183 493 492 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09740 495 494 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09741 5183 495 494 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09742 497 496 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09743 5183 497 496 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09744 499 498 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09745 5183 499 498 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09746 501 500 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09747 5183 501 500 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09748 503 502 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09749 5183 503 502 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09750 505 504 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09751 5183 505 504 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09752 507 506 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09753 5183 507 506 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09754 509 508 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09755 5183 509 508 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09756 511 510 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09757 5183 511 510 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09758 513 512 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09759 5183 513 512 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09760 515 514 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09761 5183 515 514 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09762 517 516 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09763 5183 517 516 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09764 519 518 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09765 5183 519 518 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09766 521 520 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09767 5183 521 520 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09768 523 522 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09769 5183 523 522 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09770 525 524 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09771 5183 525 524 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09772 527 526 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09773 5183 527 526 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09774 529 528 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09775 5183 529 528 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09776 531 530 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09777 5183 531 530 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09778 533 532 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09779 5183 533 532 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09780 535 534 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09781 5183 535 534 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09782 537 536 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09783 5183 537 536 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09784 539 538 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09785 5183 539 538 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09786 541 540 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09787 5183 541 540 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09788 543 542 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09789 5183 543 542 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09790 545 544 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09791 5183 545 544 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09792 547 546 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09793 5183 547 546 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09794 549 548 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09795 5183 549 548 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09796 551 550 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09797 5183 551 550 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09798 553 552 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09799 5183 553 552 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09800 555 554 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09801 5183 555 554 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09802 557 556 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09803 5183 557 556 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09804 559 558 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09805 5183 559 558 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09806 561 560 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09807 5183 561 560 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09808 563 562 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09809 5183 563 562 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09810 565 564 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09811 5183 565 564 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09812 567 566 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09813 5183 567 566 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09814 569 568 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09815 5183 569 568 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09816 571 570 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09817 5183 571 570 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09818 573 572 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09819 5183 573 572 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09820 575 574 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09821 5183 575 574 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09822 577 576 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09823 5183 577 576 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09824 579 578 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09825 5183 579 578 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09826 581 580 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09827 5183 581 580 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09828 583 582 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09829 5183 583 582 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09830 585 584 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09831 5183 585 584 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09832 587 586 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09833 5183 587 586 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09834 589 588 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09835 5183 589 588 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09836 591 590 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09837 5183 591 590 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09838 593 592 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09839 5183 593 592 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09840 595 594 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09841 5183 595 594 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09842 597 596 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09843 5183 597 596 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09844 599 598 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09845 5183 599 598 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09846 601 600 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09847 5183 601 600 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09848 603 602 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09849 5183 603 602 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09850 605 604 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09851 5183 605 604 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09852 607 606 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09853 5183 607 606 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09854 609 608 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09855 5183 609 608 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09856 611 610 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09857 5183 611 610 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09858 613 612 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09859 5183 613 612 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09860 615 614 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09861 5183 615 614 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09862 617 616 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09863 5183 617 616 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09864 619 618 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09865 5183 619 618 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09866 621 620 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09867 5183 621 620 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09868 623 622 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09869 5183 623 622 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09870 625 624 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09871 5183 625 624 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09872 627 626 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09873 5183 627 626 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09874 629 628 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09875 5183 629 628 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09876 631 630 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09877 5183 631 630 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09878 633 632 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09879 5183 633 632 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09880 635 634 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09881 5183 635 634 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09882 637 636 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09883 5183 637 636 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09884 639 638 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09885 5183 639 638 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09886 641 640 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09887 5183 641 640 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09888 643 642 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09889 5183 643 642 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09890 645 644 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09891 5183 645 644 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09892 647 646 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09893 5183 647 646 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09894 649 648 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09895 5183 649 648 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09896 651 650 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09897 5183 651 650 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09898 653 652 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09899 5183 653 652 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09900 655 654 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09901 5183 655 654 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09902 657 656 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09903 5183 657 656 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09904 659 658 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09905 5183 659 658 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09906 661 660 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09907 5183 661 660 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09908 663 662 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09909 5183 663 662 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09910 665 664 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09911 5183 665 664 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09912 667 666 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09913 5183 667 666 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09914 669 668 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09915 5183 669 668 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09916 671 670 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09917 5183 671 670 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09918 673 672 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09919 5183 673 672 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09920 675 674 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09921 5183 675 674 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09922 677 676 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09923 5183 677 676 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09924 679 678 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09925 5183 679 678 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09926 681 680 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09927 5183 681 680 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09928 683 682 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09929 5183 683 682 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09930 685 684 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09931 5183 685 684 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09932 687 686 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09933 5183 687 686 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09934 689 688 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09935 5183 689 688 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09936 691 690 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09937 5183 691 690 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09938 693 692 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09939 5183 693 692 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09940 695 694 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09941 5183 695 694 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09942 697 696 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09943 5183 697 696 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09944 699 698 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09945 5183 699 698 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09946 701 700 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09947 5183 701 700 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09948 703 702 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09949 5183 703 702 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09950 705 704 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09951 5183 705 704 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09952 707 706 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09953 5183 707 706 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09954 709 708 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09955 5183 709 708 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09956 711 710 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09957 5183 711 710 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09958 713 712 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09959 5183 713 712 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09960 715 714 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09961 5183 715 714 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09962 717 716 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09963 5183 717 716 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09964 719 718 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09965 5183 719 718 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09966 721 720 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09967 5183 721 720 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09968 723 722 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09969 5183 723 722 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09970 725 724 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09971 5183 725 724 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09972 727 726 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09973 5183 727 726 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09974 729 728 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09975 5183 729 728 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09976 731 730 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09977 5183 731 730 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09978 733 732 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09979 5183 733 732 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09980 735 734 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09981 5183 735 734 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09982 737 736 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09983 5183 737 736 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09984 739 738 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09985 5183 739 738 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09986 741 740 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09987 5183 741 740 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09988 743 742 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09989 5183 743 742 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09990 745 744 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09991 5183 745 744 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09992 747 746 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09993 5183 747 746 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09994 749 748 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09995 5183 749 748 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09996 751 750 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09997 5183 751 750 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09998 753 752 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_09999 5183 753 752 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10000 755 754 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10001 5183 755 754 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10002 757 756 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10003 5183 757 756 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10004 759 758 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10005 5183 759 758 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10006 761 760 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10007 5183 761 760 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10008 763 762 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10009 5183 763 762 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10010 765 764 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10011 5183 765 764 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10012 767 766 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10013 5183 767 766 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10014 769 768 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10015 5183 769 768 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10016 771 770 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10017 5183 771 770 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10018 773 772 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10019 5183 773 772 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10020 775 774 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10021 5183 775 774 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10022 777 776 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10023 5183 777 776 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10024 779 778 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10025 5183 779 778 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10026 781 780 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10027 5183 781 780 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10028 783 782 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10029 5183 783 782 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10030 785 784 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10031 5183 785 784 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10032 787 786 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10033 5183 787 786 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10034 789 788 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10035 5183 789 788 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10036 791 790 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10037 5183 791 790 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10038 793 792 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10039 5183 793 792 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10040 795 794 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10041 5183 795 794 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10042 797 796 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10043 5183 797 796 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10044 799 798 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10045 5183 799 798 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10046 801 800 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10047 5183 801 800 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10048 803 802 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10049 5183 803 802 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10050 805 804 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10051 5183 805 804 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10052 807 806 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10053 5183 807 806 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10054 809 808 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10055 5183 809 808 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10056 811 810 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10057 5183 811 810 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10058 813 812 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10059 5183 813 812 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10060 815 814 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10061 5183 815 814 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10062 817 816 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10063 5183 817 816 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10064 819 818 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10065 5183 819 818 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10066 821 820 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10067 5183 821 820 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10068 823 822 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10069 5183 823 822 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10070 825 824 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10071 5183 825 824 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10072 827 826 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10073 5183 827 826 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10074 829 828 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10075 5183 829 828 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10076 831 830 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10077 5183 831 830 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10078 833 832 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10079 5183 833 832 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10080 835 834 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10081 5183 835 834 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10082 837 836 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10083 5183 837 836 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10084 839 838 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10085 5183 839 838 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10086 841 840 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10087 5183 841 840 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10088 843 842 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10089 5183 843 842 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10090 845 844 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10091 5183 845 844 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10092 847 846 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10093 5183 847 846 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10094 849 848 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10095 5183 849 848 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10096 851 850 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10097 5183 851 850 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10098 853 852 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10099 5183 853 852 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10100 855 854 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10101 5183 855 854 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10102 857 856 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10103 5183 857 856 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10104 859 858 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10105 5183 859 858 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10106 861 860 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10107 5183 861 860 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10108 863 862 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10109 5183 863 862 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10110 865 864 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10111 5183 865 864 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10112 867 866 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10113 5183 867 866 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10114 869 868 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10115 5183 869 868 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10116 871 870 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10117 5183 871 870 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10118 873 872 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10119 5183 873 872 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10120 875 874 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10121 5183 875 874 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10122 877 876 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10123 5183 877 876 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10124 879 878 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10125 5183 879 878 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10126 881 880 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10127 5183 881 880 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10128 883 882 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10129 5183 883 882 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10130 885 884 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10131 5183 885 884 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10132 887 886 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10133 5183 887 886 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10134 889 888 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10135 5183 889 888 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10136 891 890 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10137 5183 891 890 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10138 893 892 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10139 5183 893 892 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10140 895 894 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10141 5183 895 894 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10142 897 896 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10143 5183 897 896 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10144 899 898 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10145 5183 899 898 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10146 901 900 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10147 5183 901 900 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10148 903 902 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10149 5183 903 902 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10150 905 904 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10151 5183 905 904 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10152 907 906 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10153 5183 907 906 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10154 909 908 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10155 5183 909 908 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10156 911 910 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10157 5183 911 910 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10158 913 912 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10159 5183 913 912 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10160 915 914 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10161 5183 915 914 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10162 917 916 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10163 5183 917 916 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10164 919 918 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10165 5183 919 918 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10166 921 920 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10167 5183 921 920 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10168 923 922 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10169 5183 923 922 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10170 925 924 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10171 5183 925 924 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10172 927 926 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10173 5183 927 926 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10174 929 928 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10175 5183 929 928 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10176 931 930 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10177 5183 931 930 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10178 933 932 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10179 5183 933 932 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10180 935 934 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10181 5183 935 934 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10182 937 936 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10183 5183 937 936 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10184 939 938 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10185 5183 939 938 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10186 941 940 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10187 5183 941 940 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10188 943 942 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10189 5183 943 942 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10190 945 944 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10191 5183 945 944 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10192 947 946 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10193 5183 947 946 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10194 956 948 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10195 5183 948 948 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10196 950 950 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10197 5183 950 949 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10198 951 952 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10199 5183 952 952 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10200 953 5192 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10201 5183 955 954 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10202 955 5192 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10203 5183 5192 955 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10204 5192 958 5183 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_10205 5183 958 5192 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_10206 5183 3074 958 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_10207 958 956 5183 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_10208 958 3077 957 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_10209 960 959 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10210 5183 960 959 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10211 962 961 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10212 5183 962 961 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10213 964 963 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10214 5183 964 963 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10215 966 965 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10216 5183 966 965 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10217 968 967 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10218 5183 968 967 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10219 970 969 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10220 5183 970 969 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10221 972 971 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10222 5183 972 971 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10223 974 973 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10224 5183 974 973 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10225 976 975 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10226 5183 976 975 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10227 978 977 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10228 5183 978 977 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10229 980 979 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10230 5183 980 979 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10231 982 981 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10232 5183 982 981 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10233 984 983 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10234 5183 984 983 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10235 986 985 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10236 5183 986 985 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10237 988 987 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10238 5183 988 987 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10239 990 989 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10240 5183 990 989 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10241 992 991 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10242 5183 992 991 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10243 994 993 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10244 5183 994 993 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10245 996 995 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10246 5183 996 995 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10247 998 997 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10248 5183 998 997 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10249 1000 999 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10250 5183 1000 999 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10251 1002 1001 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10252 5183 1002 1001 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10253 1004 1003 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10254 5183 1004 1003 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10255 1006 1005 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10256 5183 1006 1005 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10257 1008 1007 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10258 5183 1008 1007 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10259 1010 1009 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10260 5183 1010 1009 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10261 1012 1011 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10262 5183 1012 1011 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10263 1014 1013 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10264 5183 1014 1013 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10265 1016 1015 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10266 5183 1016 1015 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10267 1018 1017 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10268 5183 1018 1017 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10269 1020 1019 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10270 5183 1020 1019 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10271 1022 1021 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10272 5183 1022 1021 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10273 1024 1023 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10274 5183 1024 1023 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10275 1026 1025 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10276 5183 1026 1025 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10277 1028 1027 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10278 5183 1028 1027 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10279 1030 1029 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10280 5183 1030 1029 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10281 1032 1031 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10282 5183 1032 1031 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10283 1034 1033 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10284 5183 1034 1033 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10285 1036 1035 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10286 5183 1036 1035 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10287 1038 1037 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10288 5183 1038 1037 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10289 1040 1039 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10290 5183 1040 1039 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10291 1042 1041 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10292 5183 1042 1041 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10293 1044 1043 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10294 5183 1044 1043 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10295 1046 1045 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10296 5183 1046 1045 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10297 1048 1047 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10298 5183 1048 1047 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10299 1050 1049 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10300 5183 1050 1049 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10301 1052 1051 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10302 5183 1052 1051 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10303 1054 1053 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10304 5183 1054 1053 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10305 1056 1055 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10306 5183 1056 1055 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10307 1058 1057 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10308 5183 1058 1057 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10309 1060 1059 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10310 5183 1060 1059 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10311 1062 1061 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10312 5183 1062 1061 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10313 1064 1063 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10314 5183 1064 1063 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10315 1066 1065 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10316 5183 1066 1065 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10317 1068 1067 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10318 5183 1068 1067 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10319 1070 1069 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10320 5183 1070 1069 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10321 1072 1071 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10322 5183 1072 1071 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10323 1074 1073 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10324 5183 1074 1073 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10325 1076 1075 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10326 5183 1076 1075 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10327 1078 1077 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10328 5183 1078 1077 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10329 1080 1079 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10330 5183 1080 1079 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10331 1082 1081 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10332 5183 1082 1081 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10333 1084 1083 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10334 5183 1084 1083 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10335 1086 1085 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10336 5183 1086 1085 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10337 1088 1087 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10338 5183 1088 1087 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10339 1090 1089 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10340 5183 1090 1089 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10341 1092 1091 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10342 5183 1092 1091 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10343 1094 1093 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10344 5183 1094 1093 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10345 1096 1095 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10346 5183 1096 1095 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10347 1098 1097 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10348 5183 1098 1097 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10349 1100 1099 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10350 5183 1100 1099 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10351 1102 1101 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10352 5183 1102 1101 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10353 1104 1103 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10354 5183 1104 1103 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10355 1106 1105 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10356 5183 1106 1105 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10357 1108 1107 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10358 5183 1108 1107 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10359 1110 1109 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10360 5183 1110 1109 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10361 1112 1111 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10362 5183 1112 1111 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10363 1114 1113 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10364 5183 1114 1113 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10365 1116 1115 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10366 5183 1116 1115 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10367 1118 1117 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10368 5183 1118 1117 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10369 1120 1119 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10370 5183 1120 1119 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10371 1122 1121 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10372 5183 1122 1121 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10373 1124 1123 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10374 5183 1124 1123 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10375 1126 1125 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10376 5183 1126 1125 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10377 1128 1127 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10378 5183 1128 1127 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10379 1130 1129 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10380 5183 1130 1129 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10381 1132 1131 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10382 5183 1132 1131 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10383 1134 1133 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10384 5183 1134 1133 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10385 1136 1135 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10386 5183 1136 1135 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10387 1138 1137 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10388 5183 1138 1137 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10389 1140 1139 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10390 5183 1140 1139 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10391 1142 1141 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10392 5183 1142 1141 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10393 1144 1143 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10394 5183 1144 1143 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10395 1146 1145 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10396 5183 1146 1145 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10397 1148 1147 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10398 5183 1148 1147 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10399 1150 1149 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10400 5183 1150 1149 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10401 1152 1151 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10402 5183 1152 1151 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10403 1154 1153 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10404 5183 1154 1153 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10405 1156 1155 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10406 5183 1156 1155 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10407 1158 1157 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10408 5183 1158 1157 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10409 1160 1159 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10410 5183 1160 1159 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10411 1162 1161 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10412 5183 1162 1161 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10413 1164 1163 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10414 5183 1164 1163 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10415 1166 1165 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10416 5183 1166 1165 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10417 1168 1167 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10418 5183 1168 1167 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10419 1170 1169 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10420 5183 1170 1169 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10421 1172 1171 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10422 5183 1172 1171 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10423 1174 1173 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10424 5183 1174 1173 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10425 1176 1175 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10426 5183 1176 1175 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10427 1178 1177 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10428 5183 1178 1177 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10429 1180 1179 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10430 5183 1180 1179 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10431 1182 1181 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10432 5183 1182 1181 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10433 1184 1183 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10434 5183 1184 1183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10435 1186 1185 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10436 5183 1186 1185 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10437 1188 1187 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10438 5183 1188 1187 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10439 1190 1189 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10440 5183 1190 1189 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10441 1192 1191 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10442 5183 1192 1191 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10443 1194 1193 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10444 5183 1194 1193 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10445 1196 1195 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10446 5183 1196 1195 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10447 1198 1197 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10448 5183 1198 1197 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10449 1200 1199 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10450 5183 1200 1199 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10451 1202 1201 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10452 5183 1202 1201 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10453 1204 1203 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10454 5183 1204 1203 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10455 1206 1205 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10456 5183 1206 1205 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10457 1208 1207 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10458 5183 1208 1207 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10459 1210 1209 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10460 5183 1210 1209 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10461 1212 1211 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10462 5183 1212 1211 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10463 1214 1213 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10464 5183 1214 1213 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10465 1216 1215 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10466 5183 1216 1215 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10467 1218 1217 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10468 5183 1218 1217 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10469 1220 1219 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10470 5183 1220 1219 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10471 1222 1221 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10472 5183 1222 1221 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10473 1224 1223 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10474 5183 1224 1223 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10475 1226 1225 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10476 5183 1226 1225 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10477 1228 1227 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10478 5183 1228 1227 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10479 1230 1229 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10480 5183 1230 1229 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10481 1232 1231 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10482 5183 1232 1231 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10483 1234 1233 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10484 5183 1234 1233 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10485 1236 1235 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10486 5183 1236 1235 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10487 1238 1237 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10488 5183 1238 1237 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10489 1240 1239 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10490 5183 1240 1239 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10491 1242 1241 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10492 5183 1242 1241 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10493 1244 1243 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10494 5183 1244 1243 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10495 1246 1245 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10496 5183 1246 1245 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10497 1248 1247 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10498 5183 1248 1247 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10499 1250 1249 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10500 5183 1250 1249 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10501 1252 1251 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10502 5183 1252 1251 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10503 1254 1253 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10504 5183 1254 1253 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10505 1256 1255 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10506 5183 1256 1255 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10507 1258 1257 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10508 5183 1258 1257 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10509 1260 1259 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10510 5183 1260 1259 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10511 1262 1261 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10512 5183 1262 1261 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10513 1264 1263 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10514 5183 1264 1263 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10515 1266 1265 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10516 5183 1266 1265 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10517 1268 1267 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10518 5183 1268 1267 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10519 1270 1269 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10520 5183 1270 1269 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10521 1272 1271 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10522 5183 1272 1271 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10523 1274 1273 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10524 5183 1274 1273 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10525 1276 1275 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10526 5183 1276 1275 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10527 1278 1277 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10528 5183 1278 1277 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10529 1280 1279 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10530 5183 1280 1279 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10531 1282 1281 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10532 5183 1282 1281 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10533 1284 1283 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10534 5183 1284 1283 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10535 1286 1285 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10536 5183 1286 1285 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10537 1288 1287 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10538 5183 1288 1287 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10539 1290 1289 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10540 5183 1290 1289 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10541 1292 1291 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10542 5183 1292 1291 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10543 1294 1293 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10544 5183 1294 1293 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10545 1296 1295 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10546 5183 1296 1295 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10547 1298 1297 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10548 5183 1298 1297 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10549 1300 1299 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10550 5183 1300 1299 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10551 1302 1301 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10552 5183 1302 1301 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10553 1304 1303 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10554 5183 1304 1303 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10555 1306 1305 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10556 5183 1306 1305 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10557 1308 1307 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10558 5183 1308 1307 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10559 1310 1309 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10560 5183 1310 1309 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10561 1312 1311 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10562 5183 1312 1311 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10563 1314 1313 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10564 5183 1314 1313 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10565 1316 1315 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10566 5183 1316 1315 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10567 1318 1317 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10568 5183 1318 1317 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10569 1320 1319 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10570 5183 1320 1319 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10571 1322 1321 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10572 5183 1322 1321 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10573 1324 1323 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10574 5183 1324 1323 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10575 1326 1325 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10576 5183 1326 1325 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10577 1328 1327 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10578 5183 1328 1327 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10579 1330 1329 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10580 5183 1330 1329 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10581 1332 1331 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10582 5183 1332 1331 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10583 1334 1333 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10584 5183 1334 1333 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10585 1336 1335 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10586 5183 1336 1335 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10587 1338 1337 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10588 5183 1338 1337 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10589 1340 1339 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10590 5183 1340 1339 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10591 1342 1341 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10592 5183 1342 1341 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10593 1344 1343 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10594 5183 1344 1343 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10595 1346 1345 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10596 5183 1346 1345 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10597 1348 1347 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10598 5183 1348 1347 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10599 1350 1349 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10600 5183 1350 1349 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10601 1352 1351 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10602 5183 1352 1351 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10603 1354 1353 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10604 5183 1354 1353 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10605 1356 1355 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10606 5183 1356 1355 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10607 1358 1357 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10608 5183 1358 1357 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10609 1360 1359 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10610 5183 1360 1359 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10611 1362 1361 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10612 5183 1362 1361 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10613 1364 1363 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10614 5183 1364 1363 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10615 1366 1365 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10616 5183 1366 1365 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10617 1368 1367 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10618 5183 1368 1367 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10619 1370 1369 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10620 5183 1370 1369 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10621 1372 1371 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10622 5183 1372 1371 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10623 1374 1373 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10624 5183 1374 1373 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10625 1376 1375 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10626 5183 1376 1375 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10627 1378 1377 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10628 5183 1378 1377 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10629 1380 1379 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10630 5183 1380 1379 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10631 1382 1381 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10632 5183 1382 1381 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10633 1384 1383 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10634 5183 1384 1383 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10635 1386 1385 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10636 5183 1386 1385 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10637 1388 1387 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10638 5183 1388 1387 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10639 1390 1389 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10640 5183 1390 1389 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10641 1392 1391 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10642 5183 1392 1391 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10643 1394 1393 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10644 5183 1394 1393 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10645 1396 1395 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10646 5183 1396 1395 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10647 1398 1397 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10648 5183 1398 1397 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10649 1400 1399 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10650 5183 1400 1399 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10651 1402 1401 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10652 5183 1402 1401 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10653 1404 1403 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10654 5183 1404 1403 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10655 1406 1405 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10656 5183 1406 1405 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10657 1408 1407 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10658 5183 1408 1407 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10659 1410 1409 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10660 5183 1410 1409 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10661 1412 1411 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10662 5183 1412 1411 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10663 1414 1413 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10664 5183 1414 1413 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10665 1416 1415 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10666 5183 1416 1415 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10667 1418 1417 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10668 5183 1418 1417 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10669 1420 1419 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10670 5183 1420 1419 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10671 1422 1421 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10672 5183 1422 1421 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10673 1424 1423 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10674 5183 1424 1423 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10675 1426 1425 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10676 5183 1426 1425 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10677 1428 1427 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10678 5183 1428 1427 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10679 1430 1429 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10680 5183 1430 1429 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10681 1432 1431 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10682 5183 1432 1431 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10683 1434 1433 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10684 5183 1434 1433 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10685 1436 1435 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10686 5183 1436 1435 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10687 1438 1437 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10688 5183 1438 1437 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10689 1440 1439 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10690 5183 1440 1439 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10691 1442 1441 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10692 5183 1442 1441 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10693 1444 1443 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10694 5183 1444 1443 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10695 1446 1445 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10696 5183 1446 1445 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10697 1448 1447 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10698 5183 1448 1447 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10699 1450 1449 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10700 5183 1450 1449 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10701 1452 1451 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10702 5183 1452 1451 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10703 1454 1453 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10704 5183 1454 1453 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10705 1456 1455 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10706 5183 1456 1455 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10707 1458 1457 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10708 5183 1458 1457 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10709 1460 1459 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10710 5183 1460 1459 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10711 1462 1461 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10712 5183 1462 1461 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10713 1464 1463 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10714 5183 1464 1463 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10715 1466 1465 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10716 5183 1466 1465 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10717 1468 1467 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10718 5183 1468 1467 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10719 1470 1469 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10720 5183 1470 1469 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10721 1479 1471 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10722 5183 1471 1471 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10723 1473 1473 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10724 5183 1473 1472 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10725 1474 1475 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10726 5183 1475 1475 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10727 1476 5191 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10728 5183 1478 1477 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10729 1478 5191 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10730 5183 5191 1478 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_10731 5191 1481 5183 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_10732 5183 1481 5191 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_10733 5183 3074 1481 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_10734 1481 1479 5183 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_10735 1481 3077 1480 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_10736 1483 1482 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10737 5183 1483 1482 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10738 1485 1484 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10739 5183 1485 1484 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10740 1487 1486 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10741 5183 1487 1486 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10742 1489 1488 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10743 5183 1489 1488 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10744 1491 1490 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10745 5183 1491 1490 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10746 1493 1492 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10747 5183 1493 1492 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10748 1495 1494 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10749 5183 1495 1494 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10750 1497 1496 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10751 5183 1497 1496 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10752 1499 1498 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10753 5183 1499 1498 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10754 1501 1500 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10755 5183 1501 1500 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10756 1503 1502 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10757 5183 1503 1502 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10758 1505 1504 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10759 5183 1505 1504 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10760 1507 1506 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10761 5183 1507 1506 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10762 1509 1508 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10763 5183 1509 1508 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10764 1511 1510 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10765 5183 1511 1510 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10766 1513 1512 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10767 5183 1513 1512 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10768 1515 1514 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10769 5183 1515 1514 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10770 1517 1516 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10771 5183 1517 1516 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10772 1519 1518 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10773 5183 1519 1518 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10774 1521 1520 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10775 5183 1521 1520 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10776 1523 1522 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10777 5183 1523 1522 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10778 1525 1524 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10779 5183 1525 1524 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10780 1527 1526 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10781 5183 1527 1526 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10782 1529 1528 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10783 5183 1529 1528 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10784 1531 1530 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10785 5183 1531 1530 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10786 1533 1532 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10787 5183 1533 1532 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10788 1535 1534 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10789 5183 1535 1534 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10790 1537 1536 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10791 5183 1537 1536 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10792 1539 1538 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10793 5183 1539 1538 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10794 1541 1540 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10795 5183 1541 1540 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10796 1543 1542 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10797 5183 1543 1542 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10798 1545 1544 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10799 5183 1545 1544 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10800 1547 1546 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10801 5183 1547 1546 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10802 1549 1548 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10803 5183 1549 1548 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10804 1551 1550 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10805 5183 1551 1550 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10806 1553 1552 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10807 5183 1553 1552 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10808 1555 1554 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10809 5183 1555 1554 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10810 1557 1556 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10811 5183 1557 1556 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10812 1559 1558 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10813 5183 1559 1558 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10814 1561 1560 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10815 5183 1561 1560 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10816 1563 1562 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10817 5183 1563 1562 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10818 1565 1564 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10819 5183 1565 1564 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10820 1567 1566 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10821 5183 1567 1566 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10822 1569 1568 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10823 5183 1569 1568 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10824 1571 1570 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10825 5183 1571 1570 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10826 1573 1572 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10827 5183 1573 1572 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10828 1575 1574 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10829 5183 1575 1574 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10830 1577 1576 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10831 5183 1577 1576 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10832 1579 1578 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10833 5183 1579 1578 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10834 1581 1580 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10835 5183 1581 1580 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10836 1583 1582 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10837 5183 1583 1582 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10838 1585 1584 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10839 5183 1585 1584 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10840 1587 1586 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10841 5183 1587 1586 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10842 1589 1588 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10843 5183 1589 1588 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10844 1591 1590 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10845 5183 1591 1590 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10846 1593 1592 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10847 5183 1593 1592 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10848 1595 1594 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10849 5183 1595 1594 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10850 1597 1596 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10851 5183 1597 1596 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10852 1599 1598 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10853 5183 1599 1598 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10854 1601 1600 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10855 5183 1601 1600 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10856 1603 1602 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10857 5183 1603 1602 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10858 1605 1604 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10859 5183 1605 1604 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10860 1607 1606 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10861 5183 1607 1606 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10862 1609 1608 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10863 5183 1609 1608 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10864 1611 1610 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10865 5183 1611 1610 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10866 1613 1612 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10867 5183 1613 1612 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10868 1615 1614 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10869 5183 1615 1614 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10870 1617 1616 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10871 5183 1617 1616 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10872 1619 1618 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10873 5183 1619 1618 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10874 1621 1620 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10875 5183 1621 1620 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10876 1623 1622 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10877 5183 1623 1622 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10878 1625 1624 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10879 5183 1625 1624 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10880 1627 1626 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10881 5183 1627 1626 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10882 1629 1628 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10883 5183 1629 1628 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10884 1631 1630 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10885 5183 1631 1630 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10886 1633 1632 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10887 5183 1633 1632 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10888 1635 1634 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10889 5183 1635 1634 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10890 1637 1636 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10891 5183 1637 1636 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10892 1639 1638 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10893 5183 1639 1638 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10894 1641 1640 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10895 5183 1641 1640 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10896 1643 1642 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10897 5183 1643 1642 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10898 1645 1644 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10899 5183 1645 1644 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10900 1647 1646 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10901 5183 1647 1646 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10902 1649 1648 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10903 5183 1649 1648 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10904 1651 1650 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10905 5183 1651 1650 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10906 1653 1652 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10907 5183 1653 1652 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10908 1655 1654 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10909 5183 1655 1654 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10910 1657 1656 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10911 5183 1657 1656 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10912 1659 1658 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10913 5183 1659 1658 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10914 1661 1660 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10915 5183 1661 1660 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10916 1663 1662 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10917 5183 1663 1662 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10918 1665 1664 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10919 5183 1665 1664 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10920 1667 1666 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10921 5183 1667 1666 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10922 1669 1668 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10923 5183 1669 1668 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10924 1671 1670 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10925 5183 1671 1670 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10926 1673 1672 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10927 5183 1673 1672 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10928 1675 1674 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10929 5183 1675 1674 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10930 1677 1676 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10931 5183 1677 1676 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10932 1679 1678 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10933 5183 1679 1678 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10934 1681 1680 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10935 5183 1681 1680 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10936 1683 1682 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10937 5183 1683 1682 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10938 1685 1684 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10939 5183 1685 1684 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10940 1687 1686 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10941 5183 1687 1686 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10942 1689 1688 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10943 5183 1689 1688 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10944 1691 1690 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10945 5183 1691 1690 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10946 1693 1692 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10947 5183 1693 1692 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10948 1695 1694 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10949 5183 1695 1694 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10950 1697 1696 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10951 5183 1697 1696 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10952 1699 1698 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10953 5183 1699 1698 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10954 1701 1700 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10955 5183 1701 1700 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10956 1703 1702 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10957 5183 1703 1702 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10958 1705 1704 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10959 5183 1705 1704 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10960 1707 1706 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10961 5183 1707 1706 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10962 1709 1708 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10963 5183 1709 1708 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10964 1711 1710 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10965 5183 1711 1710 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10966 1713 1712 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10967 5183 1713 1712 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10968 1715 1714 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10969 5183 1715 1714 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10970 1717 1716 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10971 5183 1717 1716 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10972 1719 1718 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10973 5183 1719 1718 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10974 1721 1720 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10975 5183 1721 1720 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10976 1723 1722 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10977 5183 1723 1722 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10978 1725 1724 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10979 5183 1725 1724 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10980 1727 1726 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10981 5183 1727 1726 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10982 1729 1728 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10983 5183 1729 1728 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10984 1731 1730 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10985 5183 1731 1730 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10986 1733 1732 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10987 5183 1733 1732 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10988 1735 1734 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10989 5183 1735 1734 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10990 1737 1736 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10991 5183 1737 1736 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10992 1739 1738 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10993 5183 1739 1738 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10994 1741 1740 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10995 5183 1741 1740 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10996 1743 1742 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10997 5183 1743 1742 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10998 1745 1744 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_10999 5183 1745 1744 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11000 1747 1746 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11001 5183 1747 1746 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11002 1749 1748 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11003 5183 1749 1748 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11004 1751 1750 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11005 5183 1751 1750 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11006 1753 1752 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11007 5183 1753 1752 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11008 1755 1754 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11009 5183 1755 1754 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11010 1757 1756 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11011 5183 1757 1756 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11012 1759 1758 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11013 5183 1759 1758 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11014 1761 1760 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11015 5183 1761 1760 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11016 1763 1762 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11017 5183 1763 1762 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11018 1765 1764 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11019 5183 1765 1764 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11020 1767 1766 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11021 5183 1767 1766 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11022 1769 1768 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11023 5183 1769 1768 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11024 1771 1770 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11025 5183 1771 1770 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11026 1773 1772 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11027 5183 1773 1772 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11028 1775 1774 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11029 5183 1775 1774 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11030 1777 1776 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11031 5183 1777 1776 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11032 1779 1778 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11033 5183 1779 1778 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11034 1781 1780 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11035 5183 1781 1780 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11036 1783 1782 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11037 5183 1783 1782 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11038 1785 1784 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11039 5183 1785 1784 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11040 1787 1786 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11041 5183 1787 1786 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11042 1789 1788 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11043 5183 1789 1788 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11044 1791 1790 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11045 5183 1791 1790 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11046 1793 1792 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11047 5183 1793 1792 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11048 1795 1794 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11049 5183 1795 1794 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11050 1797 1796 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11051 5183 1797 1796 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11052 1799 1798 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11053 5183 1799 1798 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11054 1801 1800 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11055 5183 1801 1800 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11056 1803 1802 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11057 5183 1803 1802 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11058 1805 1804 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11059 5183 1805 1804 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11060 1807 1806 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11061 5183 1807 1806 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11062 1809 1808 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11063 5183 1809 1808 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11064 1811 1810 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11065 5183 1811 1810 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11066 1813 1812 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11067 5183 1813 1812 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11068 1815 1814 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11069 5183 1815 1814 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11070 1817 1816 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11071 5183 1817 1816 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11072 1819 1818 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11073 5183 1819 1818 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11074 1821 1820 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11075 5183 1821 1820 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11076 1823 1822 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11077 5183 1823 1822 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11078 1825 1824 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11079 5183 1825 1824 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11080 1827 1826 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11081 5183 1827 1826 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11082 1829 1828 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11083 5183 1829 1828 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11084 1831 1830 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11085 5183 1831 1830 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11086 1833 1832 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11087 5183 1833 1832 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11088 1835 1834 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11089 5183 1835 1834 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11090 1837 1836 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11091 5183 1837 1836 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11092 1839 1838 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11093 5183 1839 1838 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11094 1841 1840 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11095 5183 1841 1840 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11096 1843 1842 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11097 5183 1843 1842 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11098 1845 1844 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11099 5183 1845 1844 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11100 1847 1846 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11101 5183 1847 1846 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11102 1849 1848 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11103 5183 1849 1848 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11104 1851 1850 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11105 5183 1851 1850 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11106 1853 1852 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11107 5183 1853 1852 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11108 1855 1854 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11109 5183 1855 1854 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11110 1857 1856 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11111 5183 1857 1856 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11112 1859 1858 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11113 5183 1859 1858 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11114 1861 1860 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11115 5183 1861 1860 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11116 1863 1862 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11117 5183 1863 1862 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11118 1865 1864 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11119 5183 1865 1864 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11120 1867 1866 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11121 5183 1867 1866 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11122 1869 1868 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11123 5183 1869 1868 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11124 1871 1870 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11125 5183 1871 1870 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11126 1873 1872 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11127 5183 1873 1872 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11128 1875 1874 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11129 5183 1875 1874 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11130 1877 1876 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11131 5183 1877 1876 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11132 1879 1878 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11133 5183 1879 1878 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11134 1881 1880 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11135 5183 1881 1880 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11136 1883 1882 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11137 5183 1883 1882 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11138 1885 1884 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11139 5183 1885 1884 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11140 1887 1886 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11141 5183 1887 1886 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11142 1889 1888 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11143 5183 1889 1888 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11144 1891 1890 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11145 5183 1891 1890 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11146 1893 1892 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11147 5183 1893 1892 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11148 1895 1894 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11149 5183 1895 1894 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11150 1897 1896 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11151 5183 1897 1896 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11152 1899 1898 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11153 5183 1899 1898 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11154 1901 1900 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11155 5183 1901 1900 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11156 1903 1902 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11157 5183 1903 1902 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11158 1905 1904 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11159 5183 1905 1904 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11160 1907 1906 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11161 5183 1907 1906 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11162 1909 1908 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11163 5183 1909 1908 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11164 1911 1910 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11165 5183 1911 1910 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11166 1913 1912 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11167 5183 1913 1912 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11168 1915 1914 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11169 5183 1915 1914 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11170 1917 1916 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11171 5183 1917 1916 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11172 1919 1918 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11173 5183 1919 1918 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11174 1921 1920 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11175 5183 1921 1920 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11176 1923 1922 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11177 5183 1923 1922 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11178 1925 1924 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11179 5183 1925 1924 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11180 1927 1926 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11181 5183 1927 1926 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11182 1929 1928 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11183 5183 1929 1928 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11184 1931 1930 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11185 5183 1931 1930 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11186 1933 1932 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11187 5183 1933 1932 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11188 1935 1934 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11189 5183 1935 1934 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11190 1937 1936 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11191 5183 1937 1936 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11192 1939 1938 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11193 5183 1939 1938 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11194 1941 1940 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11195 5183 1941 1940 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11196 1943 1942 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11197 5183 1943 1942 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11198 1945 1944 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11199 5183 1945 1944 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11200 1947 1946 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11201 5183 1947 1946 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11202 1949 1948 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11203 5183 1949 1948 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11204 1951 1950 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11205 5183 1951 1950 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11206 1953 1952 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11207 5183 1953 1952 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11208 1955 1954 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11209 5183 1955 1954 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11210 1957 1956 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11211 5183 1957 1956 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11212 1959 1958 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11213 5183 1959 1958 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11214 1961 1960 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11215 5183 1961 1960 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11216 1963 1962 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11217 5183 1963 1962 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11218 1965 1964 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11219 5183 1965 1964 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11220 1967 1966 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11221 5183 1967 1966 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11222 1969 1968 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11223 5183 1969 1968 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11224 1971 1970 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11225 5183 1971 1970 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11226 1973 1972 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11227 5183 1973 1972 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11228 1975 1974 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11229 5183 1975 1974 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11230 1977 1976 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11231 5183 1977 1976 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11232 1979 1978 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11233 5183 1979 1978 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11234 1981 1980 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11235 5183 1981 1980 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11236 1983 1982 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11237 5183 1983 1982 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11238 1985 1984 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11239 5183 1985 1984 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11240 1987 1986 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11241 5183 1987 1986 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11242 1989 1988 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11243 5183 1989 1988 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11244 1991 1990 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11245 5183 1991 1990 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11246 1993 1992 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11247 5183 1993 1992 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11248 2002 1994 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11249 5183 1994 1994 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11250 1996 1996 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11251 5183 1996 1995 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11252 1997 1998 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11253 5183 1998 1998 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11254 1999 5190 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11255 5183 2001 2000 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11256 2001 5190 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11257 5183 5190 2001 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11258 5190 2004 5183 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_11259 5183 2004 5190 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_11260 5183 3074 2004 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_11261 2004 2002 5183 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_11262 2004 3077 2003 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_11263 2006 2005 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11264 5183 2006 2005 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11265 2008 2007 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11266 5183 2008 2007 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11267 2010 2009 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11268 5183 2010 2009 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11269 2012 2011 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11270 5183 2012 2011 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11271 2014 2013 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11272 5183 2014 2013 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11273 2016 2015 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11274 5183 2016 2015 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11275 2018 2017 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11276 5183 2018 2017 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11277 2020 2019 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11278 5183 2020 2019 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11279 2022 2021 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11280 5183 2022 2021 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11281 2024 2023 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11282 5183 2024 2023 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11283 2026 2025 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11284 5183 2026 2025 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11285 2028 2027 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11286 5183 2028 2027 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11287 2030 2029 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11288 5183 2030 2029 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11289 2032 2031 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11290 5183 2032 2031 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11291 2034 2033 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11292 5183 2034 2033 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11293 2036 2035 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11294 5183 2036 2035 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11295 2038 2037 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11296 5183 2038 2037 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11297 2040 2039 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11298 5183 2040 2039 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11299 2042 2041 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11300 5183 2042 2041 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11301 2044 2043 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11302 5183 2044 2043 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11303 2046 2045 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11304 5183 2046 2045 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11305 2048 2047 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11306 5183 2048 2047 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11307 2050 2049 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11308 5183 2050 2049 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11309 2052 2051 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11310 5183 2052 2051 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11311 2054 2053 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11312 5183 2054 2053 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11313 2056 2055 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11314 5183 2056 2055 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11315 2058 2057 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11316 5183 2058 2057 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11317 2060 2059 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11318 5183 2060 2059 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11319 2062 2061 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11320 5183 2062 2061 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11321 2064 2063 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11322 5183 2064 2063 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11323 2066 2065 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11324 5183 2066 2065 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11325 2068 2067 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11326 5183 2068 2067 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11327 2070 2069 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11328 5183 2070 2069 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11329 2072 2071 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11330 5183 2072 2071 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11331 2074 2073 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11332 5183 2074 2073 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11333 2076 2075 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11334 5183 2076 2075 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11335 2078 2077 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11336 5183 2078 2077 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11337 2080 2079 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11338 5183 2080 2079 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11339 2082 2081 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11340 5183 2082 2081 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11341 2084 2083 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11342 5183 2084 2083 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11343 2086 2085 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11344 5183 2086 2085 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11345 2088 2087 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11346 5183 2088 2087 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11347 2090 2089 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11348 5183 2090 2089 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11349 2092 2091 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11350 5183 2092 2091 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11351 2094 2093 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11352 5183 2094 2093 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11353 2096 2095 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11354 5183 2096 2095 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11355 2098 2097 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11356 5183 2098 2097 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11357 2100 2099 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11358 5183 2100 2099 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11359 2102 2101 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11360 5183 2102 2101 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11361 2104 2103 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11362 5183 2104 2103 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11363 2106 2105 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11364 5183 2106 2105 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11365 2108 2107 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11366 5183 2108 2107 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11367 2110 2109 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11368 5183 2110 2109 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11369 2112 2111 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11370 5183 2112 2111 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11371 2114 2113 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11372 5183 2114 2113 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11373 2116 2115 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11374 5183 2116 2115 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11375 2118 2117 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11376 5183 2118 2117 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11377 2120 2119 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11378 5183 2120 2119 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11379 2122 2121 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11380 5183 2122 2121 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11381 2124 2123 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11382 5183 2124 2123 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11383 2126 2125 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11384 5183 2126 2125 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11385 2128 2127 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11386 5183 2128 2127 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11387 2130 2129 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11388 5183 2130 2129 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11389 2132 2131 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11390 5183 2132 2131 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11391 2134 2133 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11392 5183 2134 2133 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11393 2136 2135 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11394 5183 2136 2135 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11395 2138 2137 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11396 5183 2138 2137 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11397 2140 2139 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11398 5183 2140 2139 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11399 2142 2141 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11400 5183 2142 2141 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11401 2144 2143 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11402 5183 2144 2143 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11403 2146 2145 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11404 5183 2146 2145 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11405 2148 2147 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11406 5183 2148 2147 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11407 2150 2149 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11408 5183 2150 2149 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11409 2152 2151 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11410 5183 2152 2151 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11411 2154 2153 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11412 5183 2154 2153 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11413 2156 2155 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11414 5183 2156 2155 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11415 2158 2157 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11416 5183 2158 2157 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11417 2160 2159 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11418 5183 2160 2159 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11419 2162 2161 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11420 5183 2162 2161 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11421 2164 2163 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11422 5183 2164 2163 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11423 2166 2165 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11424 5183 2166 2165 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11425 2168 2167 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11426 5183 2168 2167 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11427 2170 2169 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11428 5183 2170 2169 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11429 2172 2171 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11430 5183 2172 2171 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11431 2174 2173 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11432 5183 2174 2173 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11433 2176 2175 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11434 5183 2176 2175 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11435 2178 2177 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11436 5183 2178 2177 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11437 2180 2179 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11438 5183 2180 2179 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11439 2182 2181 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11440 5183 2182 2181 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11441 2184 2183 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11442 5183 2184 2183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11443 2186 2185 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11444 5183 2186 2185 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11445 2188 2187 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11446 5183 2188 2187 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11447 2190 2189 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11448 5183 2190 2189 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11449 2192 2191 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11450 5183 2192 2191 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11451 2194 2193 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11452 5183 2194 2193 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11453 2196 2195 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11454 5183 2196 2195 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11455 2198 2197 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11456 5183 2198 2197 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11457 2200 2199 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11458 5183 2200 2199 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11459 2202 2201 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11460 5183 2202 2201 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11461 2204 2203 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11462 5183 2204 2203 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11463 2206 2205 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11464 5183 2206 2205 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11465 2208 2207 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11466 5183 2208 2207 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11467 2210 2209 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11468 5183 2210 2209 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11469 2212 2211 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11470 5183 2212 2211 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11471 2214 2213 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11472 5183 2214 2213 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11473 2216 2215 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11474 5183 2216 2215 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11475 2218 2217 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11476 5183 2218 2217 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11477 2220 2219 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11478 5183 2220 2219 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11479 2222 2221 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11480 5183 2222 2221 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11481 2224 2223 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11482 5183 2224 2223 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11483 2226 2225 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11484 5183 2226 2225 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11485 2228 2227 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11486 5183 2228 2227 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11487 2230 2229 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11488 5183 2230 2229 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11489 2232 2231 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11490 5183 2232 2231 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11491 2234 2233 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11492 5183 2234 2233 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11493 2236 2235 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11494 5183 2236 2235 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11495 2238 2237 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11496 5183 2238 2237 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11497 2240 2239 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11498 5183 2240 2239 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11499 2242 2241 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11500 5183 2242 2241 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11501 2244 2243 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11502 5183 2244 2243 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11503 2246 2245 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11504 5183 2246 2245 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11505 2248 2247 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11506 5183 2248 2247 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11507 2250 2249 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11508 5183 2250 2249 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11509 2252 2251 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11510 5183 2252 2251 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11511 2254 2253 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11512 5183 2254 2253 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11513 2256 2255 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11514 5183 2256 2255 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11515 2258 2257 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11516 5183 2258 2257 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11517 2260 2259 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11518 5183 2260 2259 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11519 2262 2261 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11520 5183 2262 2261 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11521 2264 2263 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11522 5183 2264 2263 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11523 2266 2265 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11524 5183 2266 2265 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11525 2268 2267 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11526 5183 2268 2267 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11527 2270 2269 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11528 5183 2270 2269 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11529 2272 2271 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11530 5183 2272 2271 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11531 2274 2273 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11532 5183 2274 2273 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11533 2276 2275 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11534 5183 2276 2275 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11535 2278 2277 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11536 5183 2278 2277 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11537 2280 2279 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11538 5183 2280 2279 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11539 2282 2281 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11540 5183 2282 2281 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11541 2284 2283 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11542 5183 2284 2283 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11543 2286 2285 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11544 5183 2286 2285 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11545 2288 2287 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11546 5183 2288 2287 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11547 2290 2289 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11548 5183 2290 2289 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11549 2292 2291 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11550 5183 2292 2291 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11551 2294 2293 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11552 5183 2294 2293 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11553 2296 2295 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11554 5183 2296 2295 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11555 2298 2297 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11556 5183 2298 2297 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11557 2300 2299 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11558 5183 2300 2299 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11559 2302 2301 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11560 5183 2302 2301 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11561 2304 2303 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11562 5183 2304 2303 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11563 2306 2305 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11564 5183 2306 2305 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11565 2308 2307 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11566 5183 2308 2307 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11567 2310 2309 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11568 5183 2310 2309 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11569 2312 2311 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11570 5183 2312 2311 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11571 2314 2313 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11572 5183 2314 2313 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11573 2316 2315 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11574 5183 2316 2315 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11575 2318 2317 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11576 5183 2318 2317 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11577 2320 2319 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11578 5183 2320 2319 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11579 2322 2321 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11580 5183 2322 2321 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11581 2324 2323 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11582 5183 2324 2323 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11583 2326 2325 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11584 5183 2326 2325 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11585 2328 2327 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11586 5183 2328 2327 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11587 2330 2329 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11588 5183 2330 2329 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11589 2332 2331 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11590 5183 2332 2331 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11591 2334 2333 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11592 5183 2334 2333 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11593 2336 2335 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11594 5183 2336 2335 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11595 2338 2337 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11596 5183 2338 2337 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11597 2340 2339 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11598 5183 2340 2339 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11599 2342 2341 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11600 5183 2342 2341 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11601 2344 2343 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11602 5183 2344 2343 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11603 2346 2345 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11604 5183 2346 2345 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11605 2348 2347 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11606 5183 2348 2347 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11607 2350 2349 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11608 5183 2350 2349 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11609 2352 2351 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11610 5183 2352 2351 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11611 2354 2353 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11612 5183 2354 2353 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11613 2356 2355 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11614 5183 2356 2355 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11615 2358 2357 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11616 5183 2358 2357 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11617 2360 2359 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11618 5183 2360 2359 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11619 2362 2361 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11620 5183 2362 2361 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11621 2364 2363 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11622 5183 2364 2363 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11623 2366 2365 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11624 5183 2366 2365 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11625 2368 2367 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11626 5183 2368 2367 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11627 2370 2369 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11628 5183 2370 2369 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11629 2372 2371 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11630 5183 2372 2371 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11631 2374 2373 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11632 5183 2374 2373 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11633 2376 2375 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11634 5183 2376 2375 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11635 2378 2377 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11636 5183 2378 2377 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11637 2380 2379 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11638 5183 2380 2379 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11639 2382 2381 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11640 5183 2382 2381 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11641 2384 2383 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11642 5183 2384 2383 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11643 2386 2385 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11644 5183 2386 2385 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11645 2388 2387 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11646 5183 2388 2387 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11647 2390 2389 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11648 5183 2390 2389 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11649 2392 2391 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11650 5183 2392 2391 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11651 2394 2393 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11652 5183 2394 2393 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11653 2396 2395 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11654 5183 2396 2395 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11655 2398 2397 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11656 5183 2398 2397 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11657 2400 2399 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11658 5183 2400 2399 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11659 2402 2401 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11660 5183 2402 2401 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11661 2404 2403 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11662 5183 2404 2403 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11663 2406 2405 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11664 5183 2406 2405 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11665 2408 2407 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11666 5183 2408 2407 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11667 2410 2409 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11668 5183 2410 2409 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11669 2412 2411 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11670 5183 2412 2411 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11671 2414 2413 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11672 5183 2414 2413 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11673 2416 2415 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11674 5183 2416 2415 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11675 2418 2417 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11676 5183 2418 2417 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11677 2420 2419 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11678 5183 2420 2419 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11679 2422 2421 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11680 5183 2422 2421 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11681 2424 2423 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11682 5183 2424 2423 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11683 2426 2425 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11684 5183 2426 2425 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11685 2428 2427 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11686 5183 2428 2427 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11687 2430 2429 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11688 5183 2430 2429 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11689 2432 2431 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11690 5183 2432 2431 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11691 2434 2433 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11692 5183 2434 2433 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11693 2436 2435 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11694 5183 2436 2435 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11695 2438 2437 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11696 5183 2438 2437 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11697 2440 2439 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11698 5183 2440 2439 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11699 2442 2441 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11700 5183 2442 2441 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11701 2444 2443 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11702 5183 2444 2443 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11703 2446 2445 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11704 5183 2446 2445 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11705 2448 2447 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11706 5183 2448 2447 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11707 2450 2449 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11708 5183 2450 2449 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11709 2452 2451 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11710 5183 2452 2451 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11711 2454 2453 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11712 5183 2454 2453 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11713 2456 2455 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11714 5183 2456 2455 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11715 2458 2457 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11716 5183 2458 2457 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11717 2460 2459 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11718 5183 2460 2459 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11719 2462 2461 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11720 5183 2462 2461 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11721 2464 2463 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11722 5183 2464 2463 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11723 2466 2465 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11724 5183 2466 2465 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11725 2468 2467 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11726 5183 2468 2467 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11727 2470 2469 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11728 5183 2470 2469 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11729 2472 2471 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11730 5183 2472 2471 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11731 2474 2473 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11732 5183 2474 2473 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11733 2476 2475 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11734 5183 2476 2475 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11735 2478 2477 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11736 5183 2478 2477 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11737 2480 2479 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11738 5183 2480 2479 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11739 2482 2481 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11740 5183 2482 2481 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11741 2484 2483 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11742 5183 2484 2483 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11743 2486 2485 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11744 5183 2486 2485 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11745 2488 2487 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11746 5183 2488 2487 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11747 2490 2489 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11748 5183 2490 2489 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11749 2492 2491 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11750 5183 2492 2491 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11751 2494 2493 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11752 5183 2494 2493 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11753 2496 2495 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11754 5183 2496 2495 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11755 2498 2497 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11756 5183 2498 2497 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11757 2500 2499 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11758 5183 2500 2499 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11759 2502 2501 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11760 5183 2502 2501 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11761 2504 2503 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11762 5183 2504 2503 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11763 2506 2505 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11764 5183 2506 2505 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11765 2508 2507 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11766 5183 2508 2507 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11767 2510 2509 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11768 5183 2510 2509 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11769 2512 2511 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11770 5183 2512 2511 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11771 2514 2513 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11772 5183 2514 2513 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11773 2516 2515 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11774 5183 2516 2515 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11775 2525 2517 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11776 5183 2517 2517 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11777 2519 2519 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11778 5183 2519 2518 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11779 2520 2521 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11780 5183 2521 2521 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11781 2522 5189 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11782 5183 2524 2523 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11783 2524 5189 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11784 5183 5189 2524 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11785 5189 2527 5183 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_11786 5183 2527 5189 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_11787 5183 3074 2527 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_11788 2527 2525 5183 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_11789 2527 3077 2526 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_11790 2528 2530 5183 5183 pmos L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_11791 5183 2530 2528 5183 pmos L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_11792 2528 2530 5183 5183 pmos L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_11793 5183 2530 2528 5183 pmos L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_11794 2529 2532 5183 5183 pmos L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_11795 5183 2532 2529 5183 pmos L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_11796 2529 2532 5183 5183 pmos L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_11797 5183 2532 2529 5183 pmos L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_11798 2531 3085 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_11799 5183 2531 2530 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11800 2530 3086 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11801 5183 2531 2532 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11802 2532 3086 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11803 5183 2546 2533 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11804 5183 3085 2546 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11805 5183 2537 2546 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11806 2546 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11807 5183 2537 2544 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11808 2544 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11809 5183 3085 2544 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11810 5183 2544 2535 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11811 2542 2537 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11812 5183 3067 2542 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11813 2542 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11814 2548 2537 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11815 5183 3071 2548 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11816 2548 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11817 5183 2542 2534 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11818 2536 2548 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11819 2533 2546 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11820 2534 2542 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11821 2535 2544 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11822 5183 2548 2536 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11823 2537 2540 2538 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_11824 2538 2539 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_11825 2539 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11826 5183 3060 2539 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11827 5183 3054 2540 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11828 2540 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11829 5183 3048 2540 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11830 2541 2542 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11831 5183 2542 2541 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11832 2543 2544 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11833 5183 2544 2543 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11834 2545 2546 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11835 5183 2546 2545 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11836 2547 2548 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11837 5183 2548 2547 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11838 5183 2562 2549 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11839 5183 3085 2562 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11840 5183 2553 2562 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11841 2562 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11842 5183 2553 2560 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11843 2560 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11844 5183 3085 2560 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11845 5183 2560 2551 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11846 2558 2553 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11847 5183 3067 2558 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11848 2558 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11849 2564 2553 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11850 5183 3071 2564 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11851 2564 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11852 5183 2558 2550 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11853 2552 2564 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11854 2549 2562 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11855 2550 2558 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11856 2551 2560 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11857 5183 2564 2552 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11858 2553 2556 2554 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_11859 2554 2555 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_11860 2555 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11861 5183 3060 2555 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11862 5183 3054 2556 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11863 2556 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11864 5183 3047 2556 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11865 2557 2558 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11866 5183 2558 2557 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11867 2559 2560 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11868 5183 2560 2559 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11869 2561 2562 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11870 5183 2562 2561 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11871 2563 2564 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11872 5183 2564 2563 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11873 5183 2578 2565 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11874 5183 3085 2578 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11875 5183 2569 2578 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11876 2578 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11877 5183 2569 2576 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11878 2576 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11879 5183 3085 2576 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11880 5183 2576 2567 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11881 2574 2569 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11882 5183 3067 2574 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11883 2574 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11884 2580 2569 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11885 5183 3071 2580 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11886 2580 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11887 5183 2574 2566 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11888 2568 2580 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11889 2565 2578 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11890 2566 2574 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11891 2567 2576 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11892 5183 2580 2568 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11893 2569 2572 2570 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_11894 2570 2571 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_11895 2571 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11896 5183 3060 2571 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11897 5183 3054 2572 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11898 2572 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11899 5183 3048 2572 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11900 2573 2574 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11901 5183 2574 2573 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11902 2575 2576 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11903 5183 2576 2575 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11904 2577 2578 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11905 5183 2578 2577 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11906 2579 2580 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11907 5183 2580 2579 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11908 5183 2594 2581 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11909 5183 3085 2594 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11910 5183 2585 2594 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11911 2594 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11912 5183 2585 2592 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11913 2592 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11914 5183 3085 2592 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11915 5183 2592 2583 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11916 2590 2585 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11917 5183 3067 2590 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11918 2590 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11919 2596 2585 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11920 5183 3071 2596 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11921 2596 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11922 5183 2590 2582 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11923 2584 2596 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11924 2581 2594 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11925 2582 2590 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11926 2583 2592 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11927 5183 2596 2584 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11928 2585 2588 2586 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_11929 2586 2587 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_11930 2587 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11931 5183 3060 2587 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11932 5183 3054 2588 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11933 2588 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11934 5183 3047 2588 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11935 2589 2590 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11936 5183 2590 2589 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11937 2591 2592 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11938 5183 2592 2591 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11939 2593 2594 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11940 5183 2594 2593 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11941 2595 2596 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11942 5183 2596 2595 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11943 5183 2610 2597 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11944 5183 3085 2610 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11945 5183 2601 2610 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11946 2610 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11947 5183 2601 2608 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11948 2608 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11949 5183 3085 2608 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11950 5183 2608 2599 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11951 2606 2601 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11952 5183 3067 2606 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11953 2606 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11954 2612 2601 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11955 5183 3071 2612 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11956 2612 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11957 5183 2606 2598 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11958 2600 2612 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11959 2597 2610 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11960 2598 2606 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11961 2599 2608 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11962 5183 2612 2600 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11963 2601 2604 2602 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_11964 2602 2603 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_11965 2603 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11966 5183 3060 2603 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11967 5183 3053 2604 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11968 2604 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11969 5183 3048 2604 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_11970 2605 2606 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11971 5183 2606 2605 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11972 2607 2608 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11973 5183 2608 2607 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11974 2609 2610 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11975 5183 2610 2609 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11976 2611 2612 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11977 5183 2612 2611 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11978 5183 2626 2613 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11979 5183 3085 2626 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11980 5183 2617 2626 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11981 2626 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11982 5183 2617 2624 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11983 2624 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11984 5183 3085 2624 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11985 5183 2624 2615 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11986 2622 2617 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11987 5183 3067 2622 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11988 2622 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11989 2628 2617 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11990 5183 3071 2628 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11991 2628 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_11992 5183 2622 2614 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11993 2616 2628 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11994 2613 2626 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11995 2614 2622 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11996 2615 2624 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11997 5183 2628 2616 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_11998 2617 2620 2618 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_11999 2618 2619 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12000 2619 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12001 5183 3060 2619 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12002 5183 3053 2620 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12003 2620 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12004 5183 3047 2620 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12005 2621 2622 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12006 5183 2622 2621 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12007 2623 2624 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12008 5183 2624 2623 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12009 2625 2626 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12010 5183 2626 2625 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12011 2627 2628 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12012 5183 2628 2627 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12013 5183 2642 2629 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12014 5183 3085 2642 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12015 5183 2633 2642 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12016 2642 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12017 5183 2633 2640 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12018 2640 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12019 5183 3085 2640 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12020 5183 2640 2631 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12021 2638 2633 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12022 5183 3067 2638 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12023 2638 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12024 2644 2633 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12025 5183 3071 2644 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12026 2644 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12027 5183 2638 2630 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12028 2632 2644 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12029 2629 2642 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12030 2630 2638 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12031 2631 2640 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12032 5183 2644 2632 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12033 2633 2636 2634 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12034 2634 2635 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12035 2635 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12036 5183 3060 2635 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12037 5183 3053 2636 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12038 2636 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12039 5183 3048 2636 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12040 2637 2638 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12041 5183 2638 2637 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12042 2639 2640 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12043 5183 2640 2639 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12044 2641 2642 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12045 5183 2642 2641 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12046 2643 2644 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12047 5183 2644 2643 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12048 5183 2658 2645 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12049 5183 3085 2658 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12050 5183 2649 2658 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12051 2658 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12052 5183 2649 2656 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12053 2656 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12054 5183 3085 2656 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12055 5183 2656 2647 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12056 2654 2649 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12057 5183 3067 2654 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12058 2654 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12059 2660 2649 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12060 5183 3071 2660 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12061 2660 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12062 5183 2654 2646 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12063 2648 2660 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12064 2645 2658 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12065 2646 2654 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12066 2647 2656 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12067 5183 2660 2648 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12068 2649 2652 2650 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12069 2650 2651 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12070 2651 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12071 5183 3060 2651 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12072 5183 3053 2652 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12073 2652 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12074 5183 3047 2652 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12075 2653 2654 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12076 5183 2654 2653 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12077 2655 2656 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12078 5183 2656 2655 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12079 2657 2658 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12080 5183 2658 2657 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12081 2659 2660 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12082 5183 2660 2659 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12083 5183 2674 2661 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12084 5183 3085 2674 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12085 5183 2665 2674 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12086 2674 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12087 5183 2665 2672 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12088 2672 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12089 5183 3085 2672 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12090 5183 2672 2663 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12091 2670 2665 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12092 5183 3067 2670 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12093 2670 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12094 2676 2665 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12095 5183 3071 2676 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12096 2676 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12097 5183 2670 2662 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12098 2664 2676 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12099 2661 2674 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12100 2662 2670 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12101 2663 2672 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12102 5183 2676 2664 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12103 2665 2668 2666 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12104 2666 2667 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12105 2667 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12106 5183 3060 2667 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12107 5183 3054 2668 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12108 2668 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12109 5183 3048 2668 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12110 2669 2670 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12111 5183 2670 2669 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12112 2671 2672 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12113 5183 2672 2671 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12114 2673 2674 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12115 5183 2674 2673 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12116 2675 2676 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12117 5183 2676 2675 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12118 5183 2690 2677 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12119 5183 3085 2690 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12120 5183 2681 2690 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12121 2690 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12122 5183 2681 2688 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12123 2688 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12124 5183 3085 2688 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12125 5183 2688 2679 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12126 2686 2681 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12127 5183 3067 2686 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12128 2686 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12129 2692 2681 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12130 5183 3071 2692 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12131 2692 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12132 5183 2686 2678 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12133 2680 2692 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12134 2677 2690 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12135 2678 2686 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12136 2679 2688 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12137 5183 2692 2680 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12138 2681 2684 2682 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12139 2682 2683 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12140 2683 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12141 5183 3060 2683 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12142 5183 3054 2684 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12143 2684 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12144 5183 3047 2684 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12145 2685 2686 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12146 5183 2686 2685 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12147 2687 2688 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12148 5183 2688 2687 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12149 2689 2690 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12150 5183 2690 2689 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12151 2691 2692 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12152 5183 2692 2691 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12153 5183 2706 2693 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12154 5183 3085 2706 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12155 5183 2697 2706 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12156 2706 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12157 5183 2697 2704 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12158 2704 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12159 5183 3085 2704 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12160 5183 2704 2695 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12161 2702 2697 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12162 5183 3067 2702 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12163 2702 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12164 2708 2697 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12165 5183 3071 2708 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12166 2708 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12167 5183 2702 2694 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12168 2696 2708 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12169 2693 2706 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12170 2694 2702 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12171 2695 2704 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12172 5183 2708 2696 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12173 2697 2700 2698 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12174 2698 2699 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12175 2699 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12176 5183 3060 2699 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12177 5183 3054 2700 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12178 2700 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12179 5183 3048 2700 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12180 2701 2702 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12181 5183 2702 2701 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12182 2703 2704 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12183 5183 2704 2703 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12184 2705 2706 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12185 5183 2706 2705 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12186 2707 2708 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12187 5183 2708 2707 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12188 5183 2722 2709 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12189 5183 3085 2722 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12190 5183 2713 2722 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12191 2722 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12192 5183 2713 2720 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12193 2720 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12194 5183 3085 2720 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12195 5183 2720 2711 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12196 2718 2713 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12197 5183 3067 2718 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12198 2718 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12199 2724 2713 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12200 5183 3071 2724 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12201 2724 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12202 5183 2718 2710 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12203 2712 2724 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12204 2709 2722 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12205 2710 2718 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12206 2711 2720 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12207 5183 2724 2712 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12208 2713 2716 2714 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12209 2714 2715 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12210 2715 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12211 5183 3060 2715 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12212 5183 3054 2716 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12213 2716 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12214 5183 3047 2716 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12215 2717 2718 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12216 5183 2718 2717 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12217 2719 2720 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12218 5183 2720 2719 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12219 2721 2722 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12220 5183 2722 2721 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12221 2723 2724 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12222 5183 2724 2723 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12223 5183 2738 2725 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12224 5183 3085 2738 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12225 5183 2729 2738 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12226 2738 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12227 5183 2729 2736 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12228 2736 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12229 5183 3085 2736 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12230 5183 2736 2727 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12231 2734 2729 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12232 5183 3067 2734 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12233 2734 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12234 2740 2729 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12235 5183 3071 2740 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12236 2740 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12237 5183 2734 2726 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12238 2728 2740 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12239 2725 2738 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12240 2726 2734 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12241 2727 2736 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12242 5183 2740 2728 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12243 2729 2732 2730 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12244 2730 2731 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12245 2731 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12246 5183 3060 2731 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12247 5183 3053 2732 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12248 2732 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12249 5183 3048 2732 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12250 2733 2734 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12251 5183 2734 2733 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12252 2735 2736 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12253 5183 2736 2735 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12254 2737 2738 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12255 5183 2738 2737 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12256 2739 2740 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12257 5183 2740 2739 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12258 5183 2754 2741 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12259 5183 3085 2754 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12260 5183 2745 2754 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12261 2754 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12262 5183 2745 2752 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12263 2752 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12264 5183 3085 2752 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12265 5183 2752 2743 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12266 2750 2745 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12267 5183 3067 2750 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12268 2750 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12269 2756 2745 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12270 5183 3071 2756 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12271 2756 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12272 5183 2750 2742 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12273 2744 2756 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12274 2741 2754 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12275 2742 2750 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12276 2743 2752 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12277 5183 2756 2744 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12278 2745 2748 2746 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12279 2746 2747 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12280 2747 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12281 5183 3060 2747 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12282 5183 3053 2748 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12283 2748 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12284 5183 3047 2748 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12285 2749 2750 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12286 5183 2750 2749 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12287 2751 2752 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12288 5183 2752 2751 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12289 2753 2754 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12290 5183 2754 2753 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12291 2755 2756 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12292 5183 2756 2755 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12293 5183 2770 2757 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12294 5183 3085 2770 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12295 5183 2761 2770 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12296 2770 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12297 5183 2761 2768 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12298 2768 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12299 5183 3085 2768 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12300 5183 2768 2759 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12301 2766 2761 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12302 5183 3067 2766 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12303 2766 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12304 2772 2761 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12305 5183 3071 2772 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12306 2772 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12307 5183 2766 2758 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12308 2760 2772 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12309 2757 2770 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12310 2758 2766 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12311 2759 2768 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12312 5183 2772 2760 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12313 2761 2764 2762 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12314 2762 2763 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12315 2763 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12316 5183 3060 2763 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12317 5183 3053 2764 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12318 2764 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12319 5183 3048 2764 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12320 2765 2766 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12321 5183 2766 2765 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12322 2767 2768 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12323 5183 2768 2767 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12324 2769 2770 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12325 5183 2770 2769 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12326 2771 2772 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12327 5183 2772 2771 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12328 5183 2786 2773 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12329 5183 3085 2786 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12330 5183 2777 2786 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12331 2786 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12332 5183 2777 2784 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12333 2784 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12334 5183 3085 2784 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12335 5183 2784 2775 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12336 2782 2777 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12337 5183 3067 2782 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12338 2782 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12339 2788 2777 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12340 5183 3071 2788 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12341 2788 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12342 5183 2782 2774 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12343 2776 2788 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12344 2773 2786 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12345 2774 2782 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12346 2775 2784 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12347 5183 2788 2776 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12348 2777 2780 2778 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12349 2778 2779 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12350 2779 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12351 5183 3060 2779 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12352 5183 3053 2780 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12353 2780 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12354 5183 3047 2780 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12355 2781 2782 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12356 5183 2782 2781 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12357 2783 2784 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12358 5183 2784 2783 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12359 2785 2786 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12360 5183 2786 2785 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12361 2787 2788 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12362 5183 2788 2787 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12363 5183 2802 2789 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12364 5183 3085 2802 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12365 5183 2793 2802 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12366 2802 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12367 5183 2793 2800 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12368 2800 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12369 5183 3085 2800 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12370 5183 2800 2791 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12371 2798 2793 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12372 5183 3067 2798 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12373 2798 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12374 2804 2793 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12375 5183 3071 2804 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12376 2804 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12377 5183 2798 2790 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12378 2792 2804 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12379 2789 2802 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12380 2790 2798 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12381 2791 2800 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12382 5183 2804 2792 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12383 2793 2796 2794 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12384 2794 2795 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12385 2795 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12386 5183 3059 2795 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12387 5183 3054 2796 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12388 2796 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12389 5183 3048 2796 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12390 2797 2798 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12391 5183 2798 2797 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12392 2799 2800 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12393 5183 2800 2799 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12394 2801 2802 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12395 5183 2802 2801 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12396 2803 2804 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12397 5183 2804 2803 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12398 5183 2818 2805 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12399 5183 3085 2818 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12400 5183 2809 2818 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12401 2818 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12402 5183 2809 2816 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12403 2816 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12404 5183 3085 2816 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12405 5183 2816 2807 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12406 2814 2809 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12407 5183 3067 2814 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12408 2814 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12409 2820 2809 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12410 5183 3071 2820 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12411 2820 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12412 5183 2814 2806 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12413 2808 2820 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12414 2805 2818 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12415 2806 2814 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12416 2807 2816 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12417 5183 2820 2808 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12418 2809 2812 2810 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12419 2810 2811 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12420 2811 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12421 5183 3059 2811 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12422 5183 3054 2812 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12423 2812 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12424 5183 3047 2812 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12425 2813 2814 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12426 5183 2814 2813 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12427 2815 2816 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12428 5183 2816 2815 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12429 2817 2818 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12430 5183 2818 2817 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12431 2819 2820 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12432 5183 2820 2819 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12433 5183 2834 2821 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12434 5183 3085 2834 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12435 5183 2825 2834 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12436 2834 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12437 5183 2825 2832 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12438 2832 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12439 5183 3085 2832 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12440 5183 2832 2823 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12441 2830 2825 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12442 5183 3067 2830 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12443 2830 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12444 2836 2825 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12445 5183 3071 2836 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12446 2836 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12447 5183 2830 2822 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12448 2824 2836 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12449 2821 2834 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12450 2822 2830 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12451 2823 2832 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12452 5183 2836 2824 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12453 2825 2828 2826 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12454 2826 2827 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12455 2827 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12456 5183 3059 2827 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12457 5183 3054 2828 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12458 2828 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12459 5183 3048 2828 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12460 2829 2830 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12461 5183 2830 2829 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12462 2831 2832 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12463 5183 2832 2831 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12464 2833 2834 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12465 5183 2834 2833 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12466 2835 2836 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12467 5183 2836 2835 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12468 5183 2850 2837 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12469 5183 3085 2850 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12470 5183 2841 2850 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12471 2850 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12472 5183 2841 2848 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12473 2848 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12474 5183 3085 2848 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12475 5183 2848 2839 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12476 2846 2841 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12477 5183 3067 2846 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12478 2846 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12479 2852 2841 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12480 5183 3071 2852 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12481 2852 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12482 5183 2846 2838 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12483 2840 2852 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12484 2837 2850 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12485 2838 2846 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12486 2839 2848 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12487 5183 2852 2840 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12488 2841 2844 2842 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12489 2842 2843 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12490 2843 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12491 5183 3059 2843 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12492 5183 3054 2844 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12493 2844 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12494 5183 3047 2844 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12495 2845 2846 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12496 5183 2846 2845 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12497 2847 2848 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12498 5183 2848 2847 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12499 2849 2850 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12500 5183 2850 2849 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12501 2851 2852 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12502 5183 2852 2851 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12503 5183 2866 2853 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12504 5183 3085 2866 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12505 5183 2857 2866 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12506 2866 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12507 5183 2857 2864 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12508 2864 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12509 5183 3085 2864 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12510 5183 2864 2855 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12511 2862 2857 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12512 5183 3067 2862 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12513 2862 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12514 2868 2857 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12515 5183 3071 2868 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12516 2868 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12517 5183 2862 2854 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12518 2856 2868 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12519 2853 2866 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12520 2854 2862 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12521 2855 2864 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12522 5183 2868 2856 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12523 2857 2860 2858 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12524 2858 2859 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12525 2859 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12526 5183 3059 2859 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12527 5183 3053 2860 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12528 2860 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12529 5183 3048 2860 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12530 2861 2862 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12531 5183 2862 2861 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12532 2863 2864 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12533 5183 2864 2863 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12534 2865 2866 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12535 5183 2866 2865 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12536 2867 2868 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12537 5183 2868 2867 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12538 5183 2882 2869 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12539 5183 3085 2882 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12540 5183 2873 2882 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12541 2882 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12542 5183 2873 2880 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12543 2880 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12544 5183 3085 2880 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12545 5183 2880 2871 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12546 2878 2873 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12547 5183 3067 2878 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12548 2878 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12549 2884 2873 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12550 5183 3071 2884 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12551 2884 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12552 5183 2878 2870 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12553 2872 2884 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12554 2869 2882 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12555 2870 2878 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12556 2871 2880 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12557 5183 2884 2872 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12558 2873 2876 2874 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12559 2874 2875 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12560 2875 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12561 5183 3059 2875 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12562 5183 3053 2876 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12563 2876 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12564 5183 3047 2876 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12565 2877 2878 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12566 5183 2878 2877 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12567 2879 2880 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12568 5183 2880 2879 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12569 2881 2882 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12570 5183 2882 2881 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12571 2883 2884 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12572 5183 2884 2883 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12573 5183 2898 2885 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12574 5183 3085 2898 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12575 5183 2889 2898 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12576 2898 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12577 5183 2889 2896 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12578 2896 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12579 5183 3085 2896 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12580 5183 2896 2887 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12581 2894 2889 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12582 5183 3067 2894 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12583 2894 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12584 2900 2889 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12585 5183 3071 2900 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12586 2900 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12587 5183 2894 2886 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12588 2888 2900 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12589 2885 2898 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12590 2886 2894 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12591 2887 2896 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12592 5183 2900 2888 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12593 2889 2892 2890 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12594 2890 2891 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12595 2891 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12596 5183 3059 2891 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12597 5183 3053 2892 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12598 2892 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12599 5183 3048 2892 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12600 2893 2894 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12601 5183 2894 2893 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12602 2895 2896 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12603 5183 2896 2895 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12604 2897 2898 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12605 5183 2898 2897 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12606 2899 2900 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12607 5183 2900 2899 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12608 5183 2914 2901 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12609 5183 3085 2914 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12610 5183 2905 2914 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12611 2914 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12612 5183 2905 2912 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12613 2912 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12614 5183 3085 2912 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12615 5183 2912 2903 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12616 2910 2905 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12617 5183 3067 2910 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12618 2910 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12619 2916 2905 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12620 5183 3071 2916 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12621 2916 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12622 5183 2910 2902 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12623 2904 2916 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12624 2901 2914 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12625 2902 2910 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12626 2903 2912 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12627 5183 2916 2904 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12628 2905 2908 2906 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12629 2906 2907 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12630 2907 3057 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12631 5183 3059 2907 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12632 5183 3053 2908 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12633 2908 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12634 5183 3047 2908 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12635 2909 2910 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12636 5183 2910 2909 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12637 2911 2912 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12638 5183 2912 2911 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12639 2913 2914 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12640 5183 2914 2913 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12641 2915 2916 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12642 5183 2916 2915 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12643 5183 2930 2917 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12644 5183 3085 2930 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12645 5183 2921 2930 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12646 2930 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12647 5183 2921 2928 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12648 2928 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12649 5183 3085 2928 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12650 5183 2928 2919 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12651 2926 2921 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12652 5183 3067 2926 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12653 2926 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12654 2932 2921 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12655 5183 3071 2932 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12656 2932 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12657 5183 2926 2918 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12658 2920 2932 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12659 2917 2930 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12660 2918 2926 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12661 2919 2928 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12662 5183 2932 2920 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12663 2921 2924 2922 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12664 2922 2923 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12665 2923 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12666 5183 3059 2923 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12667 5183 3054 2924 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12668 2924 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12669 5183 3048 2924 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12670 2925 2926 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12671 5183 2926 2925 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12672 2927 2928 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12673 5183 2928 2927 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12674 2929 2930 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12675 5183 2930 2929 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12676 2931 2932 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12677 5183 2932 2931 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12678 5183 2946 2933 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12679 5183 3085 2946 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12680 5183 2937 2946 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12681 2946 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12682 5183 2937 2944 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12683 2944 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12684 5183 3085 2944 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12685 5183 2944 2935 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12686 2942 2937 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12687 5183 3067 2942 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12688 2942 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12689 2948 2937 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12690 5183 3071 2948 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12691 2948 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12692 5183 2942 2934 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12693 2936 2948 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12694 2933 2946 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12695 2934 2942 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12696 2935 2944 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12697 5183 2948 2936 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12698 2937 2940 2938 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12699 2938 2939 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12700 2939 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12701 5183 3059 2939 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12702 5183 3054 2940 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12703 2940 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12704 5183 3047 2940 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12705 2941 2942 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12706 5183 2942 2941 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12707 2943 2944 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12708 5183 2944 2943 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12709 2945 2946 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12710 5183 2946 2945 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12711 2947 2948 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12712 5183 2948 2947 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12713 5183 2962 2949 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12714 5183 3085 2962 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12715 5183 2953 2962 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12716 2962 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12717 5183 2953 2960 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12718 2960 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12719 5183 3085 2960 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12720 5183 2960 2951 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12721 2958 2953 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12722 5183 3067 2958 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12723 2958 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12724 2964 2953 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12725 5183 3071 2964 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12726 2964 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12727 5183 2958 2950 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12728 2952 2964 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12729 2949 2962 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12730 2950 2958 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12731 2951 2960 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12732 5183 2964 2952 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12733 2953 2956 2954 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12734 2954 2955 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12735 2955 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12736 5183 3059 2955 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12737 5183 3054 2956 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12738 2956 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12739 5183 3048 2956 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12740 2957 2958 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12741 5183 2958 2957 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12742 2959 2960 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12743 5183 2960 2959 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12744 2961 2962 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12745 5183 2962 2961 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12746 2963 2964 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12747 5183 2964 2963 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12748 5183 2978 2965 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12749 5183 3085 2978 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12750 5183 2969 2978 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12751 2978 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12752 5183 2969 2976 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12753 2976 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12754 5183 3085 2976 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12755 5183 2976 2967 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12756 2974 2969 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12757 5183 3067 2974 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12758 2974 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12759 2980 2969 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12760 5183 3071 2980 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12761 2980 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12762 5183 2974 2966 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12763 2968 2980 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12764 2965 2978 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12765 2966 2974 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12766 2967 2976 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12767 5183 2980 2968 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12768 2969 2972 2970 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12769 2970 2971 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12770 2971 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12771 5183 3059 2971 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12772 5183 3054 2972 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12773 2972 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12774 5183 3047 2972 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12775 2973 2974 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12776 5183 2974 2973 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12777 2975 2976 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12778 5183 2976 2975 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12779 2977 2978 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12780 5183 2978 2977 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12781 2979 2980 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12782 5183 2980 2979 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12783 5183 2994 2981 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12784 5183 3085 2994 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12785 5183 2985 2994 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12786 2994 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12787 5183 2985 2992 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12788 2992 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12789 5183 3085 2992 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12790 5183 2992 2983 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12791 2990 2985 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12792 5183 3067 2990 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12793 2990 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12794 2996 2985 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12795 5183 3071 2996 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12796 2996 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12797 5183 2990 2982 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12798 2984 2996 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12799 2981 2994 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12800 2982 2990 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12801 2983 2992 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12802 5183 2996 2984 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12803 2985 2988 2986 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12804 2986 2987 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12805 2987 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12806 5183 3059 2987 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12807 5183 3053 2988 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12808 2988 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12809 5183 3048 2988 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12810 2989 2990 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12811 5183 2990 2989 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12812 2991 2992 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12813 5183 2992 2991 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12814 2993 2994 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12815 5183 2994 2993 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12816 2995 2996 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12817 5183 2996 2995 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12818 5183 3010 2997 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12819 5183 3085 3010 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12820 5183 3001 3010 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12821 3010 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12822 5183 3001 3008 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12823 3008 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12824 5183 3085 3008 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12825 5183 3008 2999 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12826 3006 3001 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12827 5183 3067 3006 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12828 3006 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12829 3012 3001 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12830 5183 3071 3012 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12831 3012 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12832 5183 3006 2998 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12833 3000 3012 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12834 2997 3010 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12835 2998 3006 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12836 2999 3008 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12837 5183 3012 3000 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12838 3001 3004 3002 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12839 3002 3003 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12840 3003 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12841 5183 3059 3003 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12842 5183 3053 3004 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12843 3004 3051 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12844 5183 3047 3004 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12845 3005 3006 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12846 5183 3006 3005 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12847 3007 3008 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12848 5183 3008 3007 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12849 3009 3010 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12850 5183 3010 3009 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12851 3011 3012 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12852 5183 3012 3011 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12853 5183 3026 3013 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12854 5183 3085 3026 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12855 5183 3017 3026 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12856 3026 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12857 5183 3017 3024 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12858 3024 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12859 5183 3085 3024 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12860 5183 3024 3015 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12861 3022 3017 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12862 5183 3067 3022 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12863 3022 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12864 3028 3017 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12865 5183 3071 3028 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12866 3028 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12867 5183 3022 3014 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12868 3016 3028 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12869 3013 3026 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12870 3014 3022 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12871 3015 3024 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12872 5183 3028 3016 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12873 3017 3020 3018 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12874 3018 3019 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12875 3019 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12876 5183 3059 3019 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12877 5183 3053 3020 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12878 3020 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12879 5183 3048 3020 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12880 3021 3022 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12881 5183 3022 3021 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12882 3023 3024 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12883 5183 3024 3023 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12884 3025 3026 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12885 5183 3026 3025 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12886 3027 3028 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12887 5183 3028 3027 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12888 5183 3042 3029 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12889 5183 3085 3042 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12890 5183 3033 3042 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12891 3042 3064 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12892 5183 3033 3040 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12893 3040 3068 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12894 5183 3085 3040 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12895 5183 3040 3031 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12896 3038 3033 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12897 5183 3067 3038 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12898 3038 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12899 3044 3033 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12900 5183 3071 3044 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12901 3044 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12902 5183 3038 3030 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12903 3032 3044 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12904 3029 3042 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12905 3030 3038 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12906 3031 3040 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12907 5183 3044 3032 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12908 3033 3036 3034 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12909 3034 3035 5183 5183 pmos L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_12910 3035 3056 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12911 5183 3059 3035 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12912 5183 3053 3036 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12913 3036 3050 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12914 5183 3047 3036 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12915 3037 3038 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12916 5183 3038 3037 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12917 3039 3040 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12918 5183 3040 3039 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12919 3041 3042 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12920 5183 3042 3041 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12921 3043 3044 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12922 5183 3044 3043 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12923 5183 3072 3045 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12924 3046 3073 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12925 3047 5198 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12926 5183 3049 3048 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12927 5183 5198 3049 5183 pmos L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_12928 3050 5197 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12929 5183 3052 3051 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12930 5183 5197 3052 5183 pmos L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_12931 3053 5196 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12932 5183 3055 3054 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12933 5183 5196 3055 5183 pmos L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_12934 3056 5195 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12935 5183 3058 3057 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12936 5183 5195 3058 5183 pmos L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_12937 3059 5194 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12938 5183 3061 3060 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12939 5183 5194 3061 5183 pmos L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_12940 5183 5200 3062 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12941 3063 5199 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12942 5183 5200 3070 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12943 3070 5199 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12944 5183 5200 3069 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12945 3065 3063 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12946 5183 3062 3065 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12947 3066 5199 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12948 5183 3062 3066 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12949 3069 3063 5183 5183 pmos L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_12950 5183 3065 3064 5183 pmos L=1U W=38U AS=76P AD=76P PS=80U PD=80U 
Mtr_12951 3067 3066 5183 5183 pmos L=1U W=38U AS=76P AD=76P PS=80U PD=80U 
Mtr_12952 5183 3069 3068 5183 pmos L=1U W=38U AS=76P AD=76P PS=80U PD=80U 
Mtr_12953 3071 3070 5183 5183 pmos L=1U W=38U AS=76P AD=76P PS=80U PD=80U 
Mtr_12954 3072 3073 5183 5183 pmos L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_12955 5183 5201 3073 5183 pmos L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_12956 3074 3075 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12957 3075 3078 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12958 5183 3075 3074 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12959 5176 3076 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12960 3076 3079 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12961 5183 3076 5176 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12962 3077 3078 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12963 3078 5181 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12964 5183 3085 3078 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12965 5183 3078 3077 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12966 5179 3079 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12967 3079 5181 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12968 5183 3085 3079 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12969 5183 3079 5179 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12970 5183 3080 3081 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12971 5183 3086 3080 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12972 3080 3084 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12973 3081 3080 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12974 5183 3082 3083 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12975 5183 3086 3082 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12976 3082 3084 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12977 3083 3082 5183 5183 pmos L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_12978 3084 3085 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_12979 5183 3086 3085 5183 pmos L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_12980 3085 3086 5183 5183 pmos L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_12981 5183 3086 3085 5183 pmos L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_12982 3085 3086 5183 5183 pmos L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_12983 3086 5193 5183 5183 pmos L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_12984 5183 5184 3086 5183 pmos L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_12985 3088 3087 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12986 5183 3088 3087 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12987 3090 3089 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12988 5183 3090 3089 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12989 3092 3091 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12990 5183 3092 3091 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12991 3094 3093 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12992 5183 3094 3093 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12993 3096 3095 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12994 5183 3096 3095 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12995 3098 3097 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12996 5183 3098 3097 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12997 3100 3099 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12998 5183 3100 3099 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_12999 3102 3101 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13000 5183 3102 3101 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13001 3104 3103 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13002 5183 3104 3103 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13003 3106 3105 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13004 5183 3106 3105 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13005 3108 3107 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13006 5183 3108 3107 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13007 3110 3109 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13008 5183 3110 3109 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13009 3112 3111 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13010 5183 3112 3111 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13011 3114 3113 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13012 5183 3114 3113 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13013 3116 3115 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13014 5183 3116 3115 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13015 3118 3117 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13016 5183 3118 3117 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13017 3120 3119 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13018 5183 3120 3119 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13019 3122 3121 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13020 5183 3122 3121 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13021 3124 3123 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13022 5183 3124 3123 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13023 3126 3125 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13024 5183 3126 3125 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13025 3128 3127 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13026 5183 3128 3127 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13027 3130 3129 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13028 5183 3130 3129 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13029 3132 3131 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13030 5183 3132 3131 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13031 3134 3133 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13032 5183 3134 3133 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13033 3136 3135 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13034 5183 3136 3135 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13035 3138 3137 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13036 5183 3138 3137 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13037 3140 3139 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13038 5183 3140 3139 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13039 3142 3141 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13040 5183 3142 3141 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13041 3144 3143 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13042 5183 3144 3143 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13043 3146 3145 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13044 5183 3146 3145 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13045 3148 3147 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13046 5183 3148 3147 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13047 3150 3149 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13048 5183 3150 3149 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13049 3152 3151 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13050 5183 3152 3151 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13051 3154 3153 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13052 5183 3154 3153 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13053 3156 3155 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13054 5183 3156 3155 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13055 3158 3157 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13056 5183 3158 3157 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13057 3160 3159 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13058 5183 3160 3159 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13059 3162 3161 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13060 5183 3162 3161 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13061 3164 3163 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13062 5183 3164 3163 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13063 3166 3165 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13064 5183 3166 3165 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13065 3168 3167 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13066 5183 3168 3167 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13067 3170 3169 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13068 5183 3170 3169 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13069 3172 3171 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13070 5183 3172 3171 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13071 3174 3173 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13072 5183 3174 3173 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13073 3176 3175 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13074 5183 3176 3175 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13075 3178 3177 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13076 5183 3178 3177 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13077 3180 3179 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13078 5183 3180 3179 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13079 3182 3181 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13080 5183 3182 3181 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13081 3184 3183 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13082 5183 3184 3183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13083 3186 3185 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13084 5183 3186 3185 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13085 3188 3187 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13086 5183 3188 3187 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13087 3190 3189 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13088 5183 3190 3189 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13089 3192 3191 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13090 5183 3192 3191 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13091 3194 3193 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13092 5183 3194 3193 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13093 3196 3195 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13094 5183 3196 3195 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13095 3198 3197 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13096 5183 3198 3197 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13097 3200 3199 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13098 5183 3200 3199 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13099 3202 3201 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13100 5183 3202 3201 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13101 3204 3203 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13102 5183 3204 3203 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13103 3206 3205 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13104 5183 3206 3205 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13105 3208 3207 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13106 5183 3208 3207 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13107 3210 3209 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13108 5183 3210 3209 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13109 3212 3211 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13110 5183 3212 3211 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13111 3214 3213 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13112 5183 3214 3213 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13113 3216 3215 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13114 5183 3216 3215 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13115 3218 3217 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13116 5183 3218 3217 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13117 3220 3219 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13118 5183 3220 3219 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13119 3222 3221 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13120 5183 3222 3221 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13121 3224 3223 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13122 5183 3224 3223 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13123 3226 3225 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13124 5183 3226 3225 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13125 3228 3227 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13126 5183 3228 3227 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13127 3230 3229 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13128 5183 3230 3229 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13129 3232 3231 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13130 5183 3232 3231 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13131 3234 3233 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13132 5183 3234 3233 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13133 3236 3235 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13134 5183 3236 3235 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13135 3238 3237 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13136 5183 3238 3237 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13137 3240 3239 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13138 5183 3240 3239 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13139 3242 3241 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13140 5183 3242 3241 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13141 3244 3243 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13142 5183 3244 3243 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13143 3246 3245 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13144 5183 3246 3245 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13145 3248 3247 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13146 5183 3248 3247 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13147 3250 3249 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13148 5183 3250 3249 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13149 3252 3251 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13150 5183 3252 3251 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13151 3254 3253 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13152 5183 3254 3253 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13153 3256 3255 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13154 5183 3256 3255 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13155 3258 3257 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13156 5183 3258 3257 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13157 3260 3259 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13158 5183 3260 3259 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13159 3262 3261 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13160 5183 3262 3261 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13161 3264 3263 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13162 5183 3264 3263 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13163 3266 3265 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13164 5183 3266 3265 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13165 3268 3267 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13166 5183 3268 3267 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13167 3270 3269 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13168 5183 3270 3269 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13169 3272 3271 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13170 5183 3272 3271 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13171 3274 3273 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13172 5183 3274 3273 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13173 3276 3275 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13174 5183 3276 3275 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13175 3278 3277 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13176 5183 3278 3277 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13177 3280 3279 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13178 5183 3280 3279 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13179 3282 3281 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13180 5183 3282 3281 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13181 3284 3283 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13182 5183 3284 3283 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13183 3286 3285 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13184 5183 3286 3285 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13185 3288 3287 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13186 5183 3288 3287 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13187 3290 3289 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13188 5183 3290 3289 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13189 3292 3291 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13190 5183 3292 3291 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13191 3294 3293 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13192 5183 3294 3293 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13193 3296 3295 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13194 5183 3296 3295 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13195 3298 3297 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13196 5183 3298 3297 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13197 3300 3299 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13198 5183 3300 3299 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13199 3302 3301 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13200 5183 3302 3301 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13201 3304 3303 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13202 5183 3304 3303 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13203 3306 3305 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13204 5183 3306 3305 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13205 3308 3307 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13206 5183 3308 3307 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13207 3310 3309 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13208 5183 3310 3309 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13209 3312 3311 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13210 5183 3312 3311 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13211 3314 3313 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13212 5183 3314 3313 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13213 3316 3315 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13214 5183 3316 3315 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13215 3318 3317 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13216 5183 3318 3317 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13217 3320 3319 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13218 5183 3320 3319 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13219 3322 3321 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13220 5183 3322 3321 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13221 3324 3323 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13222 5183 3324 3323 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13223 3326 3325 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13224 5183 3326 3325 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13225 3328 3327 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13226 5183 3328 3327 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13227 3330 3329 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13228 5183 3330 3329 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13229 3332 3331 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13230 5183 3332 3331 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13231 3334 3333 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13232 5183 3334 3333 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13233 3336 3335 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13234 5183 3336 3335 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13235 3338 3337 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13236 5183 3338 3337 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13237 3340 3339 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13238 5183 3340 3339 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13239 3342 3341 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13240 5183 3342 3341 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13241 3344 3343 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13242 5183 3344 3343 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13243 3346 3345 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13244 5183 3346 3345 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13245 3348 3347 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13246 5183 3348 3347 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13247 3350 3349 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13248 5183 3350 3349 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13249 3352 3351 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13250 5183 3352 3351 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13251 3354 3353 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13252 5183 3354 3353 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13253 3356 3355 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13254 5183 3356 3355 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13255 3358 3357 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13256 5183 3358 3357 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13257 3360 3359 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13258 5183 3360 3359 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13259 3362 3361 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13260 5183 3362 3361 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13261 3364 3363 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13262 5183 3364 3363 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13263 3366 3365 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13264 5183 3366 3365 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13265 3368 3367 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13266 5183 3368 3367 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13267 3370 3369 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13268 5183 3370 3369 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13269 3372 3371 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13270 5183 3372 3371 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13271 3374 3373 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13272 5183 3374 3373 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13273 3376 3375 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13274 5183 3376 3375 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13275 3378 3377 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13276 5183 3378 3377 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13277 3380 3379 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13278 5183 3380 3379 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13279 3382 3381 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13280 5183 3382 3381 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13281 3384 3383 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13282 5183 3384 3383 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13283 3386 3385 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13284 5183 3386 3385 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13285 3388 3387 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13286 5183 3388 3387 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13287 3390 3389 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13288 5183 3390 3389 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13289 3392 3391 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13290 5183 3392 3391 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13291 3394 3393 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13292 5183 3394 3393 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13293 3396 3395 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13294 5183 3396 3395 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13295 3398 3397 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13296 5183 3398 3397 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13297 3400 3399 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13298 5183 3400 3399 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13299 3402 3401 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13300 5183 3402 3401 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13301 3404 3403 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13302 5183 3404 3403 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13303 3406 3405 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13304 5183 3406 3405 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13305 3408 3407 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13306 5183 3408 3407 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13307 3410 3409 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13308 5183 3410 3409 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13309 3412 3411 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13310 5183 3412 3411 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13311 3414 3413 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13312 5183 3414 3413 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13313 3416 3415 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13314 5183 3416 3415 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13315 3418 3417 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13316 5183 3418 3417 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13317 3420 3419 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13318 5183 3420 3419 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13319 3422 3421 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13320 5183 3422 3421 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13321 3424 3423 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13322 5183 3424 3423 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13323 3426 3425 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13324 5183 3426 3425 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13325 3428 3427 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13326 5183 3428 3427 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13327 3430 3429 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13328 5183 3430 3429 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13329 3432 3431 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13330 5183 3432 3431 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13331 3434 3433 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13332 5183 3434 3433 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13333 3436 3435 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13334 5183 3436 3435 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13335 3438 3437 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13336 5183 3438 3437 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13337 3440 3439 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13338 5183 3440 3439 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13339 3442 3441 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13340 5183 3442 3441 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13341 3444 3443 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13342 5183 3444 3443 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13343 3446 3445 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13344 5183 3446 3445 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13345 3448 3447 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13346 5183 3448 3447 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13347 3450 3449 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13348 5183 3450 3449 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13349 3452 3451 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13350 5183 3452 3451 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13351 3454 3453 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13352 5183 3454 3453 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13353 3456 3455 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13354 5183 3456 3455 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13355 3458 3457 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13356 5183 3458 3457 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13357 3460 3459 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13358 5183 3460 3459 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13359 3462 3461 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13360 5183 3462 3461 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13361 3464 3463 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13362 5183 3464 3463 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13363 3466 3465 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13364 5183 3466 3465 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13365 3468 3467 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13366 5183 3468 3467 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13367 3470 3469 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13368 5183 3470 3469 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13369 3472 3471 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13370 5183 3472 3471 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13371 3474 3473 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13372 5183 3474 3473 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13373 3476 3475 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13374 5183 3476 3475 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13375 3478 3477 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13376 5183 3478 3477 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13377 3480 3479 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13378 5183 3480 3479 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13379 3482 3481 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13380 5183 3482 3481 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13381 3484 3483 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13382 5183 3484 3483 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13383 3486 3485 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13384 5183 3486 3485 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13385 3488 3487 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13386 5183 3488 3487 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13387 3490 3489 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13388 5183 3490 3489 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13389 3492 3491 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13390 5183 3492 3491 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13391 3494 3493 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13392 5183 3494 3493 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13393 3496 3495 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13394 5183 3496 3495 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13395 3498 3497 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13396 5183 3498 3497 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13397 3500 3499 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13398 5183 3500 3499 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13399 3502 3501 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13400 5183 3502 3501 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13401 3504 3503 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13402 5183 3504 3503 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13403 3506 3505 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13404 5183 3506 3505 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13405 3508 3507 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13406 5183 3508 3507 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13407 3510 3509 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13408 5183 3510 3509 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13409 3512 3511 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13410 5183 3512 3511 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13411 3514 3513 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13412 5183 3514 3513 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13413 3516 3515 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13414 5183 3516 3515 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13415 3518 3517 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13416 5183 3518 3517 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13417 3520 3519 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13418 5183 3520 3519 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13419 3522 3521 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13420 5183 3522 3521 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13421 3524 3523 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13422 5183 3524 3523 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13423 3526 3525 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13424 5183 3526 3525 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13425 3528 3527 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13426 5183 3528 3527 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13427 3530 3529 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13428 5183 3530 3529 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13429 3532 3531 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13430 5183 3532 3531 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13431 3534 3533 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13432 5183 3534 3533 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13433 3536 3535 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13434 5183 3536 3535 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13435 3538 3537 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13436 5183 3538 3537 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13437 3540 3539 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13438 5183 3540 3539 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13439 3542 3541 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13440 5183 3542 3541 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13441 3544 3543 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13442 5183 3544 3543 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13443 3546 3545 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13444 5183 3546 3545 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13445 3548 3547 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13446 5183 3548 3547 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13447 3550 3549 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13448 5183 3550 3549 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13449 3552 3551 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13450 5183 3552 3551 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13451 3554 3553 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13452 5183 3554 3553 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13453 3556 3555 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13454 5183 3556 3555 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13455 3558 3557 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13456 5183 3558 3557 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13457 3560 3559 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13458 5183 3560 3559 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13459 3562 3561 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13460 5183 3562 3561 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13461 3564 3563 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13462 5183 3564 3563 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13463 3566 3565 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13464 5183 3566 3565 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13465 3568 3567 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13466 5183 3568 3567 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13467 3570 3569 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13468 5183 3570 3569 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13469 3572 3571 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13470 5183 3572 3571 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13471 3574 3573 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13472 5183 3574 3573 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13473 3576 3575 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13474 5183 3576 3575 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13475 3578 3577 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13476 5183 3578 3577 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13477 3580 3579 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13478 5183 3580 3579 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13479 3582 3581 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13480 5183 3582 3581 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13481 3584 3583 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13482 5183 3584 3583 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13483 3586 3585 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13484 5183 3586 3585 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13485 3588 3587 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13486 5183 3588 3587 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13487 3590 3589 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13488 5183 3590 3589 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13489 3592 3591 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13490 5183 3592 3591 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13491 3594 3593 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13492 5183 3594 3593 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13493 3596 3595 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13494 5183 3596 3595 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13495 3598 3597 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13496 5183 3598 3597 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13497 3607 3599 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_13498 5183 3599 3599 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_13499 3601 3601 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_13500 5183 3601 3600 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_13501 3602 3603 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_13502 5183 3603 3603 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_13503 3604 5188 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_13504 5183 3606 3605 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_13505 3606 5188 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_13506 5183 5188 3606 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_13507 5188 3609 5183 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_13508 5183 3609 5188 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_13509 5183 5176 3609 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_13510 3609 3607 5183 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_13511 3609 5179 3608 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_13512 3611 3610 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13513 5183 3611 3610 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13514 3613 3612 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13515 5183 3613 3612 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13516 3615 3614 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13517 5183 3615 3614 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13518 3617 3616 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13519 5183 3617 3616 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13520 3619 3618 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13521 5183 3619 3618 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13522 3621 3620 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13523 5183 3621 3620 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13524 3623 3622 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13525 5183 3623 3622 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13526 3625 3624 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13527 5183 3625 3624 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13528 3627 3626 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13529 5183 3627 3626 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13530 3629 3628 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13531 5183 3629 3628 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13532 3631 3630 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13533 5183 3631 3630 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13534 3633 3632 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13535 5183 3633 3632 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13536 3635 3634 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13537 5183 3635 3634 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13538 3637 3636 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13539 5183 3637 3636 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13540 3639 3638 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13541 5183 3639 3638 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13542 3641 3640 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13543 5183 3641 3640 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13544 3643 3642 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13545 5183 3643 3642 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13546 3645 3644 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13547 5183 3645 3644 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13548 3647 3646 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13549 5183 3647 3646 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13550 3649 3648 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13551 5183 3649 3648 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13552 3651 3650 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13553 5183 3651 3650 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13554 3653 3652 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13555 5183 3653 3652 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13556 3655 3654 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13557 5183 3655 3654 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13558 3657 3656 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13559 5183 3657 3656 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13560 3659 3658 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13561 5183 3659 3658 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13562 3661 3660 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13563 5183 3661 3660 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13564 3663 3662 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13565 5183 3663 3662 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13566 3665 3664 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13567 5183 3665 3664 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13568 3667 3666 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13569 5183 3667 3666 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13570 3669 3668 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13571 5183 3669 3668 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13572 3671 3670 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13573 5183 3671 3670 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13574 3673 3672 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13575 5183 3673 3672 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13576 3675 3674 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13577 5183 3675 3674 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13578 3677 3676 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13579 5183 3677 3676 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13580 3679 3678 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13581 5183 3679 3678 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13582 3681 3680 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13583 5183 3681 3680 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13584 3683 3682 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13585 5183 3683 3682 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13586 3685 3684 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13587 5183 3685 3684 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13588 3687 3686 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13589 5183 3687 3686 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13590 3689 3688 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13591 5183 3689 3688 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13592 3691 3690 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13593 5183 3691 3690 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13594 3693 3692 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13595 5183 3693 3692 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13596 3695 3694 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13597 5183 3695 3694 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13598 3697 3696 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13599 5183 3697 3696 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13600 3699 3698 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13601 5183 3699 3698 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13602 3701 3700 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13603 5183 3701 3700 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13604 3703 3702 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13605 5183 3703 3702 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13606 3705 3704 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13607 5183 3705 3704 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13608 3707 3706 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13609 5183 3707 3706 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13610 3709 3708 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13611 5183 3709 3708 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13612 3711 3710 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13613 5183 3711 3710 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13614 3713 3712 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13615 5183 3713 3712 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13616 3715 3714 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13617 5183 3715 3714 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13618 3717 3716 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13619 5183 3717 3716 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13620 3719 3718 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13621 5183 3719 3718 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13622 3721 3720 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13623 5183 3721 3720 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13624 3723 3722 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13625 5183 3723 3722 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13626 3725 3724 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13627 5183 3725 3724 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13628 3727 3726 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13629 5183 3727 3726 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13630 3729 3728 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13631 5183 3729 3728 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13632 3731 3730 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13633 5183 3731 3730 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13634 3733 3732 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13635 5183 3733 3732 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13636 3735 3734 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13637 5183 3735 3734 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13638 3737 3736 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13639 5183 3737 3736 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13640 3739 3738 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13641 5183 3739 3738 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13642 3741 3740 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13643 5183 3741 3740 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13644 3743 3742 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13645 5183 3743 3742 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13646 3745 3744 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13647 5183 3745 3744 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13648 3747 3746 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13649 5183 3747 3746 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13650 3749 3748 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13651 5183 3749 3748 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13652 3751 3750 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13653 5183 3751 3750 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13654 3753 3752 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13655 5183 3753 3752 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13656 3755 3754 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13657 5183 3755 3754 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13658 3757 3756 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13659 5183 3757 3756 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13660 3759 3758 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13661 5183 3759 3758 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13662 3761 3760 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13663 5183 3761 3760 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13664 3763 3762 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13665 5183 3763 3762 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13666 3765 3764 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13667 5183 3765 3764 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13668 3767 3766 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13669 5183 3767 3766 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13670 3769 3768 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13671 5183 3769 3768 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13672 3771 3770 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13673 5183 3771 3770 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13674 3773 3772 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13675 5183 3773 3772 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13676 3775 3774 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13677 5183 3775 3774 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13678 3777 3776 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13679 5183 3777 3776 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13680 3779 3778 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13681 5183 3779 3778 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13682 3781 3780 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13683 5183 3781 3780 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13684 3783 3782 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13685 5183 3783 3782 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13686 3785 3784 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13687 5183 3785 3784 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13688 3787 3786 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13689 5183 3787 3786 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13690 3789 3788 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13691 5183 3789 3788 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13692 3791 3790 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13693 5183 3791 3790 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13694 3793 3792 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13695 5183 3793 3792 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13696 3795 3794 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13697 5183 3795 3794 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13698 3797 3796 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13699 5183 3797 3796 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13700 3799 3798 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13701 5183 3799 3798 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13702 3801 3800 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13703 5183 3801 3800 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13704 3803 3802 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13705 5183 3803 3802 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13706 3805 3804 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13707 5183 3805 3804 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13708 3807 3806 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13709 5183 3807 3806 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13710 3809 3808 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13711 5183 3809 3808 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13712 3811 3810 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13713 5183 3811 3810 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13714 3813 3812 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13715 5183 3813 3812 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13716 3815 3814 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13717 5183 3815 3814 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13718 3817 3816 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13719 5183 3817 3816 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13720 3819 3818 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13721 5183 3819 3818 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13722 3821 3820 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13723 5183 3821 3820 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13724 3823 3822 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13725 5183 3823 3822 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13726 3825 3824 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13727 5183 3825 3824 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13728 3827 3826 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13729 5183 3827 3826 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13730 3829 3828 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13731 5183 3829 3828 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13732 3831 3830 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13733 5183 3831 3830 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13734 3833 3832 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13735 5183 3833 3832 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13736 3835 3834 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13737 5183 3835 3834 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13738 3837 3836 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13739 5183 3837 3836 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13740 3839 3838 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13741 5183 3839 3838 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13742 3841 3840 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13743 5183 3841 3840 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13744 3843 3842 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13745 5183 3843 3842 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13746 3845 3844 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13747 5183 3845 3844 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13748 3847 3846 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13749 5183 3847 3846 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13750 3849 3848 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13751 5183 3849 3848 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13752 3851 3850 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13753 5183 3851 3850 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13754 3853 3852 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13755 5183 3853 3852 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13756 3855 3854 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13757 5183 3855 3854 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13758 3857 3856 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13759 5183 3857 3856 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13760 3859 3858 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13761 5183 3859 3858 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13762 3861 3860 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13763 5183 3861 3860 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13764 3863 3862 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13765 5183 3863 3862 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13766 3865 3864 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13767 5183 3865 3864 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13768 3867 3866 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13769 5183 3867 3866 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13770 3869 3868 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13771 5183 3869 3868 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13772 3871 3870 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13773 5183 3871 3870 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13774 3873 3872 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13775 5183 3873 3872 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13776 3875 3874 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13777 5183 3875 3874 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13778 3877 3876 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13779 5183 3877 3876 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13780 3879 3878 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13781 5183 3879 3878 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13782 3881 3880 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13783 5183 3881 3880 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13784 3883 3882 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13785 5183 3883 3882 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13786 3885 3884 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13787 5183 3885 3884 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13788 3887 3886 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13789 5183 3887 3886 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13790 3889 3888 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13791 5183 3889 3888 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13792 3891 3890 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13793 5183 3891 3890 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13794 3893 3892 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13795 5183 3893 3892 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13796 3895 3894 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13797 5183 3895 3894 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13798 3897 3896 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13799 5183 3897 3896 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13800 3899 3898 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13801 5183 3899 3898 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13802 3901 3900 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13803 5183 3901 3900 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13804 3903 3902 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13805 5183 3903 3902 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13806 3905 3904 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13807 5183 3905 3904 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13808 3907 3906 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13809 5183 3907 3906 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13810 3909 3908 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13811 5183 3909 3908 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13812 3911 3910 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13813 5183 3911 3910 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13814 3913 3912 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13815 5183 3913 3912 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13816 3915 3914 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13817 5183 3915 3914 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13818 3917 3916 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13819 5183 3917 3916 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13820 3919 3918 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13821 5183 3919 3918 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13822 3921 3920 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13823 5183 3921 3920 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13824 3923 3922 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13825 5183 3923 3922 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13826 3925 3924 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13827 5183 3925 3924 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13828 3927 3926 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13829 5183 3927 3926 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13830 3929 3928 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13831 5183 3929 3928 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13832 3931 3930 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13833 5183 3931 3930 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13834 3933 3932 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13835 5183 3933 3932 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13836 3935 3934 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13837 5183 3935 3934 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13838 3937 3936 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13839 5183 3937 3936 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13840 3939 3938 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13841 5183 3939 3938 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13842 3941 3940 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13843 5183 3941 3940 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13844 3943 3942 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13845 5183 3943 3942 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13846 3945 3944 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13847 5183 3945 3944 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13848 3947 3946 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13849 5183 3947 3946 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13850 3949 3948 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13851 5183 3949 3948 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13852 3951 3950 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13853 5183 3951 3950 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13854 3953 3952 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13855 5183 3953 3952 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13856 3955 3954 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13857 5183 3955 3954 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13858 3957 3956 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13859 5183 3957 3956 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13860 3959 3958 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13861 5183 3959 3958 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13862 3961 3960 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13863 5183 3961 3960 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13864 3963 3962 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13865 5183 3963 3962 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13866 3965 3964 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13867 5183 3965 3964 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13868 3967 3966 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13869 5183 3967 3966 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13870 3969 3968 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13871 5183 3969 3968 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13872 3971 3970 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13873 5183 3971 3970 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13874 3973 3972 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13875 5183 3973 3972 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13876 3975 3974 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13877 5183 3975 3974 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13878 3977 3976 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13879 5183 3977 3976 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13880 3979 3978 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13881 5183 3979 3978 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13882 3981 3980 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13883 5183 3981 3980 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13884 3983 3982 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13885 5183 3983 3982 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13886 3985 3984 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13887 5183 3985 3984 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13888 3987 3986 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13889 5183 3987 3986 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13890 3989 3988 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13891 5183 3989 3988 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13892 3991 3990 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13893 5183 3991 3990 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13894 3993 3992 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13895 5183 3993 3992 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13896 3995 3994 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13897 5183 3995 3994 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13898 3997 3996 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13899 5183 3997 3996 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13900 3999 3998 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13901 5183 3999 3998 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13902 4001 4000 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13903 5183 4001 4000 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13904 4003 4002 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13905 5183 4003 4002 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13906 4005 4004 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13907 5183 4005 4004 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13908 4007 4006 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13909 5183 4007 4006 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13910 4009 4008 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13911 5183 4009 4008 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13912 4011 4010 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13913 5183 4011 4010 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13914 4013 4012 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13915 5183 4013 4012 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13916 4015 4014 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13917 5183 4015 4014 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13918 4017 4016 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13919 5183 4017 4016 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13920 4019 4018 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13921 5183 4019 4018 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13922 4021 4020 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13923 5183 4021 4020 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13924 4023 4022 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13925 5183 4023 4022 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13926 4025 4024 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13927 5183 4025 4024 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13928 4027 4026 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13929 5183 4027 4026 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13930 4029 4028 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13931 5183 4029 4028 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13932 4031 4030 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13933 5183 4031 4030 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13934 4033 4032 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13935 5183 4033 4032 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13936 4035 4034 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13937 5183 4035 4034 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13938 4037 4036 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13939 5183 4037 4036 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13940 4039 4038 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13941 5183 4039 4038 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13942 4041 4040 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13943 5183 4041 4040 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13944 4043 4042 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13945 5183 4043 4042 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13946 4045 4044 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13947 5183 4045 4044 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13948 4047 4046 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13949 5183 4047 4046 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13950 4049 4048 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13951 5183 4049 4048 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13952 4051 4050 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13953 5183 4051 4050 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13954 4053 4052 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13955 5183 4053 4052 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13956 4055 4054 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13957 5183 4055 4054 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13958 4057 4056 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13959 5183 4057 4056 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13960 4059 4058 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13961 5183 4059 4058 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13962 4061 4060 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13963 5183 4061 4060 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13964 4063 4062 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13965 5183 4063 4062 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13966 4065 4064 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13967 5183 4065 4064 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13968 4067 4066 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13969 5183 4067 4066 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13970 4069 4068 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13971 5183 4069 4068 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13972 4071 4070 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13973 5183 4071 4070 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13974 4073 4072 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13975 5183 4073 4072 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13976 4075 4074 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13977 5183 4075 4074 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13978 4077 4076 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13979 5183 4077 4076 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13980 4079 4078 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13981 5183 4079 4078 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13982 4081 4080 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13983 5183 4081 4080 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13984 4083 4082 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13985 5183 4083 4082 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13986 4085 4084 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13987 5183 4085 4084 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13988 4087 4086 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13989 5183 4087 4086 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13990 4089 4088 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13991 5183 4089 4088 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13992 4091 4090 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13993 5183 4091 4090 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13994 4093 4092 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13995 5183 4093 4092 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13996 4095 4094 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13997 5183 4095 4094 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13998 4097 4096 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_13999 5183 4097 4096 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14000 4099 4098 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14001 5183 4099 4098 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14002 4101 4100 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14003 5183 4101 4100 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14004 4103 4102 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14005 5183 4103 4102 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14006 4105 4104 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14007 5183 4105 4104 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14008 4107 4106 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14009 5183 4107 4106 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14010 4109 4108 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14011 5183 4109 4108 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14012 4111 4110 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14013 5183 4111 4110 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14014 4113 4112 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14015 5183 4113 4112 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14016 4115 4114 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14017 5183 4115 4114 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14018 4117 4116 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14019 5183 4117 4116 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14020 4119 4118 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14021 5183 4119 4118 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14022 4121 4120 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14023 5183 4121 4120 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14024 4130 4122 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14025 5183 4122 4122 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14026 4124 4124 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14027 5183 4124 4123 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14028 4125 4126 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14029 5183 4126 4126 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14030 4127 5187 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14031 5183 4129 4128 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14032 4129 5187 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14033 5183 5187 4129 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14034 5187 4132 5183 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_14035 5183 4132 5187 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_14036 5183 5176 4132 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_14037 4132 4130 5183 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_14038 4132 5179 4131 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_14039 4134 4133 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14040 5183 4134 4133 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14041 4136 4135 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14042 5183 4136 4135 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14043 4138 4137 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14044 5183 4138 4137 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14045 4140 4139 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14046 5183 4140 4139 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14047 4142 4141 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14048 5183 4142 4141 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14049 4144 4143 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14050 5183 4144 4143 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14051 4146 4145 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14052 5183 4146 4145 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14053 4148 4147 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14054 5183 4148 4147 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14055 4150 4149 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14056 5183 4150 4149 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14057 4152 4151 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14058 5183 4152 4151 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14059 4154 4153 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14060 5183 4154 4153 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14061 4156 4155 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14062 5183 4156 4155 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14063 4158 4157 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14064 5183 4158 4157 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14065 4160 4159 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14066 5183 4160 4159 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14067 4162 4161 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14068 5183 4162 4161 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14069 4164 4163 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14070 5183 4164 4163 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14071 4166 4165 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14072 5183 4166 4165 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14073 4168 4167 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14074 5183 4168 4167 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14075 4170 4169 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14076 5183 4170 4169 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14077 4172 4171 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14078 5183 4172 4171 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14079 4174 4173 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14080 5183 4174 4173 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14081 4176 4175 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14082 5183 4176 4175 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14083 4178 4177 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14084 5183 4178 4177 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14085 4180 4179 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14086 5183 4180 4179 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14087 4182 4181 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14088 5183 4182 4181 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14089 4184 4183 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14090 5183 4184 4183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14091 4186 4185 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14092 5183 4186 4185 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14093 4188 4187 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14094 5183 4188 4187 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14095 4190 4189 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14096 5183 4190 4189 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14097 4192 4191 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14098 5183 4192 4191 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14099 4194 4193 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14100 5183 4194 4193 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14101 4196 4195 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14102 5183 4196 4195 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14103 4198 4197 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14104 5183 4198 4197 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14105 4200 4199 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14106 5183 4200 4199 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14107 4202 4201 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14108 5183 4202 4201 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14109 4204 4203 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14110 5183 4204 4203 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14111 4206 4205 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14112 5183 4206 4205 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14113 4208 4207 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14114 5183 4208 4207 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14115 4210 4209 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14116 5183 4210 4209 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14117 4212 4211 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14118 5183 4212 4211 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14119 4214 4213 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14120 5183 4214 4213 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14121 4216 4215 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14122 5183 4216 4215 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14123 4218 4217 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14124 5183 4218 4217 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14125 4220 4219 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14126 5183 4220 4219 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14127 4222 4221 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14128 5183 4222 4221 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14129 4224 4223 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14130 5183 4224 4223 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14131 4226 4225 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14132 5183 4226 4225 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14133 4228 4227 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14134 5183 4228 4227 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14135 4230 4229 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14136 5183 4230 4229 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14137 4232 4231 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14138 5183 4232 4231 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14139 4234 4233 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14140 5183 4234 4233 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14141 4236 4235 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14142 5183 4236 4235 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14143 4238 4237 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14144 5183 4238 4237 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14145 4240 4239 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14146 5183 4240 4239 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14147 4242 4241 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14148 5183 4242 4241 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14149 4244 4243 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14150 5183 4244 4243 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14151 4246 4245 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14152 5183 4246 4245 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14153 4248 4247 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14154 5183 4248 4247 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14155 4250 4249 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14156 5183 4250 4249 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14157 4252 4251 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14158 5183 4252 4251 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14159 4254 4253 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14160 5183 4254 4253 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14161 4256 4255 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14162 5183 4256 4255 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14163 4258 4257 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14164 5183 4258 4257 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14165 4260 4259 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14166 5183 4260 4259 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14167 4262 4261 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14168 5183 4262 4261 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14169 4264 4263 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14170 5183 4264 4263 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14171 4266 4265 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14172 5183 4266 4265 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14173 4268 4267 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14174 5183 4268 4267 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14175 4270 4269 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14176 5183 4270 4269 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14177 4272 4271 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14178 5183 4272 4271 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14179 4274 4273 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14180 5183 4274 4273 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14181 4276 4275 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14182 5183 4276 4275 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14183 4278 4277 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14184 5183 4278 4277 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14185 4280 4279 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14186 5183 4280 4279 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14187 4282 4281 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14188 5183 4282 4281 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14189 4284 4283 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14190 5183 4284 4283 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14191 4286 4285 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14192 5183 4286 4285 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14193 4288 4287 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14194 5183 4288 4287 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14195 4290 4289 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14196 5183 4290 4289 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14197 4292 4291 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14198 5183 4292 4291 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14199 4294 4293 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14200 5183 4294 4293 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14201 4296 4295 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14202 5183 4296 4295 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14203 4298 4297 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14204 5183 4298 4297 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14205 4300 4299 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14206 5183 4300 4299 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14207 4302 4301 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14208 5183 4302 4301 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14209 4304 4303 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14210 5183 4304 4303 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14211 4306 4305 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14212 5183 4306 4305 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14213 4308 4307 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14214 5183 4308 4307 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14215 4310 4309 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14216 5183 4310 4309 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14217 4312 4311 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14218 5183 4312 4311 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14219 4314 4313 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14220 5183 4314 4313 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14221 4316 4315 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14222 5183 4316 4315 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14223 4318 4317 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14224 5183 4318 4317 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14225 4320 4319 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14226 5183 4320 4319 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14227 4322 4321 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14228 5183 4322 4321 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14229 4324 4323 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14230 5183 4324 4323 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14231 4326 4325 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14232 5183 4326 4325 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14233 4328 4327 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14234 5183 4328 4327 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14235 4330 4329 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14236 5183 4330 4329 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14237 4332 4331 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14238 5183 4332 4331 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14239 4334 4333 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14240 5183 4334 4333 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14241 4336 4335 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14242 5183 4336 4335 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14243 4338 4337 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14244 5183 4338 4337 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14245 4340 4339 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14246 5183 4340 4339 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14247 4342 4341 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14248 5183 4342 4341 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14249 4344 4343 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14250 5183 4344 4343 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14251 4346 4345 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14252 5183 4346 4345 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14253 4348 4347 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14254 5183 4348 4347 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14255 4350 4349 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14256 5183 4350 4349 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14257 4352 4351 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14258 5183 4352 4351 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14259 4354 4353 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14260 5183 4354 4353 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14261 4356 4355 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14262 5183 4356 4355 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14263 4358 4357 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14264 5183 4358 4357 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14265 4360 4359 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14266 5183 4360 4359 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14267 4362 4361 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14268 5183 4362 4361 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14269 4364 4363 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14270 5183 4364 4363 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14271 4366 4365 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14272 5183 4366 4365 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14273 4368 4367 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14274 5183 4368 4367 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14275 4370 4369 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14276 5183 4370 4369 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14277 4372 4371 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14278 5183 4372 4371 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14279 4374 4373 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14280 5183 4374 4373 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14281 4376 4375 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14282 5183 4376 4375 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14283 4378 4377 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14284 5183 4378 4377 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14285 4380 4379 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14286 5183 4380 4379 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14287 4382 4381 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14288 5183 4382 4381 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14289 4384 4383 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14290 5183 4384 4383 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14291 4386 4385 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14292 5183 4386 4385 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14293 4388 4387 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14294 5183 4388 4387 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14295 4390 4389 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14296 5183 4390 4389 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14297 4392 4391 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14298 5183 4392 4391 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14299 4394 4393 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14300 5183 4394 4393 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14301 4396 4395 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14302 5183 4396 4395 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14303 4398 4397 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14304 5183 4398 4397 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14305 4400 4399 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14306 5183 4400 4399 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14307 4402 4401 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14308 5183 4402 4401 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14309 4404 4403 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14310 5183 4404 4403 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14311 4406 4405 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14312 5183 4406 4405 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14313 4408 4407 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14314 5183 4408 4407 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14315 4410 4409 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14316 5183 4410 4409 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14317 4412 4411 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14318 5183 4412 4411 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14319 4414 4413 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14320 5183 4414 4413 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14321 4416 4415 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14322 5183 4416 4415 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14323 4418 4417 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14324 5183 4418 4417 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14325 4420 4419 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14326 5183 4420 4419 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14327 4422 4421 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14328 5183 4422 4421 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14329 4424 4423 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14330 5183 4424 4423 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14331 4426 4425 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14332 5183 4426 4425 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14333 4428 4427 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14334 5183 4428 4427 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14335 4430 4429 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14336 5183 4430 4429 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14337 4432 4431 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14338 5183 4432 4431 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14339 4434 4433 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14340 5183 4434 4433 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14341 4436 4435 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14342 5183 4436 4435 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14343 4438 4437 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14344 5183 4438 4437 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14345 4440 4439 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14346 5183 4440 4439 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14347 4442 4441 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14348 5183 4442 4441 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14349 4444 4443 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14350 5183 4444 4443 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14351 4446 4445 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14352 5183 4446 4445 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14353 4448 4447 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14354 5183 4448 4447 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14355 4450 4449 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14356 5183 4450 4449 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14357 4452 4451 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14358 5183 4452 4451 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14359 4454 4453 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14360 5183 4454 4453 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14361 4456 4455 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14362 5183 4456 4455 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14363 4458 4457 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14364 5183 4458 4457 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14365 4460 4459 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14366 5183 4460 4459 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14367 4462 4461 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14368 5183 4462 4461 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14369 4464 4463 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14370 5183 4464 4463 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14371 4466 4465 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14372 5183 4466 4465 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14373 4468 4467 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14374 5183 4468 4467 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14375 4470 4469 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14376 5183 4470 4469 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14377 4472 4471 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14378 5183 4472 4471 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14379 4474 4473 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14380 5183 4474 4473 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14381 4476 4475 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14382 5183 4476 4475 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14383 4478 4477 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14384 5183 4478 4477 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14385 4480 4479 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14386 5183 4480 4479 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14387 4482 4481 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14388 5183 4482 4481 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14389 4484 4483 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14390 5183 4484 4483 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14391 4486 4485 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14392 5183 4486 4485 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14393 4488 4487 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14394 5183 4488 4487 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14395 4490 4489 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14396 5183 4490 4489 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14397 4492 4491 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14398 5183 4492 4491 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14399 4494 4493 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14400 5183 4494 4493 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14401 4496 4495 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14402 5183 4496 4495 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14403 4498 4497 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14404 5183 4498 4497 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14405 4500 4499 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14406 5183 4500 4499 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14407 4502 4501 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14408 5183 4502 4501 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14409 4504 4503 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14410 5183 4504 4503 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14411 4506 4505 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14412 5183 4506 4505 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14413 4508 4507 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14414 5183 4508 4507 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14415 4510 4509 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14416 5183 4510 4509 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14417 4512 4511 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14418 5183 4512 4511 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14419 4514 4513 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14420 5183 4514 4513 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14421 4516 4515 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14422 5183 4516 4515 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14423 4518 4517 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14424 5183 4518 4517 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14425 4520 4519 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14426 5183 4520 4519 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14427 4522 4521 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14428 5183 4522 4521 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14429 4524 4523 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14430 5183 4524 4523 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14431 4526 4525 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14432 5183 4526 4525 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14433 4528 4527 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14434 5183 4528 4527 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14435 4530 4529 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14436 5183 4530 4529 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14437 4532 4531 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14438 5183 4532 4531 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14439 4534 4533 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14440 5183 4534 4533 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14441 4536 4535 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14442 5183 4536 4535 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14443 4538 4537 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14444 5183 4538 4537 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14445 4540 4539 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14446 5183 4540 4539 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14447 4542 4541 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14448 5183 4542 4541 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14449 4544 4543 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14450 5183 4544 4543 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14451 4546 4545 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14452 5183 4546 4545 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14453 4548 4547 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14454 5183 4548 4547 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14455 4550 4549 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14456 5183 4550 4549 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14457 4552 4551 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14458 5183 4552 4551 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14459 4554 4553 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14460 5183 4554 4553 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14461 4556 4555 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14462 5183 4556 4555 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14463 4558 4557 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14464 5183 4558 4557 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14465 4560 4559 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14466 5183 4560 4559 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14467 4562 4561 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14468 5183 4562 4561 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14469 4564 4563 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14470 5183 4564 4563 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14471 4566 4565 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14472 5183 4566 4565 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14473 4568 4567 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14474 5183 4568 4567 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14475 4570 4569 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14476 5183 4570 4569 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14477 4572 4571 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14478 5183 4572 4571 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14479 4574 4573 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14480 5183 4574 4573 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14481 4576 4575 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14482 5183 4576 4575 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14483 4578 4577 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14484 5183 4578 4577 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14485 4580 4579 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14486 5183 4580 4579 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14487 4582 4581 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14488 5183 4582 4581 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14489 4584 4583 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14490 5183 4584 4583 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14491 4586 4585 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14492 5183 4586 4585 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14493 4588 4587 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14494 5183 4588 4587 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14495 4590 4589 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14496 5183 4590 4589 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14497 4592 4591 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14498 5183 4592 4591 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14499 4594 4593 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14500 5183 4594 4593 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14501 4596 4595 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14502 5183 4596 4595 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14503 4598 4597 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14504 5183 4598 4597 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14505 4600 4599 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14506 5183 4600 4599 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14507 4602 4601 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14508 5183 4602 4601 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14509 4604 4603 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14510 5183 4604 4603 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14511 4606 4605 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14512 5183 4606 4605 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14513 4608 4607 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14514 5183 4608 4607 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14515 4610 4609 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14516 5183 4610 4609 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14517 4612 4611 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14518 5183 4612 4611 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14519 4614 4613 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14520 5183 4614 4613 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14521 4616 4615 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14522 5183 4616 4615 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14523 4618 4617 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14524 5183 4618 4617 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14525 4620 4619 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14526 5183 4620 4619 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14527 4622 4621 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14528 5183 4622 4621 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14529 4624 4623 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14530 5183 4624 4623 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14531 4626 4625 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14532 5183 4626 4625 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14533 4628 4627 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14534 5183 4628 4627 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14535 4630 4629 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14536 5183 4630 4629 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14537 4632 4631 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14538 5183 4632 4631 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14539 4634 4633 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14540 5183 4634 4633 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14541 4636 4635 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14542 5183 4636 4635 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14543 4638 4637 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14544 5183 4638 4637 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14545 4640 4639 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14546 5183 4640 4639 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14547 4642 4641 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14548 5183 4642 4641 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14549 4644 4643 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14550 5183 4644 4643 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14551 4653 4645 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14552 5183 4645 4645 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14553 4647 4647 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14554 5183 4647 4646 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14555 4648 4649 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14556 5183 4649 4649 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14557 4650 5186 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14558 5183 4652 4651 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14559 4652 5186 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14560 5183 5186 4652 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_14561 5186 4655 5183 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_14562 5183 4655 5186 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_14563 5183 5176 4655 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_14564 4655 4653 5183 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_14565 4655 5179 4654 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_14566 4657 4656 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14567 5183 4657 4656 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14568 4659 4658 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14569 5183 4659 4658 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14570 4661 4660 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14571 5183 4661 4660 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14572 4663 4662 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14573 5183 4663 4662 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14574 4665 4664 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14575 5183 4665 4664 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14576 4667 4666 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14577 5183 4667 4666 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14578 4669 4668 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14579 5183 4669 4668 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14580 4671 4670 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14581 5183 4671 4670 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14582 4673 4672 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14583 5183 4673 4672 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14584 4675 4674 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14585 5183 4675 4674 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14586 4677 4676 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14587 5183 4677 4676 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14588 4679 4678 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14589 5183 4679 4678 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14590 4681 4680 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14591 5183 4681 4680 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14592 4683 4682 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14593 5183 4683 4682 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14594 4685 4684 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14595 5183 4685 4684 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14596 4687 4686 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14597 5183 4687 4686 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14598 4689 4688 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14599 5183 4689 4688 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14600 4691 4690 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14601 5183 4691 4690 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14602 4693 4692 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14603 5183 4693 4692 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14604 4695 4694 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14605 5183 4695 4694 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14606 4697 4696 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14607 5183 4697 4696 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14608 4699 4698 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14609 5183 4699 4698 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14610 4701 4700 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14611 5183 4701 4700 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14612 4703 4702 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14613 5183 4703 4702 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14614 4705 4704 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14615 5183 4705 4704 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14616 4707 4706 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14617 5183 4707 4706 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14618 4709 4708 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14619 5183 4709 4708 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14620 4711 4710 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14621 5183 4711 4710 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14622 4713 4712 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14623 5183 4713 4712 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14624 4715 4714 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14625 5183 4715 4714 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14626 4717 4716 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14627 5183 4717 4716 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14628 4719 4718 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14629 5183 4719 4718 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14630 4721 4720 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14631 5183 4721 4720 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14632 4723 4722 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14633 5183 4723 4722 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14634 4725 4724 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14635 5183 4725 4724 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14636 4727 4726 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14637 5183 4727 4726 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14638 4729 4728 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14639 5183 4729 4728 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14640 4731 4730 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14641 5183 4731 4730 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14642 4733 4732 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14643 5183 4733 4732 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14644 4735 4734 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14645 5183 4735 4734 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14646 4737 4736 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14647 5183 4737 4736 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14648 4739 4738 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14649 5183 4739 4738 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14650 4741 4740 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14651 5183 4741 4740 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14652 4743 4742 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14653 5183 4743 4742 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14654 4745 4744 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14655 5183 4745 4744 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14656 4747 4746 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14657 5183 4747 4746 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14658 4749 4748 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14659 5183 4749 4748 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14660 4751 4750 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14661 5183 4751 4750 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14662 4753 4752 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14663 5183 4753 4752 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14664 4755 4754 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14665 5183 4755 4754 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14666 4757 4756 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14667 5183 4757 4756 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14668 4759 4758 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14669 5183 4759 4758 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14670 4761 4760 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14671 5183 4761 4760 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14672 4763 4762 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14673 5183 4763 4762 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14674 4765 4764 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14675 5183 4765 4764 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14676 4767 4766 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14677 5183 4767 4766 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14678 4769 4768 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14679 5183 4769 4768 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14680 4771 4770 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14681 5183 4771 4770 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14682 4773 4772 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14683 5183 4773 4772 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14684 4775 4774 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14685 5183 4775 4774 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14686 4777 4776 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14687 5183 4777 4776 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14688 4779 4778 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14689 5183 4779 4778 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14690 4781 4780 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14691 5183 4781 4780 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14692 4783 4782 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14693 5183 4783 4782 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14694 4785 4784 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14695 5183 4785 4784 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14696 4787 4786 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14697 5183 4787 4786 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14698 4789 4788 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14699 5183 4789 4788 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14700 4791 4790 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14701 5183 4791 4790 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14702 4793 4792 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14703 5183 4793 4792 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14704 4795 4794 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14705 5183 4795 4794 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14706 4797 4796 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14707 5183 4797 4796 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14708 4799 4798 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14709 5183 4799 4798 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14710 4801 4800 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14711 5183 4801 4800 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14712 4803 4802 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14713 5183 4803 4802 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14714 4805 4804 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14715 5183 4805 4804 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14716 4807 4806 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14717 5183 4807 4806 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14718 4809 4808 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14719 5183 4809 4808 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14720 4811 4810 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14721 5183 4811 4810 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14722 4813 4812 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14723 5183 4813 4812 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14724 4815 4814 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14725 5183 4815 4814 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14726 4817 4816 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14727 5183 4817 4816 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14728 4819 4818 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14729 5183 4819 4818 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14730 4821 4820 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14731 5183 4821 4820 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14732 4823 4822 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14733 5183 4823 4822 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14734 4825 4824 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14735 5183 4825 4824 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14736 4827 4826 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14737 5183 4827 4826 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14738 4829 4828 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14739 5183 4829 4828 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14740 4831 4830 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14741 5183 4831 4830 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14742 4833 4832 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14743 5183 4833 4832 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14744 4835 4834 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14745 5183 4835 4834 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14746 4837 4836 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14747 5183 4837 4836 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14748 4839 4838 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14749 5183 4839 4838 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14750 4841 4840 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14751 5183 4841 4840 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14752 4843 4842 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14753 5183 4843 4842 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14754 4845 4844 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14755 5183 4845 4844 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14756 4847 4846 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14757 5183 4847 4846 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14758 4849 4848 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14759 5183 4849 4848 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14760 4851 4850 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14761 5183 4851 4850 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14762 4853 4852 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14763 5183 4853 4852 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14764 4855 4854 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14765 5183 4855 4854 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14766 4857 4856 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14767 5183 4857 4856 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14768 4859 4858 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14769 5183 4859 4858 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14770 4861 4860 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14771 5183 4861 4860 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14772 4863 4862 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14773 5183 4863 4862 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14774 4865 4864 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14775 5183 4865 4864 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14776 4867 4866 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14777 5183 4867 4866 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14778 4869 4868 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14779 5183 4869 4868 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14780 4871 4870 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14781 5183 4871 4870 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14782 4873 4872 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14783 5183 4873 4872 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14784 4875 4874 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14785 5183 4875 4874 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14786 4877 4876 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14787 5183 4877 4876 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14788 4879 4878 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14789 5183 4879 4878 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14790 4881 4880 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14791 5183 4881 4880 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14792 4883 4882 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14793 5183 4883 4882 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14794 4885 4884 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14795 5183 4885 4884 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14796 4887 4886 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14797 5183 4887 4886 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14798 4889 4888 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14799 5183 4889 4888 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14800 4891 4890 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14801 5183 4891 4890 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14802 4893 4892 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14803 5183 4893 4892 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14804 4895 4894 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14805 5183 4895 4894 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14806 4897 4896 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14807 5183 4897 4896 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14808 4899 4898 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14809 5183 4899 4898 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14810 4901 4900 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14811 5183 4901 4900 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14812 4903 4902 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14813 5183 4903 4902 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14814 4905 4904 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14815 5183 4905 4904 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14816 4907 4906 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14817 5183 4907 4906 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14818 4909 4908 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14819 5183 4909 4908 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14820 4911 4910 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14821 5183 4911 4910 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14822 4913 4912 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14823 5183 4913 4912 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14824 4915 4914 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14825 5183 4915 4914 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14826 4917 4916 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14827 5183 4917 4916 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14828 4919 4918 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14829 5183 4919 4918 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14830 4921 4920 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14831 5183 4921 4920 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14832 4923 4922 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14833 5183 4923 4922 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14834 4925 4924 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14835 5183 4925 4924 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14836 4927 4926 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14837 5183 4927 4926 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14838 4929 4928 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14839 5183 4929 4928 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14840 4931 4930 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14841 5183 4931 4930 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14842 4933 4932 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14843 5183 4933 4932 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14844 4935 4934 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14845 5183 4935 4934 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14846 4937 4936 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14847 5183 4937 4936 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14848 4939 4938 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14849 5183 4939 4938 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14850 4941 4940 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14851 5183 4941 4940 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14852 4943 4942 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14853 5183 4943 4942 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14854 4945 4944 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14855 5183 4945 4944 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14856 4947 4946 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14857 5183 4947 4946 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14858 4949 4948 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14859 5183 4949 4948 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14860 4951 4950 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14861 5183 4951 4950 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14862 4953 4952 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14863 5183 4953 4952 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14864 4955 4954 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14865 5183 4955 4954 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14866 4957 4956 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14867 5183 4957 4956 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14868 4959 4958 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14869 5183 4959 4958 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14870 4961 4960 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14871 5183 4961 4960 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14872 4963 4962 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14873 5183 4963 4962 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14874 4965 4964 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14875 5183 4965 4964 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14876 4967 4966 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14877 5183 4967 4966 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14878 4969 4968 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14879 5183 4969 4968 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14880 4971 4970 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14881 5183 4971 4970 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14882 4973 4972 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14883 5183 4973 4972 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14884 4975 4974 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14885 5183 4975 4974 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14886 4977 4976 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14887 5183 4977 4976 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14888 4979 4978 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14889 5183 4979 4978 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14890 4981 4980 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14891 5183 4981 4980 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14892 4983 4982 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14893 5183 4983 4982 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14894 4985 4984 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14895 5183 4985 4984 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14896 4987 4986 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14897 5183 4987 4986 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14898 4989 4988 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14899 5183 4989 4988 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14900 4991 4990 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14901 5183 4991 4990 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14902 4993 4992 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14903 5183 4993 4992 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14904 4995 4994 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14905 5183 4995 4994 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14906 4997 4996 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14907 5183 4997 4996 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14908 4999 4998 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14909 5183 4999 4998 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14910 5001 5000 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14911 5183 5001 5000 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14912 5003 5002 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14913 5183 5003 5002 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14914 5005 5004 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14915 5183 5005 5004 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14916 5007 5006 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14917 5183 5007 5006 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14918 5009 5008 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14919 5183 5009 5008 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14920 5011 5010 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14921 5183 5011 5010 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14922 5013 5012 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14923 5183 5013 5012 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14924 5015 5014 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14925 5183 5015 5014 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14926 5017 5016 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14927 5183 5017 5016 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14928 5019 5018 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14929 5183 5019 5018 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14930 5021 5020 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14931 5183 5021 5020 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14932 5023 5022 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14933 5183 5023 5022 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14934 5025 5024 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14935 5183 5025 5024 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14936 5027 5026 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14937 5183 5027 5026 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14938 5029 5028 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14939 5183 5029 5028 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14940 5031 5030 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14941 5183 5031 5030 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14942 5033 5032 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14943 5183 5033 5032 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14944 5035 5034 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14945 5183 5035 5034 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14946 5037 5036 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14947 5183 5037 5036 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14948 5039 5038 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14949 5183 5039 5038 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14950 5041 5040 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14951 5183 5041 5040 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14952 5043 5042 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14953 5183 5043 5042 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14954 5045 5044 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14955 5183 5045 5044 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14956 5047 5046 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14957 5183 5047 5046 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14958 5049 5048 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14959 5183 5049 5048 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14960 5051 5050 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14961 5183 5051 5050 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14962 5053 5052 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14963 5183 5053 5052 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14964 5055 5054 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14965 5183 5055 5054 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14966 5057 5056 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14967 5183 5057 5056 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14968 5059 5058 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14969 5183 5059 5058 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14970 5061 5060 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14971 5183 5061 5060 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14972 5063 5062 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14973 5183 5063 5062 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14974 5065 5064 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14975 5183 5065 5064 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14976 5067 5066 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14977 5183 5067 5066 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14978 5069 5068 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14979 5183 5069 5068 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14980 5071 5070 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14981 5183 5071 5070 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14982 5073 5072 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14983 5183 5073 5072 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14984 5075 5074 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14985 5183 5075 5074 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14986 5077 5076 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14987 5183 5077 5076 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14988 5079 5078 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14989 5183 5079 5078 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14990 5081 5080 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14991 5183 5081 5080 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14992 5083 5082 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14993 5183 5083 5082 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14994 5085 5084 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14995 5183 5085 5084 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14996 5087 5086 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14997 5183 5087 5086 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14998 5089 5088 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_14999 5183 5089 5088 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15000 5091 5090 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15001 5183 5091 5090 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15002 5093 5092 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15003 5183 5093 5092 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15004 5095 5094 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15005 5183 5095 5094 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15006 5097 5096 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15007 5183 5097 5096 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15008 5099 5098 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15009 5183 5099 5098 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15010 5101 5100 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15011 5183 5101 5100 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15012 5103 5102 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15013 5183 5103 5102 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15014 5105 5104 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15015 5183 5105 5104 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15016 5107 5106 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15017 5183 5107 5106 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15018 5109 5108 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15019 5183 5109 5108 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15020 5111 5110 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15021 5183 5111 5110 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15022 5113 5112 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15023 5183 5113 5112 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15024 5115 5114 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15025 5183 5115 5114 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15026 5117 5116 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15027 5183 5117 5116 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15028 5119 5118 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15029 5183 5119 5118 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15030 5121 5120 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15031 5183 5121 5120 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15032 5123 5122 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15033 5183 5123 5122 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15034 5125 5124 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15035 5183 5125 5124 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15036 5127 5126 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15037 5183 5127 5126 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15038 5129 5128 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15039 5183 5129 5128 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15040 5131 5130 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15041 5183 5131 5130 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15042 5133 5132 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15043 5183 5133 5132 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15044 5135 5134 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15045 5183 5135 5134 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15046 5137 5136 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15047 5183 5137 5136 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15048 5139 5138 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15049 5183 5139 5138 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15050 5141 5140 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15051 5183 5141 5140 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15052 5143 5142 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15053 5183 5143 5142 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15054 5145 5144 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15055 5183 5145 5144 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15056 5147 5146 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15057 5183 5147 5146 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15058 5149 5148 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15059 5183 5149 5148 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15060 5151 5150 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15061 5183 5151 5150 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15062 5153 5152 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15063 5183 5153 5152 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15064 5155 5154 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15065 5183 5155 5154 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15066 5157 5156 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15067 5183 5157 5156 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15068 5159 5158 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15069 5183 5159 5158 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15070 5161 5160 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15071 5183 5161 5160 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15072 5163 5162 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15073 5183 5163 5162 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15074 5165 5164 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15075 5183 5165 5164 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15076 5167 5166 5183 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15077 5183 5167 5166 5183 pmos L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_15078 5177 5168 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_15079 5183 5168 5168 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_15080 5170 5170 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_15081 5183 5170 5169 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_15082 5171 5172 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_15083 5183 5172 5172 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_15084 5173 5185 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_15085 5183 5175 5174 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_15086 5175 5185 5183 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_15087 5183 5185 5175 5183 pmos L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_15088 5185 5180 5183 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_15089 5183 5180 5185 5183 pmos L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_15090 5183 5176 5180 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_15091 5180 5177 5183 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_15092 5180 5179 5178 5183 pmos L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
.ends ram8x256

