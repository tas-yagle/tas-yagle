
.subckt ff i ck t vdd vss 
M1 s5 i vdd vdd TP L=0.18U W=2.232U AS=0.80352P AD=0.80352P PS=5.184U 
+ PD=5.184U 
M2 ms s4 vdd vdd TP L=0.72U W=0.432U AS=0.15552P AD=0.15552P PS=1.584U 
+ PD=1.584U 
M3 t sl vdd vdd TP L=0.18U W=4.212U AS=1.51632P AD=1.51632P PS=9.144U 
+ PD=9.144U 
M4 vdd sl s3 vdd TP L=0.18U W=0.972U AS=0.34992P AD=0.34992P PS=2.664U 
+ PD=2.664U 
M5 sl s3 vdd vdd TP L=0.72U W=0.432U AS=0.15552P AD=0.15552P PS=1.584U 
+ PD=1.584U 
M6 s1 ck vdd vdd TP L=0.18U W=3.312U AS=1.19232P AD=1.19232P PS=7.344U 
+ PD=7.344U 
M7 vdd ms s4 vdd TP L=0.18U W=0.972U AS=0.34992P AD=0.34992P PS=2.664U 
+ PD=2.664U 
M8 s2 s4 vdd vdd TP L=0.18U W=2.232U AS=0.80352P AD=0.80352P PS=5.184U 
+ PD=5.184U 
M9 s5 i vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P PS=3.024U 
+ PD=3.024U 
M10 t sl vss vss TN L=0.18U W=2.232U AS=0.80352P AD=0.80352P PS=5.184U 
+ PD=5.184U 
M11 vss sl s3 vss TN L=0.18U W=0.972U AS=0.34992P AD=0.34992P PS=2.664U 
+ PD=2.664U 
M12 s1 ck vss vss TN L=0.18U W=1.692U AS=0.60912P AD=0.60912P PS=4.104U 
+ PD=4.104U 
M13 ms ck s5 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P PS=3.024U 
+ PD=3.024U 
M14 vss ms s4 vss TN L=0.18U W=0.972U AS=0.34992P AD=0.34992P PS=2.664U 
+ PD=2.664U 
M15 vss s3 sl vss TN L=1.26U W=0.612U AS=0.22032P AD=0.22032P PS=1.944U 
+ PD=1.944U 
M16 sl s1 s2 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P PS=3.024U 
+ PD=3.024U 
M17 s2 s4 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P PS=3.024U 
+ PD=3.024U 
M18 vss s4 ms vss TN L=1.26U W=0.612U AS=0.22032P AD=0.22032P PS=1.944U 
+ PD=1.944U 
C0 i vss 1.15344e-15

C1 ck vss 1.6848e-15

C2 t vss 1.17936e-15

C3 s1 vss 1.2312e-15
C4 s3 vss 1.4256e-15
C5 sl vss 1.04976e-15
C6 s4 vss 2.3328e-15
C7 s5 vss 4.536e-16
C8 ms vss 9.72e-16

C9 s2 vss 6.0912e-16

.ends ff

