* Spice description of r256x8_6
* Spice driver version 700
* Date ( dd/mm/yyyy hh:mm:ss ): 20/09/2002 at 17:50:09

* INTERF adr[0] adr[1] adr[2] adr[3] adr[4] adr[5] adr[6] adr[7] ck[0] ck[1] 
* INTERF f[0] f[1] f[2] f[3] f[4] f[5] f[6] f[7] vdd vss 


.subckt r256x8_6 2356 2350 2351 2352 2344 2345 2346 2342 2258 1 2374 
+ 2371 2369 2367 2365 2363 2361 2359 2372 2375 
* NET 1 = ck[1] 
* NET 5 = rl/7.w1 
* NET 66 = rbl4/1/2.e0 
* NET 67 = rck.ckp 
* NET 77 = rl/7.e1 
* NET 78 = rl/7.tr_p 
* NET 79 = rl/7.w2 
* NET 80 = rl/7.w3 
* NET 81 = rl/7.w4 
* NET 262 = rbl4/1/2.e1 
* NET 263 = rbl4/1/2.e2 
* NET 264 = rbl4/1/2.e3 
* NET 282 = rl/6.e1 
* NET 283 = rl/6.tr_p 
* NET 284 = rl/6.w1 
* NET 285 = rl/6.w2 
* NET 286 = rl/6.w3 
* NET 287 = rl/6.w4 
* NET 528 = rbl4/1/2.e7 
* NET 529 = rbl4/1/2.e6 
* NET 530 = umf.e31 
* NET 531 = rbl4/1/2.e5 
* NET 552 = rl/5.w1 
* NET 553 = rl/5.w2 
* NET 554 = rl/5.w3 
* NET 735 = rbl4/1/2.e10 
* NET 736 = rbl4/1/2.e8 
* NET 737 = rbl4/1/2.e9 
* NET 754 = rl/5.e1 
* NET 755 = rl/5.tr_p 
* NET 756 = rl/5.w4 
* NET 757 = rl/4.w1 
* NET 758 = rl/4.w2 
* NET 983 = rbl4/1/2.e11 
* NET 1000 = rbl4/1/2.e14 
* NET 1001 = rbl4/1/2.e13 
* NET 1002 = rbl4/1/2.e12 
* NET 1023 = rl/4.e1 
* NET 1024 = rl/4.tr_p 
* NET 1025 = rl/4.w3 
* NET 1026 = rl/4.w4 
* NET 1027 = rl/3.w1 
* NET 1028 = rl/3.w2 
* NET 1209 = umf.e0 
* NET 1210 = rbl4/1/2.e15 
* NET 1211 = umf.e1 
* NET 1229 = rl/3.e1 
* NET 1230 = rl/3.tr_p 
* NET 1231 = rl/3.w3 
* NET 1232 = rl/3.w4 
* NET 1233 = rl/2.w1 
* NET 1234 = rl/2.w2 
* NET 1475 = umf.e2 
* NET 1476 = umf.e5 
* NET 1477 = umf.e4 
* NET 1478 = umf.e3 
* NET 1500 = rl/2.e1 
* NET 1501 = rl/2.tr_p 
* NET 1502 = rl/2.w3 
* NET 1503 = rl/2.w4 
* NET 1504 = rl/1.w1 
* NET 1685 = umf.e8 
* NET 1686 = umf.e7 
* NET 1687 = umf.e6 
* NET 1703 = rl/1.e1 
* NET 1704 = rl/1.tr_p 
* NET 1705 = rl/1.w2 
* NET 1706 = rl/1.w3 
* NET 1707 = rl/1.w4 
* NET 1708 = rl/0.w1 
* NET 1933 = umf.e9 
* NET 1950 = umf.e12 
* NET 1951 = umf.e11 
* NET 1952 = umf.e10 
* NET 1971 = rck.ck_02 
* NET 1975 = rl/0.e1 
* NET 1976 = rl/0.tr_p 
* NET 1977 = rck.ck_03 
* NET 1978 = rl/0.w2 
* NET 1979 = rl/0.w3 
* NET 1980 = rl/0.w4 
* NET 2161 = umf.e14 
* NET 2162 = umf.e13 
* NET 2163 = umf.e15 
* NET 2176 = rw2.n1 
* NET 2177 = rw3.n1 
* NET 2178 = rw1.n1 
* NET 2179 = rw0.n1 
* NET 2180 = rc116.n2 
* NET 2191 = rp4/15.s3 
* NET 2192 = rmx4/15.bl0_p 
* NET 2193 = rp4/14.s2 
* NET 2194 = rp4/14.s1 
* NET 2195 = rp4/15.s2 
* NET 2196 = rp4/15.s1 
* NET 2197 = rp4/14.s3 
* NET 2198 = rmx4/14.bl0_p 
* NET 2199 = rp4/13.s3 
* NET 2200 = rmx4/13.bl0_p 
* NET 2201 = rp4/12.s2 
* NET 2202 = rp4/13.s2 
* NET 2203 = rp4/12.s3 
* NET 2204 = rp4/12.s1 
* NET 2205 = rp4/13.s1 
* NET 2206 = rp4/11.s3 
* NET 2207 = rmx4/11.bl0_p 
* NET 2208 = rp4/11.s2 
* NET 2209 = rp4/11.s1 
* NET 2210 = rmx4/12.bl0_p 
* NET 2211 = rp4/10.s2 
* NET 2212 = rp4/10.s3 
* NET 2213 = rp4/10.s1 
* NET 2214 = rmx4/10.bl0_p 
* NET 2215 = rp4/9.s3 
* NET 2216 = rmx4/9.bl0_p 
* NET 2217 = rp4/9.s2 
* NET 2218 = rp4/9.s1 
* NET 2219 = rmx4/7.bl0_p 
* NET 2220 = rp4/7.s3 
* NET 2221 = rp4/8.s3 
* NET 2222 = rmx4/8.bl0_p 
* NET 2223 = rp4/8.s2 
* NET 2224 = rp4/8.s1 
* NET 2225 = rp4/6.s2 
* NET 2226 = rp4/6.s1 
* NET 2227 = rp4/7.s2 
* NET 2228 = rp4/7.s1 
* NET 2229 = rp4/5.s3 
* NET 2230 = rmx4/5.bl0_p 
* NET 2231 = rp4/6.s3 
* NET 2232 = rmx4/6.bl0_p 
* NET 2233 = rp4/4.s2 
* NET 2234 = rp4/4.s1 
* NET 2235 = rp4/5.s2 
* NET 2236 = rp4/5.s1 
* NET 2237 = rp4/3.s2 
* NET 2238 = rp4/3.s3 
* NET 2239 = rp4/3.s1 
* NET 2240 = rmx4/3.bl0_p 
* NET 2241 = rp4/4.s3 
* NET 2242 = rmx4/4.bl0_p 
* NET 2243 = rp4/2.s2 
* NET 2244 = rp4/2.s3 
* NET 2245 = rp4/2.s1 
* NET 2246 = rmx4/2.bl0_p 
* NET 2247 = rp4/1.s2 
* NET 2248 = rp4/1.s3 
* NET 2249 = rp4/1.s1 
* NET 2250 = rmx4/1.bl0_p 
* NET 2251 = x0.w2 
* NET 2252 = x0.w1 
* NET 2253 = x0.w0 
* NET 2254 = rp4/0.s2 
* NET 2255 = rp4/0.s3 
* NET 2256 = rp4/0.s1 
* NET 2257 = rmx4/0.bl0_p 
* NET 2258 = ck[0] 
* NET 2265 = rw1.inv 
* NET 2268 = x2.ck_11 
* NET 2270 = x1.w3 
* NET 2271 = rmx4/15.bit_p 
* NET 2272 = rmx4/14.bit_p 
* NET 2273 = rmx4/13.bit_p 
* NET 2274 = rmx4/12.bit_p 
* NET 2275 = rmx4/11.bit_p 
* NET 2276 = rmx4/10.bit_p 
* NET 2277 = rmx4/9.bit_p 
* NET 2278 = rmx4/8.bit_p 
* NET 2279 = rmx4/7.bit_p 
* NET 2280 = rmx4/6.bit_p 
* NET 2281 = rmx4/5.bit_p 
* NET 2282 = rmx4/4.bit_p 
* NET 2283 = rmx4/3.bit_p 
* NET 2284 = rmx4/2.bit_p 
* NET 2285 = rmx4/1.bit_p 
* NET 2286 = x1.ck_13 
* NET 2287 = rmx4/0.bit_p 
* NET 2290 = x2.n3b 
* NET 2292 = rmx2/7.i1 
* NET 2294 = rmx2/7.i0 
* NET 2296 = rmx2/7.s_p 
* NET 2300 = rmx2/6.s_p 
* NET 2302 = rmx2/5.i1 
* NET 2305 = rmx2/5.i0 
* NET 2306 = rmx2/5.s_p 
* NET 2308 = rmx2/3.i1 
* NET 2313 = rmx2/4.s_p 
* NET 2314 = rmx2/3.i0 
* NET 2316 = rmx2/3.s_p 
* NET 2321 = rmx2/1.i1 
* NET 2322 = rmx2/2.s_p 
* NET 2325 = rmx2/1.i0 
* NET 2326 = rmx2/1.s_p 
* NET 2329 = bf.e1 
* NET 2330 = bf.e0 
* NET 2332 = rmx2/0.s_p 
* NET 2342 = adr[7] 
* NET 2343 = rli/0.f 
* NET 2344 = adr[4] 
* NET 2345 = adr[5] 
* NET 2346 = adr[6] 
* NET 2347 = rw3.e1 
* NET 2348 = rli/2.f 
* NET 2349 = rli/1.f 
* NET 2350 = adr[1] 
* NET 2351 = adr[2] 
* NET 2352 = adr[3] 
* NET 2353 = x1.s5 
* NET 2354 = x2.s0 
* NET 2355 = rw3.e3 
* NET 2356 = adr[0] 
* NET 2357 = x0.s7 
* NET 2358 = rob/7.vss1 
* NET 2359 = f[7] 
* NET 2360 = rob/6.vss1 
* NET 2361 = f[6] 
* NET 2362 = rob/5.vss1 
* NET 2363 = f[5] 
* NET 2364 = rob/4.vss1 
* NET 2365 = f[4] 
* NET 2366 = rob/3.vss1 
* NET 2367 = f[3] 
* NET 2368 = rob/2.vss1 
* NET 2369 = f[2] 
* NET 2370 = rob/1.vss1 
* NET 2371 = f[1] 
* NET 2372 = vdd 
* NET 2373 = rob/0.vss1 
* NET 2374 = f[0] 
* NET 2375 = vss 
Mtr_02885 2 1 2372 2372 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02884 1971 2 2372 2372 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02883 2372 2 1971 2372 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02882 1971 2 2372 2372 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02881 2372 1971 1977 2372 tp L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02880 2372 1977 3 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02879 2372 3 4 2372 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02878 67 4 2372 2372 tp L=1U W=54U AS=108P AD=108P PS=112U PD=112U 
Mtr_02877 75 2342 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02876 2372 75 73 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02875 75 2345 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02874 72 2375 77 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02873 73 1971 72 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02872 2372 2346 75 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02871 78 1977 2372 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02870 2372 5 66 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02869 262 79 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02868 262 79 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02867 2372 66 5 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02866 79 262 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02865 2372 1977 5 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02864 79 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02863 2372 80 263 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02862 264 81 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02861 2372 80 263 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02860 264 81 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02859 2372 1977 80 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02858 81 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02857 81 264 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02856 2372 263 80 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02855 2372 5 66 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02854 281 2342 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02853 2372 281 278 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02852 281 2348 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02851 277 2375 282 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02850 278 1971 277 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02849 2372 2346 281 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02848 283 1977 2372 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02847 2372 284 530 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02846 531 285 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02845 531 285 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02844 2372 530 284 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02843 285 531 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02842 2372 1977 284 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02841 285 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02840 2372 286 529 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02839 528 287 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02838 2372 286 529 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02837 528 287 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02836 2372 1977 286 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02835 287 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02834 287 528 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02833 2372 529 286 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02832 2372 284 530 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02831 753 2342 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02830 2372 753 549 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02829 753 2345 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02828 548 2375 754 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02827 549 1971 548 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02826 2372 2349 753 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02825 755 1977 2372 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02824 2372 552 736 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02823 737 553 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02822 737 553 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02821 2372 736 552 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02820 553 737 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02819 2372 1977 552 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02818 553 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02817 2372 554 735 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02816 983 756 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02815 2372 554 735 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02814 983 756 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02813 2372 1977 554 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02812 756 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02811 756 983 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02810 2372 735 554 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02809 2372 552 736 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02808 1021 2342 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02807 2372 1021 751 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02806 1021 2348 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02805 750 2375 1023 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02804 751 1971 750 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02803 2372 2349 1021 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02802 1024 1977 2372 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02801 2372 757 1002 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02800 1001 758 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02799 1001 758 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02798 2372 1002 757 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02797 758 1001 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02796 2372 1977 757 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02795 758 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02794 2372 1025 1000 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02793 1210 1026 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02792 2372 1025 1000 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02791 1210 1026 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02790 2372 1977 1025 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02789 1026 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02788 1026 1210 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02787 2372 1000 1025 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02786 2372 757 1002 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02785 1226 2343 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02784 2372 1226 1020 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02783 1226 2345 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02782 1019 2375 1229 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02781 1020 1971 1019 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02780 2372 2346 1226 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02779 1230 1977 2372 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02778 2372 1027 1209 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02777 1211 1028 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02776 1211 1028 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02775 2372 1209 1027 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02774 1028 1211 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02773 2372 1977 1027 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02772 1028 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02771 2372 1231 1475 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02770 1478 1232 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02769 2372 1231 1475 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02768 1478 1232 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02767 2372 1977 1231 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02766 1232 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02765 1232 1478 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02764 2372 1475 1231 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02763 2372 1027 1209 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02762 1497 2343 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02761 2372 1497 1224 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02760 1497 2348 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02759 1225 2375 1500 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02758 1224 1971 1225 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02757 2372 2346 1497 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02756 1501 1977 2372 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02755 2372 1233 1477 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02754 1476 1234 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02753 1476 1234 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02752 2372 1477 1233 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02751 1234 1476 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02750 2372 1977 1233 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02749 1234 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02748 2372 1502 1687 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02747 1686 1503 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02746 2372 1502 1687 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02745 1686 1503 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02744 2372 1977 1502 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02743 1503 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02742 1503 1686 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02741 2372 1687 1502 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02740 2372 1233 1477 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02739 1700 2343 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02738 2372 1700 1495 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02737 1700 2345 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02736 1496 2375 1703 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02735 1495 1971 1496 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02734 2372 2349 1700 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02733 1704 1977 2372 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02732 2372 1504 1685 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02731 1933 1705 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02730 1933 1705 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02729 2372 1685 1504 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02728 1705 1933 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02727 2372 1977 1504 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02726 1705 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02725 2372 1706 1952 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02724 1951 1707 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02723 2372 1706 1952 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02722 1951 1707 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02721 2372 1977 1706 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02720 1707 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02719 1707 1951 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02718 2372 1952 1706 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02717 2372 1504 1685 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02716 1974 2343 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02715 2372 1974 1970 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02714 1974 2348 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02713 1969 2375 1975 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02712 1970 1971 1969 2372 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02711 2372 2349 1974 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02710 1976 1977 2372 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02709 2372 1708 1950 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02708 2162 1978 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02707 2162 1978 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02706 2372 1950 1708 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02705 1978 2162 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02704 2372 1977 1708 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02703 1978 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02702 2372 1979 2161 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02701 2163 1980 2372 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02700 2372 1979 2161 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02699 2163 1980 2372 2372 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02698 2372 1977 1979 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02697 1980 1977 2372 2372 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02696 1980 2163 2372 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02695 2372 2161 1979 2372 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02694 2372 1708 1950 2372 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02693 2268 2258 2372 2372 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02692 2372 2260 2177 2372 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02691 2177 2260 2372 2372 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02690 2260 2344 2372 2372 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02689 2372 2352 2260 2372 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02688 2372 2261 2176 2372 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02687 2176 2261 2372 2372 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02686 2372 2344 2261 2372 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02685 2261 2355 2372 2372 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02684 2372 2265 2178 2372 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02683 2178 2265 2372 2372 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02682 2265 2347 2372 2372 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02681 2372 2352 2265 2372 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02680 2372 2266 2179 2372 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02679 2179 2266 2372 2372 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02678 2372 2347 2266 2372 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02677 2266 2355 2372 2372 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02676 2372 2268 2180 2372 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02675 2286 2180 2372 2372 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02674 2372 2180 2286 2372 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02673 2286 2180 2372 2372 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02672 2372 2180 2286 2372 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02671 2372 2190 2253 2372 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02670 2252 2189 2372 2372 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02669 2372 2268 2189 2372 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02668 2189 2357 2372 2372 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02667 2372 2350 2189 2372 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02666 2190 2356 2372 2372 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02665 2372 2350 2190 2372 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02664 2372 2268 2190 2372 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02663 2372 2267 2251 2372 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02662 2270 2269 2372 2372 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02661 2267 2268 2372 2372 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02660 2267 2356 2372 2372 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02659 2269 2268 2372 2372 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02658 2372 2353 2269 2372 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02657 2269 2357 2372 2372 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02656 2372 2353 2267 2372 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02655 2372 2354 2290 2372 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02654 2290 2268 2372 2372 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02653 2372 2351 2291 2372 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02652 2291 2268 2372 2372 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02651 2330 2290 2372 2372 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02650 2372 2291 2329 2372 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02649 2271 2292 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02648 2372 2286 2271 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02647 2372 2271 2292 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02646 2272 2294 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02645 2372 2286 2272 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02644 2372 2272 2294 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02643 2273 2297 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02642 2372 2286 2273 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02641 2372 2273 2297 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02640 2274 2298 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02639 2372 2286 2274 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02638 2372 2274 2298 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02637 2275 2302 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02636 2372 2286 2275 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02635 2372 2275 2302 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02634 2276 2305 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02633 2372 2286 2276 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02632 2372 2276 2305 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02631 2277 2307 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02630 2372 2286 2277 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02629 2372 2277 2307 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02628 2278 2309 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02627 2372 2286 2278 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02626 2372 2278 2309 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02625 2279 2308 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02624 2372 2286 2279 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02623 2372 2279 2308 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02622 2280 2314 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02621 2372 2286 2280 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02620 2372 2280 2314 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02619 2281 2317 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02618 2372 2286 2281 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02617 2372 2281 2317 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02616 2282 2318 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02615 2372 2286 2282 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02614 2372 2282 2318 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02613 2283 2321 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02612 2372 2286 2283 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02611 2372 2283 2321 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02610 2284 2325 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02609 2372 2286 2284 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02608 2372 2284 2325 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02607 2285 2327 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02606 2372 2286 2285 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02605 2372 2285 2327 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02604 2287 2328 2372 2372 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02603 2372 2286 2287 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02602 2372 2287 2328 2372 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02601 2372 2342 2343 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02600 2343 2342 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02599 2343 2342 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02598 2372 2342 2343 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02597 2343 2342 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02596 2343 2342 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02595 2372 2346 2349 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02594 2349 2346 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02593 2349 2346 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02592 2372 2346 2349 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02591 2349 2346 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02590 2349 2346 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02589 2372 2345 2348 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02588 2348 2345 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02587 2348 2345 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02586 2372 2345 2348 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02585 2348 2345 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02584 2348 2345 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02583 2372 2344 2347 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02582 2347 2344 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02581 2347 2344 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02580 2372 2344 2347 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02579 2347 2344 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02578 2347 2344 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02577 2372 2352 2355 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02576 2355 2352 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02575 2355 2352 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02574 2372 2352 2355 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02573 2355 2352 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02572 2355 2352 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02571 2372 2351 2354 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02570 2354 2351 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02569 2354 2351 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02568 2372 2351 2354 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02567 2354 2351 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02566 2354 2351 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02565 2372 2350 2353 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02564 2353 2350 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02563 2353 2350 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02562 2372 2350 2353 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02561 2353 2350 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02560 2353 2350 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02559 2372 2356 2357 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02558 2357 2356 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02557 2357 2356 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02556 2372 2356 2357 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02555 2357 2356 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02554 2357 2356 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02553 2296 2286 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02552 2296 2334 2372 2372 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02551 2334 2296 2372 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02550 2372 2296 2334 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02549 2372 2358 2359 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02548 2359 2358 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02547 2372 2358 2359 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02546 2372 2358 2359 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02545 2359 2358 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02544 2372 2358 2359 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02543 2372 2334 2358 2372 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02542 2300 2286 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02541 2300 2335 2372 2372 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02540 2335 2300 2372 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02539 2372 2300 2335 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02538 2372 2360 2361 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02537 2361 2360 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02536 2372 2360 2361 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02535 2372 2360 2361 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02534 2361 2360 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02533 2372 2360 2361 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02532 2372 2335 2360 2372 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02531 2306 2286 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02530 2306 2336 2372 2372 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02529 2336 2306 2372 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02528 2372 2306 2336 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02527 2372 2362 2363 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02526 2363 2362 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02525 2372 2362 2363 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02524 2372 2362 2363 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02523 2363 2362 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02522 2372 2362 2363 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02521 2372 2336 2362 2372 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02520 2313 2286 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02519 2313 2337 2372 2372 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02518 2337 2313 2372 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02517 2372 2313 2337 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02516 2372 2364 2365 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02515 2365 2364 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02514 2372 2364 2365 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02513 2372 2364 2365 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02512 2365 2364 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02511 2372 2364 2365 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02510 2372 2337 2364 2372 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02509 2316 2286 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02508 2316 2338 2372 2372 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02507 2338 2316 2372 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02506 2372 2316 2338 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02505 2372 2366 2367 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02504 2367 2366 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02503 2372 2366 2367 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02502 2372 2366 2367 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02501 2367 2366 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02500 2372 2366 2367 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02499 2372 2338 2366 2372 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02498 2322 2286 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02497 2322 2339 2372 2372 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02496 2339 2322 2372 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02495 2372 2322 2339 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02494 2372 2368 2369 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02493 2369 2368 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02492 2372 2368 2369 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02491 2372 2368 2369 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02490 2369 2368 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02489 2372 2368 2369 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02488 2372 2339 2368 2372 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02487 2326 2286 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02486 2326 2340 2372 2372 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02485 2340 2326 2372 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02484 2372 2326 2340 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02483 2372 2370 2371 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02482 2371 2370 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02481 2372 2370 2371 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02480 2372 2370 2371 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02479 2371 2370 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02478 2372 2370 2371 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02477 2372 2340 2370 2372 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02476 2332 2286 2372 2372 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02475 2332 2341 2372 2372 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02474 2341 2332 2372 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02473 2372 2332 2341 2372 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02472 2372 2373 2374 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02471 2374 2373 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02470 2372 2373 2374 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02469 2372 2373 2374 2372 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02468 2374 2373 2372 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02467 2372 2373 2374 2372 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02466 2372 2341 2373 2372 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02465 2 1 2375 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02464 1971 2 2375 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02463 2375 2 1971 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02462 2375 1977 3 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02461 1977 1971 2375 2375 tn L=1U W=18U AS=36P AD=36P PS=40U PD=40U 
Mtr_02460 2375 3 4 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02459 67 4 2375 2375 tn L=1U W=28U AS=56P AD=56P PS=60U PD=60U 
Mtr_02458 2375 2375 77 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02457 75 2345 74 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02456 74 2346 76 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02455 76 2342 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02454 2375 75 77 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02453 77 1971 2375 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02452 78 2177 5 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02451 79 2176 78 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02450 78 2178 80 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02449 81 2179 78 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02448 2375 77 78 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02447 78 77 2375 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02446 2375 5 66 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02445 262 79 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02444 2375 80 263 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02443 264 81 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02442 2375 2375 282 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02441 281 2348 279 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02440 279 2346 280 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02439 280 2342 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02438 2375 281 282 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02437 282 1971 2375 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02436 283 2177 284 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02435 285 2176 283 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02434 283 2178 286 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02433 287 2179 283 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02432 2375 282 283 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02431 283 282 2375 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02430 2375 284 530 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02429 531 285 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02428 2375 286 529 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02427 528 287 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02426 2375 2375 754 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02425 753 2345 551 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02424 551 2349 550 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02423 550 2342 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02422 2375 753 754 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02421 754 1971 2375 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02420 755 2177 552 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02419 553 2176 755 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02418 755 2178 554 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02417 756 2179 755 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02416 2375 754 755 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02415 755 754 2375 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02414 2375 552 736 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02413 737 553 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02412 2375 554 735 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02411 983 756 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02410 2375 2375 1023 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02409 1021 2348 1022 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02408 1022 2349 752 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02407 752 2342 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02406 2375 1021 1023 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02405 1023 1971 2375 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02404 1024 2177 757 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02403 758 2176 1024 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02402 1024 2178 1025 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02401 1026 2179 1024 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02400 2375 1023 1024 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02399 1024 1023 2375 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02398 2375 757 1002 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02397 1001 758 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02396 2375 1025 1000 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02395 1210 1026 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02394 2375 2375 1229 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02393 1226 2345 1227 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02392 1227 2346 1228 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02391 1228 2343 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02390 2375 1226 1229 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02389 1229 1971 2375 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02388 1230 2177 1027 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02387 1028 2176 1230 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02386 1230 2178 1231 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02385 1232 2179 1230 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02384 2375 1229 1230 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02383 1230 1229 2375 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02382 2375 1027 1209 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02381 1211 1028 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02380 2375 1231 1475 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02379 1478 1232 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02378 2375 2375 1500 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02377 1497 2348 1499 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02376 1499 2346 1498 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02375 1498 2343 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02374 2375 1497 1500 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02373 1500 1971 2375 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02372 1501 2177 1233 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02371 1234 2176 1501 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02370 1501 2178 1502 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02369 1503 2179 1501 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02368 2375 1500 1501 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02367 1501 1500 2375 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02366 2375 1233 1477 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02365 1476 1234 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02364 2375 1502 1687 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02363 1686 1503 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02362 2375 2375 1703 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02361 1700 2345 1701 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02360 1701 2349 1702 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02359 1702 2343 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02358 2375 1700 1703 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02357 1703 1971 2375 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02356 1704 2177 1504 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02355 1705 2176 1704 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02354 1704 2178 1706 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02353 1707 2179 1704 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02352 2375 1703 1704 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02351 1704 1703 2375 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02350 2375 1504 1685 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02349 1933 1705 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02348 2375 1706 1952 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02347 1951 1707 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02346 2375 2375 1975 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02345 1974 2348 1972 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02344 1972 2349 1973 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02343 1973 2343 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02342 2375 1974 1975 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02341 1975 1971 2375 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02340 1976 2177 1708 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02339 1978 2176 1976 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02338 1976 2178 1979 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02337 1980 2179 1976 2375 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02336 2375 1975 1976 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02335 1976 1975 2375 2375 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02334 2375 1708 1950 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02333 2162 1978 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02332 2375 1979 2161 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02331 2163 1980 2375 2375 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02330 2375 2258 2268 2375 tn L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02329 2177 2260 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02328 2375 2260 2177 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02327 2260 2352 2259 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02326 2259 2344 2375 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02325 2176 2261 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02324 2375 2261 2176 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02323 2262 2355 2261 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02322 2375 2344 2262 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02321 2178 2265 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02320 2375 2265 2178 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02319 2264 2347 2375 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02318 2265 2352 2264 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02317 2375 2266 2179 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02316 2263 2355 2266 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02315 2375 2347 2263 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02314 2179 2266 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02313 2180 2268 2375 2375 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02312 2375 2180 2286 2375 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02311 2286 2180 2375 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02310 2187 2268 2189 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02309 2188 2357 2187 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02308 2375 2350 2188 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02307 2252 2189 2375 2375 tn L=1U W=26U AS=52P AD=52P PS=56U PD=56U 
Mtr_02306 2185 2268 2190 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02305 2186 2356 2185 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02304 2375 2350 2186 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02303 2375 2190 2253 2375 tn L=1U W=26U AS=52P AD=52P PS=56U PD=56U 
Mtr_02302 2183 2268 2375 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02301 2184 2353 2183 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02300 2267 2356 2184 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02299 2375 2267 2251 2375 tn L=1U W=26U AS=52P AD=52P PS=56U PD=56U 
Mtr_02298 2270 2269 2375 2375 tn L=1U W=26U AS=52P AD=52P PS=56U PD=56U 
Mtr_02297 2181 2268 2375 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02296 2182 2353 2181 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02295 2269 2357 2182 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02294 2290 2354 2288 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02293 2288 2268 2375 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02292 2330 2290 2375 2375 tn L=1U W=18U AS=36P AD=36P PS=40U PD=40U 
Mtr_02291 2375 2291 2329 2375 tn L=1U W=18U AS=36P AD=36P PS=40U PD=40U 
Mtr_02290 2291 2351 2289 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02289 2289 2268 2375 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02288 2192 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02287 2191 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02286 2195 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02285 2196 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02284 313 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02283 295 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02282 2375 530 312 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02281 2375 530 294 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02280 101 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02279 89 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02278 2375 263 102 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02277 2375 263 83 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02276 2375 66 12 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02275 2375 66 6 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02274 100 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02273 86 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02272 296 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02271 2375 530 288 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02270 90 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02269 2375 263 84 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02268 87 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02267 2375 66 7 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02266 297 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02265 2375 530 289 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02264 82 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02263 2375 263 85 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02262 88 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02261 2375 66 8 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02260 574 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02259 562 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02258 2375 736 575 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02257 2375 736 558 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02256 298 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02255 314 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02254 2375 529 315 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02253 2375 529 291 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02252 2375 529 292 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02251 299 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02250 2375 736 556 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02249 563 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02248 2375 529 293 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02247 290 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02246 2375 736 557 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02245 555 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02244 2375 735 573 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02243 2375 735 559 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02242 785 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02241 760 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02240 2375 735 560 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02239 2375 735 561 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02238 761 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02237 762 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02236 2375 1002 786 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02235 2375 1002 769 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02234 2375 1002 770 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02233 2375 1002 759 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02232 784 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02231 766 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02230 767 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02229 768 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02228 1049 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02227 2375 1000 783 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02226 1037 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02225 2375 1000 763 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02224 1035 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02223 2375 1000 764 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02222 2375 1000 765 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02221 1036 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02220 1260 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02219 1242 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02218 2375 1477 1261 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02217 2375 1477 1245 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02216 1262 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02215 1239 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02214 2375 1475 1259 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02213 2375 1475 1237 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02212 2375 1209 1048 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02211 2375 1209 1032 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02210 1047 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02209 1029 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02208 1243 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02207 2375 1477 1246 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02206 1240 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02205 2375 1475 1236 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02204 1030 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02203 2375 1209 1033 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02202 1244 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02201 2375 1477 1238 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02200 1241 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02199 2375 1475 1235 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02198 1031 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02197 2375 1209 1034 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02196 1735 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02195 1710 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02194 2375 1685 1525 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02193 2375 1685 1509 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02192 1512 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02191 1523 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02190 2375 1687 1524 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02189 2375 1687 1506 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02188 2375 1687 1507 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02187 1513 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02186 2375 1685 1510 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02185 1711 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02184 2375 1687 1508 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02183 1505 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02182 2375 1685 1511 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02181 1712 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02180 2375 1952 1736 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02179 2375 1952 1719 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02178 1734 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02177 1716 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02176 2375 1952 1720 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02175 2375 1952 1709 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02174 1717 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02173 1718 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02172 2375 1950 1733 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02171 2375 1950 1713 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02170 2375 1950 1714 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02169 2375 1950 1715 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02168 1999 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02167 1989 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02166 1981 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02165 1982 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02164 2001 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02163 2375 2161 2000 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02162 1983 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02161 2375 2161 1986 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02160 1984 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02159 2375 2161 1987 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02158 2375 2161 1988 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02157 1985 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02156 2271 2253 2192 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02155 2375 2271 2292 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02154 2195 2251 2271 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02153 2271 2270 2196 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02152 2271 2252 2191 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02151 2198 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02150 2197 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02149 2193 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02148 2194 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02147 309 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02146 310 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02145 2375 530 301 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02144 2375 530 302 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02143 94 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02142 95 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02141 2375 263 97 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02140 2375 263 98 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02139 2375 66 11 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02138 2375 66 9 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02137 91 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02136 92 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02135 311 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02134 2375 530 300 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02133 96 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02132 2375 263 99 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02131 93 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02130 2375 66 10 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02129 329 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02128 2375 530 330 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02127 114 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02126 2375 263 112 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02125 113 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02124 2375 66 16 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02123 564 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02122 565 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02121 2375 736 567 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02120 2375 736 568 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02119 304 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02118 303 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02117 2375 529 306 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02116 2375 529 307 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02115 2375 529 308 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02114 305 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02113 2375 736 569 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02112 566 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02111 2375 529 331 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02110 328 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02109 2375 736 587 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02108 586 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02107 2375 735 570 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02106 2375 735 571 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02105 774 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02104 775 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02103 2375 735 572 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02102 2375 735 585 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02101 776 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02100 802 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02099 2375 1002 771 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02098 2375 1002 772 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02097 2375 1002 773 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02096 2375 1002 801 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02095 780 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02094 781 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02093 782 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02092 800 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02091 1044 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02090 2375 1000 777 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02089 1045 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02088 2375 1000 778 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02087 1046 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02086 2375 1000 779 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02085 2375 1000 799 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02084 1059 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02083 1256 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02082 1257 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02081 2375 1477 1250 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02080 2375 1477 1251 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02079 1253 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02078 1254 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02077 2375 1475 1248 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02076 2375 1475 1249 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02075 2375 1209 1039 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02074 2375 1209 1040 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02073 1042 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02072 1043 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02071 1258 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02070 2375 1477 1252 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02069 1255 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02068 2375 1475 1247 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02067 1038 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02066 2375 1209 1041 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02065 1277 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02064 2375 1477 1278 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02063 1276 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02062 2375 1475 1272 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02061 1060 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02060 2375 1209 1061 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02059 1724 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02058 1725 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02057 2375 1685 1520 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02056 2375 1685 1521 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02055 1515 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02054 1514 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02053 2375 1687 1517 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02052 2375 1687 1518 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02051 2375 1687 1519 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02050 1516 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02049 2375 1685 1522 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02048 1726 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02047 2375 1687 1537 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02046 1536 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02045 2375 1685 1535 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02044 1752 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02043 2375 1952 1721 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02042 2375 1952 1722 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02041 1730 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02040 1731 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02039 2375 1952 1723 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02038 2375 1952 1751 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02037 1732 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02036 1750 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02035 2375 1950 1727 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02034 2375 1950 1728 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02033 2375 1950 1729 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02032 2375 1950 1749 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02031 1993 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02030 1994 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02029 1995 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02028 2012 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02027 1996 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02026 2375 2161 1990 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02025 1997 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02024 2375 2161 1991 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02023 1998 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02022 2375 2161 1992 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02021 2375 2161 2013 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02020 2011 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02019 2272 2253 2198 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02018 2375 2272 2294 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02017 2193 2251 2272 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02016 2272 2270 2194 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02015 2272 2252 2197 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02014 2200 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02013 2199 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02012 2202 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02011 2205 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02010 345 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02009 325 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02008 2375 530 344 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02007 2375 530 317 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02006 125 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02005 104 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02004 2375 263 126 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02003 2375 263 107 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02002 2375 66 20 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02001 2375 66 15 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02000 124 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01999 110 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01998 326 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01997 2375 530 318 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01996 105 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01995 2375 263 108 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01994 111 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01993 2375 66 13 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01992 327 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01991 2375 530 316 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01990 106 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01989 2375 263 109 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01988 103 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01987 2375 66 14 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01986 598 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01985 581 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01984 2375 736 599 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01983 2375 736 578 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01982 319 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01981 346 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01980 2375 529 347 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01979 2375 529 322 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01978 2375 529 323 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01977 320 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01976 2375 736 579 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01975 576 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01974 2375 529 324 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01973 321 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01972 2375 736 580 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01971 577 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01970 2375 735 597 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01969 2375 735 582 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01968 817 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01967 791 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01966 2375 735 583 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01965 2375 735 584 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01964 792 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01963 790 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01962 2375 1002 818 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01961 2375 1002 787 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01960 2375 1002 788 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01959 2375 1002 789 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01958 816 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01957 796 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01956 797 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01955 798 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01954 1073 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01953 2375 1000 815 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01952 1056 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01951 2375 1000 793 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01950 1057 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01949 2375 1000 794 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01948 2375 1000 795 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01947 1058 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01946 1292 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01945 1273 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01944 2375 1477 1293 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01943 2375 1477 1266 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01942 1294 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01941 1269 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01940 2375 1475 1291 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01939 2375 1475 1265 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01938 2375 1209 1072 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01937 2375 1209 1053 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01936 1071 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01935 1050 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01934 1274 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01933 2375 1477 1267 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01932 1270 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01931 2375 1475 1264 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01930 1051 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01929 2375 1209 1054 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01928 1275 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01927 2375 1477 1268 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01926 1271 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01925 2375 1475 1263 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01924 1052 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01923 2375 1209 1055 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01922 1767 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01921 1741 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01920 2375 1685 1549 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01919 2375 1685 1532 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01918 1526 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01917 1547 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01916 2375 1687 1548 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01915 2375 1687 1529 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01914 2375 1687 1530 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01913 1527 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01912 2375 1685 1533 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01911 1742 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01910 2375 1687 1531 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01909 1528 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01908 2375 1685 1534 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01907 1740 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01906 2375 1952 1768 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01905 2375 1952 1737 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01904 1766 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01903 1746 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01902 2375 1952 1738 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01901 2375 1952 1739 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01900 1747 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01899 1748 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01898 2375 1950 1765 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01897 2375 1950 1743 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01896 2375 1950 1744 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01895 2375 1950 1745 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01894 2023 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01893 2004 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01892 2005 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01891 2003 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01890 2025 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01889 2375 2161 2024 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01888 2006 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01887 2375 2161 2009 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01886 2007 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01885 2375 2161 2010 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01884 2375 2161 2002 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01883 2008 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01882 2273 2253 2200 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01881 2375 2273 2297 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01880 2202 2251 2273 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01879 2273 2270 2205 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01878 2273 2252 2199 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01877 2210 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01876 2203 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01875 2201 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01874 2204 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01873 341 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01872 342 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01871 2375 530 333 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01870 2375 530 334 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01869 118 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01868 119 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01867 2375 263 121 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01866 2375 263 122 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01865 2375 66 19 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01864 2375 66 17 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01863 115 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01862 116 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01861 343 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01860 2375 530 332 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01859 120 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01858 2375 263 123 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01857 117 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01856 2375 66 18 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01855 365 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01854 2375 530 366 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01853 141 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01852 2375 263 139 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01851 140 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01850 2375 66 25 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01849 588 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01848 589 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01847 2375 736 591 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01846 2375 736 592 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01845 336 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01844 335 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01843 2375 529 338 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01842 2375 529 339 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01841 2375 529 340 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01840 337 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01839 2375 736 593 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01838 590 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01837 2375 529 367 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01836 364 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01835 2375 736 614 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01834 613 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01833 2375 735 594 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01832 2375 735 595 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01831 806 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01830 807 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01829 2375 735 596 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01828 2375 735 612 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01827 808 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01826 837 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01825 2375 1002 803 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01824 2375 1002 804 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01823 2375 1002 805 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01822 2375 1002 838 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01821 812 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01820 813 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01819 814 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01818 836 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01817 1068 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01816 2375 1000 809 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01815 1069 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01814 2375 1000 810 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01813 1070 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01812 2375 1000 811 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01811 2375 1000 835 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01810 1086 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01809 1288 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01808 1289 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01807 2375 1477 1282 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01806 2375 1477 1283 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01805 1285 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01804 1286 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01803 2375 1475 1280 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01802 2375 1475 1281 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01801 2375 1209 1063 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01800 2375 1209 1064 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01799 1066 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01798 1067 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01797 1290 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01796 2375 1477 1284 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01795 1287 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01794 2375 1475 1279 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01793 1062 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01792 2375 1209 1065 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01791 1313 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01790 2375 1477 1314 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01789 1312 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01788 2375 1475 1308 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01787 1087 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01786 2375 1209 1088 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01785 1756 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01784 1757 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01783 2375 1685 1544 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01782 2375 1685 1545 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01781 1539 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01780 1538 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01779 2375 1687 1541 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01778 2375 1687 1542 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01777 2375 1687 1543 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01776 1540 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01775 2375 1685 1546 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01774 1758 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01773 2375 1687 1564 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01772 1563 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01771 2375 1685 1562 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01770 1787 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01769 2375 1952 1753 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01768 2375 1952 1754 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01767 1762 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01766 1763 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01765 2375 1952 1755 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01764 2375 1952 1788 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01763 1764 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01762 1786 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01761 2375 1950 1759 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01760 2375 1950 1760 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01759 2375 1950 1761 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01758 2375 1950 1785 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01757 2017 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01756 2018 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01755 2019 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01754 2040 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01753 2020 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01752 2375 2161 2014 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01751 2021 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01750 2375 2161 2015 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01749 2022 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01748 2375 2161 2016 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01747 2375 2161 2039 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01746 2038 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01745 2274 2253 2210 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01744 2375 2274 2298 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01743 2201 2251 2274 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01742 2274 2270 2204 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01741 2274 2252 2203 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01740 2207 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01739 2206 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01738 2208 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01737 2209 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01736 361 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01735 362 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01734 2375 530 351 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01733 2375 530 352 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01732 132 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01731 133 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01730 2375 263 136 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01729 2375 263 137 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01728 2375 66 23 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01727 2375 66 24 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01726 128 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01725 129 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01724 363 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01723 2375 530 348 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01722 134 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01721 2375 263 138 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01720 130 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01719 2375 66 21 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01718 353 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01717 2375 530 349 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01716 135 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01715 2375 263 127 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01714 131 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01713 2375 66 22 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01712 600 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01711 601 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01710 2375 736 604 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01709 2375 736 605 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01708 355 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01707 354 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01706 2375 529 358 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01705 2375 529 359 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01704 2375 529 360 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01703 356 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01702 2375 736 606 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01701 602 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01700 2375 529 350 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01699 357 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01698 2375 736 607 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01697 603 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01696 2375 735 608 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01695 2375 735 609 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01694 823 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01693 824 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01692 2375 735 610 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01691 2375 735 611 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01690 825 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01689 826 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01688 2375 1002 819 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01687 2375 1002 820 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01686 2375 1002 821 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01685 2375 1002 822 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01684 831 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01683 832 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01682 833 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01681 834 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01680 1083 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01679 2375 1000 827 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01678 1084 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01677 2375 1000 828 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01676 1085 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01675 2375 1000 829 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01674 2375 1000 830 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01673 1082 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01672 1309 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01671 1310 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01670 2375 1477 1301 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01669 2375 1477 1302 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01668 1305 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01667 1306 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01666 2375 1475 1297 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01665 2375 1475 1298 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01664 2375 1209 1077 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01663 2375 1209 1078 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01662 1081 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01661 1074 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01660 1311 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01659 2375 1477 1303 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01658 1307 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01657 2375 1475 1296 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01656 1075 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01655 2375 1209 1079 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01654 1300 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01653 2375 1477 1304 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01652 1299 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01651 2375 1475 1295 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01650 1076 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01649 2375 1209 1080 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01648 1773 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01647 1774 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01646 2375 1685 1558 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01645 2375 1685 1559 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01644 1551 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01643 1550 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01642 2375 1687 1554 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01641 2375 1687 1555 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01640 2375 1687 1556 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01639 1552 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01638 2375 1685 1560 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01637 1775 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01636 2375 1687 1557 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01635 1553 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01634 2375 1685 1561 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01633 1776 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01632 2375 1952 1769 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01631 2375 1952 1770 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01630 1781 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01629 1782 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01628 2375 1952 1771 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01627 2375 1952 1772 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01626 1783 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01625 1784 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01624 2375 1950 1777 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01623 2375 1950 1778 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01622 2375 1950 1779 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01621 2375 1950 1780 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01620 2036 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01619 2028 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01618 2026 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01617 2027 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01616 2037 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01615 2375 2161 2032 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01614 2029 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01613 2375 2161 2033 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01612 2030 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01611 2375 2161 2034 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01610 2375 2161 2035 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01609 2031 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01608 2275 2253 2207 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01607 2375 2275 2302 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01606 2208 2251 2275 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01605 2275 2270 2209 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01604 2275 2252 2206 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01603 2214 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01602 2212 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01601 2211 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01600 2213 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01599 378 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01598 379 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01597 2375 530 370 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01596 2375 530 371 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01595 152 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01594 153 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01593 2375 263 146 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01592 2375 263 147 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01591 2375 66 29 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01590 2375 66 28 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01589 150 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01588 151 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01587 380 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01586 2375 530 368 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01585 144 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01584 2375 263 148 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01583 142 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01582 2375 66 26 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01581 381 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01580 2375 530 369 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01579 145 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01578 2375 263 149 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01577 143 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01576 2375 66 27 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01575 625 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01574 626 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01573 2375 736 617 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01572 2375 736 618 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01571 383 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01570 382 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01569 2375 529 374 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01568 2375 529 375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01567 2375 529 376 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01566 372 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01565 2375 736 619 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01564 615 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01563 2375 529 377 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01562 373 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01561 2375 736 620 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01560 616 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01559 2375 735 621 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01558 2375 735 622 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01557 843 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01556 844 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01555 2375 735 623 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01554 2375 735 624 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01553 841 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01552 842 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01551 2375 1002 851 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01550 2375 1002 852 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01549 2375 1002 839 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01548 2375 1002 840 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01547 847 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01546 848 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01545 849 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01544 850 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01543 1100 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01542 2375 1000 853 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01541 1097 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01540 2375 1000 854 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01539 1098 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01538 2375 1000 845 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01537 2375 1000 846 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01536 1099 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01535 1325 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01534 1326 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01533 2375 1477 1329 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01532 2375 1477 1330 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01531 1321 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01530 1322 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01529 2375 1475 1317 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01528 2375 1475 1318 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01527 2375 1209 1096 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01526 2375 1209 1089 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01525 1092 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01524 1093 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01523 1327 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01522 2375 1477 1319 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01521 1323 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01520 2375 1475 1316 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01519 1094 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01518 2375 1209 1090 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01517 1328 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01516 2375 1477 1320 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01515 1324 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01514 2375 1475 1315 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01513 1095 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01512 2375 1209 1091 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01511 1793 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01510 1794 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01509 2375 1685 1571 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01508 2375 1685 1572 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01507 1576 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01506 1575 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01505 2375 1687 1567 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01504 2375 1687 1568 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01503 2375 1687 1569 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01502 1565 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01501 2375 1685 1573 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01500 1791 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01499 2375 1687 1570 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01498 1566 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01497 2375 1685 1574 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01496 1792 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01495 2375 1952 1801 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01494 2375 1952 1802 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01493 1797 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01492 1798 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01491 2375 1952 1789 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01490 2375 1952 1790 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01489 1799 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01488 1800 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01487 2375 1950 1803 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01486 2375 1950 1804 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01485 2375 1950 1795 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01484 2375 1950 1796 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01483 2046 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01482 2043 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01481 2044 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01480 2045 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01479 2047 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01478 2375 2161 2051 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01477 2048 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01476 2375 2161 2052 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01475 2049 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01474 2375 2161 2041 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01473 2375 2161 2042 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01472 2050 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01471 2276 2253 2214 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01470 2375 2276 2305 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01469 2211 2251 2276 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01468 2276 2270 2213 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01467 2276 2252 2212 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01466 2216 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01465 2215 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01464 2217 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01463 2218 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01462 397 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01461 398 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01460 2375 530 387 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01459 2375 530 388 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01458 159 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01457 160 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01456 2375 263 163 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01455 2375 263 164 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01454 2375 66 33 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01453 2375 66 30 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01452 155 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01451 156 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01450 399 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01449 2375 530 384 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01448 161 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01447 2375 263 165 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01446 157 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01445 2375 66 31 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01444 389 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01443 2375 530 385 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01442 162 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01441 2375 263 154 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01440 158 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01439 2375 66 32 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01438 627 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01437 628 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01436 2375 736 631 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01435 2375 736 632 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01434 391 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01433 390 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01432 2375 529 394 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01431 2375 529 395 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01430 2375 529 396 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01429 392 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01428 2375 736 633 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01427 629 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01426 2375 529 386 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01425 393 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01424 2375 736 634 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01423 630 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01422 2375 735 635 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01421 2375 735 636 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01420 859 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01419 860 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01418 2375 735 637 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01417 2375 735 638 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01416 861 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01415 862 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01414 2375 1002 855 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01413 2375 1002 856 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01412 2375 1002 857 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01411 2375 1002 858 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01410 867 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01409 868 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01408 869 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01407 870 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01406 1110 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01405 2375 1000 863 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01404 1111 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01403 2375 1000 864 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01402 1112 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01401 2375 1000 865 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01400 2375 1000 866 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01399 1109 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01398 1344 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01397 1345 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01396 2375 1477 1337 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01395 2375 1477 1338 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01394 1341 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01393 1342 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01392 2375 1475 1333 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01391 2375 1475 1334 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01390 2375 1209 1104 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01389 2375 1209 1105 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01388 1108 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01387 1101 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01386 1346 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01385 2375 1477 1339 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01384 1343 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01383 2375 1475 1332 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01382 1102 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01381 2375 1209 1106 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01380 1336 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01379 2375 1477 1340 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01378 1335 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01377 2375 1475 1331 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01376 1103 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01375 2375 1209 1107 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01374 1809 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01373 1810 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01372 2375 1685 1585 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01371 2375 1685 1586 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01370 1578 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01369 1577 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01368 2375 1687 1581 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01367 2375 1687 1582 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01366 2375 1687 1583 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01365 1579 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01364 2375 1685 1587 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01363 1811 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01362 2375 1687 1584 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01361 1580 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01360 2375 1685 1588 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01359 1812 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01358 2375 1952 1805 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01357 2375 1952 1806 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01356 1817 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01355 1818 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01354 2375 1952 1807 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01353 2375 1952 1808 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01352 1819 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01351 1820 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01350 2375 1950 1813 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01349 2375 1950 1814 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01348 2375 1950 1815 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01347 2375 1950 1816 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01346 2063 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01345 2055 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01344 2053 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01343 2054 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01342 2064 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01341 2375 2161 2059 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01340 2056 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01339 2375 2161 2060 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01338 2057 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01337 2375 2161 2061 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01336 2375 2161 2062 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01335 2058 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01334 2277 2253 2216 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01333 2375 2277 2307 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01332 2217 2251 2277 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01331 2277 2270 2218 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01330 2277 2252 2215 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01329 2222 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01328 2221 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01327 2223 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01326 2224 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01325 418 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01324 419 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01323 2375 530 410 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01322 2375 530 411 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01321 182 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01320 183 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01319 2375 263 176 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01318 2375 263 177 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01317 2375 66 38 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01316 2375 66 39 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01315 180 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01314 181 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01313 420 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01312 2375 530 408 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01311 174 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01310 2375 263 178 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01309 172 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01308 2375 66 36 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01307 421 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01306 2375 530 409 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01305 175 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01304 2375 263 179 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01303 173 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01302 2375 66 37 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01301 653 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01300 654 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01299 2375 736 645 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01298 2375 736 646 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01297 423 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01296 422 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01295 2375 529 414 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01294 2375 529 415 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01293 2375 529 416 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01292 412 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01291 2375 736 647 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01290 655 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01289 2375 529 417 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01288 413 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01287 2375 736 648 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01286 656 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01285 2375 735 649 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01284 2375 735 650 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01283 879 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01282 880 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01281 2375 735 651 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01280 2375 735 652 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01279 881 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01278 882 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01277 2375 1002 887 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01276 2375 1002 888 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01275 2375 1002 889 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01274 2375 1002 890 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01273 883 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01272 884 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01271 885 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01270 886 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01269 1130 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01268 2375 1000 891 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01267 1127 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01266 2375 1000 892 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01265 1128 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01264 2375 1000 893 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01263 2375 1000 894 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01262 1129 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01261 1365 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01260 1366 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01259 2375 1477 1369 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01258 2375 1477 1370 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01257 1361 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01256 1362 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01255 2375 1475 1357 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01254 2375 1475 1358 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01253 2375 1209 1126 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01252 2375 1209 1119 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01251 1122 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01250 1123 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01249 1367 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01248 2375 1477 1359 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01247 1363 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01246 2375 1475 1356 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01245 1124 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01244 2375 1209 1120 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01243 1368 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01242 2375 1477 1360 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01241 1364 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01240 2375 1475 1355 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01239 1125 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01238 2375 1209 1121 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01237 1829 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01236 1830 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01235 2375 1685 1599 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01234 2375 1685 1600 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01233 1604 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01232 1603 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01231 2375 1687 1595 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01230 2375 1687 1596 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01229 2375 1687 1597 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01228 1605 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01227 2375 1685 1601 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01226 1831 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01225 2375 1687 1598 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01224 1606 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01223 2375 1685 1602 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01222 1832 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01221 2375 1952 1837 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01220 2375 1952 1838 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01219 1833 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01218 1834 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01217 2375 1952 1839 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01216 2375 1952 1840 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01215 1835 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01214 1836 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01213 2375 1950 1841 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01212 2375 1950 1842 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01211 2375 1950 1843 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01210 2375 1950 1844 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01209 2079 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01208 2080 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01207 2072 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01206 2071 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01205 2081 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01204 2375 2161 2075 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01203 2082 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01202 2375 2161 2076 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01201 2073 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01200 2375 2161 2077 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01199 2375 2161 2078 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01198 2074 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01197 2278 2253 2222 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01196 2375 2278 2309 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01195 2223 2251 2278 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01194 2278 2270 2224 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01193 2278 2252 2221 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01192 2219 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01191 2220 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01190 2227 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01189 2228 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01188 437 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01187 438 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01186 2375 530 436 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01185 2375 530 432 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01184 195 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01183 190 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01182 2375 263 191 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01181 2375 263 192 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01180 2375 66 42 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01179 2375 66 43 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01178 193 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01177 194 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01176 407 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01175 2375 530 400 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01174 166 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01173 2375 263 168 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01172 170 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01171 2375 66 35 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01170 402 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01169 2375 530 401 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01168 167 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01167 2375 263 169 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01166 171 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01165 2375 66 34 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01164 665 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01163 666 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01162 2375 736 667 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01161 2375 736 668 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01160 433 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01159 439 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01158 2375 529 434 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01157 2375 529 435 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01156 2375 529 405 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01155 403 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01154 2375 736 644 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01153 641 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01152 2375 529 406 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01151 404 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01150 2375 736 643 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01149 642 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01148 2375 735 663 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01147 2375 735 664 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01146 909 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01145 910 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01144 2375 735 639 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01143 2375 735 640 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01142 875 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01141 876 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01140 2375 1002 907 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01139 2375 1002 908 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01138 2375 1002 873 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01137 2375 1002 874 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01136 905 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01135 906 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01134 871 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01133 872 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01132 1141 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01131 2375 1000 903 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01130 1142 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01129 2375 1000 904 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01128 1117 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01127 2375 1000 877 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01126 2375 1000 878 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01125 1118 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01124 1384 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01123 1385 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01122 2375 1477 1386 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01121 2375 1477 1381 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01120 1382 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01119 1383 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01118 2375 1475 1380 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01117 2375 1475 1378 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01116 2375 1209 1139 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01115 2375 1209 1138 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01114 1140 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01113 1137 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01112 1354 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01111 2375 1477 1350 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01110 1352 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01109 2375 1475 1348 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01108 1113 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01107 2375 1209 1115 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01106 1349 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01105 2375 1477 1351 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01104 1353 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01103 2375 1475 1347 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01102 1114 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01101 2375 1209 1116 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01100 1859 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01099 1860 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01098 2375 1685 1613 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01097 2375 1685 1614 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01096 1616 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01095 1615 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01094 2375 1687 1617 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01093 2375 1687 1618 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01092 2375 1687 1594 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01091 1591 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01090 2375 1685 1589 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01089 1825 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01088 2375 1687 1593 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01087 1592 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01086 2375 1685 1590 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01085 1826 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01084 2375 1952 1857 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01083 2375 1952 1858 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01082 1855 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01081 1856 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01080 2375 1952 1823 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01079 2375 1952 1824 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01078 1821 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01077 1822 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01076 2375 1950 1853 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01075 2375 1950 1854 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01074 2375 1950 1827 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01073 2375 1950 1828 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01072 2093 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01071 2092 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01070 2065 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01069 2066 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01068 2094 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01067 2375 2161 2090 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01066 2089 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01065 2375 2161 2091 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01064 2067 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01063 2375 2161 2069 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01062 2375 2161 2070 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01061 2068 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01060 2279 2253 2219 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01059 2375 2279 2308 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01058 2227 2251 2279 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01057 2279 2270 2228 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01056 2279 2252 2220 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01055 2232 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01054 2231 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01053 2225 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01052 2226 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01051 431 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01050 426 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01049 2375 530 424 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01048 2375 530 425 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01047 186 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01046 187 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01045 2375 263 188 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01044 2375 263 189 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01043 2375 66 40 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01042 2375 66 41 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01041 184 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01040 185 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01039 453 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01038 2375 530 452 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01037 207 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01036 2375 263 203 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01035 205 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01034 2375 66 47 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01033 454 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01032 2375 530 448 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01031 202 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01030 2375 263 204 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01029 206 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01028 2375 66 46 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01027 658 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01026 659 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01025 2375 736 660 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01024 2375 736 661 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01023 428 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01022 427 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01021 2375 529 429 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01020 2375 529 430 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01019 2375 529 450 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01018 455 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01017 2375 736 679 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01016 677 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01015 2375 529 451 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01014 449 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01013 2375 736 680 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01012 678 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01011 2375 735 662 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01010 2375 735 657 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01009 898 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01008 899 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01007 2375 735 675 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01006 2375 735 676 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01005 925 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01004 926 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01003 2375 1002 896 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01002 2375 1002 897 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01001 2375 1002 923 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01000 2375 1002 924 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00999 902 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00998 895 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00997 921 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00996 922 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00995 1136 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00994 2375 1000 900 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00993 1135 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00992 2375 1000 901 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00991 1153 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00990 2375 1000 919 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00989 2375 1000 920 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00988 1154 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00987 1379 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00986 1373 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00985 2375 1477 1374 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00984 2375 1477 1375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00983 1376 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00982 1377 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00981 2375 1475 1371 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00980 2375 1475 1372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00979 2375 1209 1132 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00978 2375 1209 1131 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00977 1133 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00976 1134 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00975 1400 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00974 2375 1477 1402 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00973 1398 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00972 2375 1475 1396 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00971 1151 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00970 2375 1209 1150 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00969 1401 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00968 2375 1477 1397 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00967 1399 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00966 2375 1475 1393 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00965 1152 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00964 2375 1209 1149 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00963 1848 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00962 1849 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00961 2375 1685 1612 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00960 2375 1685 1607 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00959 1609 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00958 1608 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00957 2375 1687 1610 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00956 2375 1687 1611 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00955 2375 1687 1629 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00954 1627 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00953 2375 1685 1625 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00952 1875 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00951 2375 1687 1630 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00950 1628 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00949 2375 1685 1626 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00948 1876 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00947 2375 1952 1846 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00946 2375 1952 1847 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00945 1852 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00944 1845 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00943 2375 1952 1873 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00942 2375 1952 1874 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00941 1871 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00940 1872 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00939 2375 1950 1850 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00938 2375 1950 1851 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00937 2375 1950 1869 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00936 2375 1950 1870 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00935 2086 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00934 2085 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00933 2105 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00932 2104 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00931 2087 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00930 2375 2161 2083 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00929 2088 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00928 2375 2161 2084 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00927 2106 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00926 2375 2161 2102 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00925 2375 2161 2103 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00924 2101 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00923 2280 2253 2232 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00922 2375 2280 2314 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00921 2225 2251 2280 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00920 2280 2270 2226 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00919 2280 2252 2231 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00918 2230 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00917 2229 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00916 2235 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00915 2236 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00914 473 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00913 474 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00912 2375 530 472 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00911 2375 530 468 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00910 222 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00909 217 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00908 2375 263 218 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00907 2375 263 219 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00906 2375 66 51 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00905 2375 66 52 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00904 220 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00903 221 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00902 446 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00901 2375 530 441 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00900 197 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00899 2375 263 199 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00898 201 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00897 2375 66 44 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00896 447 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00895 2375 530 440 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00894 198 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00893 2375 263 200 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00892 196 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00891 2375 66 45 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00890 692 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00889 693 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00888 2375 736 694 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00887 2375 736 695 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00886 469 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00885 475 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00884 2375 529 470 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00883 2375 529 471 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00882 2375 529 444 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00881 442 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00880 2375 736 671 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00879 669 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00878 2375 529 445 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00877 443 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00876 2375 736 672 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00875 670 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00874 2375 735 690 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00873 2375 735 691 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00872 945 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00871 946 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00870 2375 735 673 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00869 2375 735 674 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00868 914 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00867 913 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00866 2375 1002 943 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00865 2375 1002 944 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00864 2375 1002 911 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00863 2375 1002 912 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00862 941 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00861 942 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00860 917 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00859 918 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00858 1168 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00857 2375 1000 939 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00856 1169 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00855 2375 1000 940 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00854 1147 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00853 2375 1000 915 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00852 2375 1000 916 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00851 1148 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00850 1420 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00849 1421 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00848 2375 1477 1422 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00847 2375 1477 1417 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00846 1418 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00845 1419 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00844 2375 1475 1416 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00843 2375 1475 1414 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00842 2375 1209 1166 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00841 2375 1209 1165 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00840 1167 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00839 1164 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00838 1394 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00837 2375 1477 1389 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00836 1391 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00835 2375 1475 1388 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00834 1143 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00833 2375 1209 1145 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00832 1395 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00831 2375 1477 1390 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00830 1392 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00829 2375 1475 1387 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00828 1144 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00827 2375 1209 1146 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00826 1895 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00825 1896 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00824 2375 1685 1640 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00823 2375 1685 1641 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00822 1643 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00821 1642 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00820 2375 1687 1644 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00819 2375 1687 1645 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00818 2375 1687 1621 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00817 1619 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00816 2375 1685 1623 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00815 1864 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00814 2375 1687 1622 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00813 1620 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00812 2375 1685 1624 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00811 1863 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00810 2375 1952 1893 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00809 2375 1952 1894 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00808 1891 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00807 1892 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00806 2375 1952 1861 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00805 2375 1952 1862 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00804 1867 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00803 1868 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00802 2375 1950 1889 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00801 2375 1950 1890 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00800 2375 1950 1865 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00799 2375 1950 1866 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00798 2120 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00797 2119 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00796 2097 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00795 2096 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00794 2121 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00793 2375 2161 2117 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00792 2116 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00791 2375 2161 2118 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00790 2098 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00789 2375 2161 2100 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00788 2375 2161 2095 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00787 2099 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00786 2281 2253 2230 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00785 2375 2281 2317 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00784 2235 2251 2281 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00783 2281 2270 2236 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00782 2281 2252 2229 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00781 2242 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00780 2241 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00779 2233 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00778 2234 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00777 467 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00776 459 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00775 2375 530 457 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00774 2375 530 458 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00773 211 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00772 212 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00771 2375 263 214 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00770 2375 263 215 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00769 2375 66 49 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00768 2375 66 50 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00767 208 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00766 209 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00765 460 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00764 2375 530 456 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00763 213 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00762 2375 263 216 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00761 210 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00760 2375 66 48 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00759 495 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00758 2375 530 493 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00757 236 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00756 2375 263 237 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00755 235 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00754 2375 66 57 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00753 683 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00752 684 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00751 2375 736 686 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00750 2375 736 687 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00749 462 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00748 461 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00747 2375 529 464 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00746 2375 529 465 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00745 2375 529 466 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00744 463 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00743 2375 736 688 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00742 685 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00741 2375 529 494 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00740 492 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00739 2375 736 710 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00738 709 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00737 2375 735 689 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00736 2375 735 681 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00735 932 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00734 933 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00733 2375 735 682 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00732 2375 735 708 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00731 934 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00730 965 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00729 2375 1002 929 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00728 2375 1002 930 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00727 2375 1002 931 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00726 2375 1002 966 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00725 938 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00724 927 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00723 928 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00722 964 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00721 1163 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00720 2375 1000 935 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00719 1161 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00718 2375 1000 936 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00717 1162 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00716 2375 1000 937 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00715 2375 1000 963 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00714 1184 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00713 1415 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00712 1406 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00711 2375 1477 1408 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00710 2375 1477 1409 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00709 1411 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00708 1412 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00707 2375 1475 1404 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00706 2375 1475 1405 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00705 2375 1209 1157 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00704 2375 1209 1155 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00703 1158 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00702 1159 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00701 1407 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00700 2375 1477 1410 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00699 1413 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00698 2375 1475 1403 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00697 1160 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00696 2375 1209 1156 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00695 1442 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00694 2375 1477 1440 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00693 1441 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00692 2375 1475 1435 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00691 1182 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00690 2375 1209 1183 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00689 1882 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00688 1883 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00687 2375 1685 1639 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00686 2375 1685 1631 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00685 1634 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00684 1633 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00683 2375 1687 1636 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00682 2375 1687 1637 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00681 2375 1687 1638 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00680 1635 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00679 2375 1685 1632 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00678 1884 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00677 2375 1687 1660 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00676 1659 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00675 2375 1685 1658 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00674 1915 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00673 2375 1952 1879 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00672 2375 1952 1880 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00671 1888 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00670 1877 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00669 2375 1952 1881 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00668 2375 1952 1916 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00667 1878 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00666 1914 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00665 2375 1950 1885 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00664 2375 1950 1886 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00663 2375 1950 1887 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00662 2375 1950 1913 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00661 2112 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00660 2110 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00659 2111 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00658 2135 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00657 2113 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00656 2375 2161 2107 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00655 2114 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00654 2375 2161 2108 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00653 2115 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00652 2375 2161 2109 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00651 2375 2161 2136 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00650 2134 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00649 2282 2253 2242 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00648 2375 2282 2318 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00647 2233 2251 2282 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00646 2282 2270 2234 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00645 2282 2252 2241 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00644 2240 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00643 2238 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00642 2237 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00641 2239 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00640 488 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00639 489 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00638 2375 530 478 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00637 2375 530 479 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00636 227 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00635 228 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00634 2375 263 231 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00633 2375 263 232 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00632 2375 66 56 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00631 2375 66 53 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00630 223 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00629 224 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00628 490 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00627 2375 530 476 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00626 229 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00625 2375 263 233 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00624 225 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00623 2375 66 54 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00622 491 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00621 2375 530 477 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00620 230 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00619 2375 263 234 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00618 226 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00617 2375 66 55 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00616 696 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00615 697 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00614 2375 736 700 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00613 2375 736 701 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00612 481 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00611 480 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00610 2375 529 484 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00609 2375 529 485 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00608 2375 529 486 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00607 482 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00606 2375 736 702 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00605 698 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00604 2375 529 487 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00603 483 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00602 2375 736 703 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00601 699 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00600 2375 735 704 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00599 2375 735 705 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00598 951 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00597 952 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00596 2375 735 706 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00595 2375 735 707 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00594 953 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00593 954 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00592 2375 1002 947 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00591 2375 1002 948 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00590 2375 1002 949 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00589 2375 1002 950 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00588 959 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00587 960 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00586 961 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00585 962 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00584 1178 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00583 2375 1000 955 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00582 1179 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00581 2375 1000 956 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00580 1180 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00579 2375 1000 957 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00578 2375 1000 958 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00577 1181 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00576 1436 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00575 1437 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00574 2375 1477 1427 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00573 2375 1477 1428 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00572 1431 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00571 1432 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00570 2375 1475 1425 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00569 2375 1475 1426 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00568 2375 1209 1172 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00567 2375 1209 1173 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00566 1176 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00565 1177 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00564 1438 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00563 2375 1477 1429 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00562 1433 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00561 2375 1475 1424 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00560 1170 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00559 2375 1209 1174 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00558 1439 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00557 2375 1477 1430 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00556 1434 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00555 2375 1475 1423 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00554 1171 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00553 2375 1209 1175 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00552 1901 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00551 1902 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00550 2375 1685 1654 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00549 2375 1685 1655 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00548 1647 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00547 1646 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00546 2375 1687 1650 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00545 2375 1687 1651 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00544 2375 1687 1652 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00543 1648 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00542 2375 1685 1656 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00541 1903 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00540 2375 1687 1653 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00539 1649 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00538 2375 1685 1657 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00537 1904 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00536 2375 1952 1897 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00535 2375 1952 1898 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00534 1909 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00533 1910 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00532 2375 1952 1899 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00531 2375 1952 1900 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00530 1911 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00529 1912 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00528 2375 1950 1905 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00527 2375 1950 1906 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00526 2375 1950 1907 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00525 2375 1950 1908 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00524 2126 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00523 2127 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00522 2128 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00521 2129 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00520 2130 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00519 2375 2161 2122 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00518 2131 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00517 2375 2161 2123 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00516 2132 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00515 2375 2161 2124 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00514 2375 2161 2125 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00513 2133 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00512 2283 2253 2240 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00511 2375 2283 2321 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00510 2237 2251 2283 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00509 2283 2270 2239 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00508 2283 2252 2238 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00507 2246 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00506 2244 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00505 2243 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00504 2245 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00503 508 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00502 509 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00501 2375 530 498 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00500 2375 530 499 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00499 242 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00498 243 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00497 2375 263 246 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00496 2375 263 247 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00495 2375 66 58 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00494 2375 66 59 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00493 238 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00492 239 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00491 510 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00490 2375 530 496 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00489 244 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00488 2375 263 248 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00487 240 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00486 2375 66 60 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00485 511 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00484 2375 530 497 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00483 245 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00482 2375 263 249 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00481 241 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00480 2375 66 61 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00479 711 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00478 712 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00477 2375 736 715 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00476 2375 736 716 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00475 501 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00474 500 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00473 2375 529 504 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00472 2375 529 505 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00471 2375 529 506 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00470 502 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00469 2375 736 717 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00468 713 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00467 2375 529 507 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00466 503 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00465 2375 736 718 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00464 714 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00463 2375 735 719 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00462 2375 735 720 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00461 971 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00460 972 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00459 2375 735 721 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00458 2375 735 722 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00457 973 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00456 974 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00455 2375 1002 967 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00454 2375 1002 968 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00453 2375 1002 969 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00452 2375 1002 970 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00451 979 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00450 980 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00449 981 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00448 982 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00447 1193 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00446 2375 1000 975 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00445 1194 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00444 2375 1000 976 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00443 1195 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00442 2375 1000 977 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00441 2375 1000 978 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00440 1196 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00439 1455 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00438 1456 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00437 2375 1477 1447 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00436 2375 1477 1448 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00435 1451 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00434 1452 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00433 2375 1475 1445 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00432 2375 1475 1446 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00431 2375 1209 1187 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00430 2375 1209 1188 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00429 1191 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00428 1192 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00427 1457 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00426 2375 1477 1449 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00425 1453 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00424 2375 1475 1444 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00423 1185 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00422 2375 1209 1189 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00421 1458 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00420 2375 1477 1450 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00419 1454 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00418 2375 1475 1443 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00417 1186 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00416 2375 1209 1190 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00415 1921 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00414 1922 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00413 2375 1685 1669 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00412 2375 1685 1670 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00411 1662 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00410 1661 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00409 2375 1687 1665 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00408 2375 1687 1666 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00407 2375 1687 1667 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00406 1663 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00405 2375 1685 1671 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00404 1923 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00403 2375 1687 1668 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00402 1664 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00401 2375 1685 1672 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00400 1924 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00399 2375 1952 1917 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00398 2375 1952 1918 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00397 1929 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00396 1930 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00395 2375 1952 1919 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00394 2375 1952 1920 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00393 1931 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00392 1932 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00391 2375 1950 1925 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00390 2375 1950 1926 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00389 2375 1950 1927 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00388 2375 1950 1928 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00387 2141 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00386 2142 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00385 2143 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00384 2144 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00383 2145 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00382 2375 2161 2137 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00381 2146 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00380 2375 2161 2138 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00379 2147 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00378 2375 2161 2139 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00377 2375 2161 2140 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00376 2148 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00375 2284 2253 2246 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00374 2375 2284 2325 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00373 2243 2251 2284 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00372 2284 2270 2245 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00371 2284 2252 2244 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00370 2250 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00369 2248 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00368 2247 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00367 2249 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00366 520 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00365 521 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00364 2375 530 513 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00363 2375 530 514 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00362 258 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00361 259 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00360 2375 263 250 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00359 2375 263 251 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00358 2375 66 65 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00357 2375 66 62 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00356 254 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00355 255 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00354 522 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00353 2375 530 515 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00352 260 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00351 2375 263 252 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00350 256 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00349 2375 66 63 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00348 523 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00347 2375 530 512 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00346 261 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00345 2375 263 253 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00344 257 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00343 2375 66 64 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00342 731 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00341 732 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00340 2375 736 723 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00339 2375 736 724 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00338 525 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00337 524 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00336 2375 529 516 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00335 2375 529 517 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00334 2375 529 518 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00333 526 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00332 2375 736 725 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00331 733 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00330 2375 529 519 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00329 527 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00328 2375 736 726 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00327 734 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00326 2375 735 727 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00325 2375 735 728 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00324 984 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00323 985 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00322 2375 735 729 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00321 2375 735 730 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00320 986 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00319 987 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00318 2375 1002 992 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00317 2375 1002 993 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00316 2375 1002 994 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00315 2375 1002 995 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00314 988 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00313 989 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00312 990 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00311 991 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00310 1207 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00309 2375 1000 996 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00308 1208 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00307 2375 1000 997 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00306 1205 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00305 2375 1000 998 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00304 2375 1000 999 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00303 1206 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00302 1467 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00301 1468 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00300 2375 1477 1471 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00299 2375 1477 1472 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00298 1463 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00297 1464 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00296 2375 1475 1461 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00295 2375 1475 1462 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00294 2375 1209 1203 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00293 2375 1209 1204 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00292 1199 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00291 1200 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00290 1469 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00289 2375 1477 1473 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00288 1465 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00287 2375 1475 1460 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00286 1201 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00285 2375 1209 1197 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00284 1470 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00283 2375 1477 1474 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00282 1466 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00281 2375 1475 1459 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00280 1202 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00279 2375 1209 1198 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00278 1934 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00277 1935 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00276 2375 1685 1677 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00275 2375 1685 1678 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00274 1682 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00273 1681 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00272 2375 1687 1673 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00271 2375 1687 1674 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00270 2375 1687 1675 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00269 1683 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00268 2375 1685 1679 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00267 1936 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00266 2375 1687 1676 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00265 1684 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00264 2375 1685 1680 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00263 1937 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00262 2375 1952 1942 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00261 2375 1952 1943 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00260 1938 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00259 1939 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00258 2375 1952 1944 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00257 2375 1952 1945 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00256 1940 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00255 1941 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00254 2375 1950 1946 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00253 2375 1950 1947 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00252 2375 1950 1948 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00251 2375 1950 1949 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00250 2151 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00249 2152 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00248 2149 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00247 2150 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00246 2153 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00245 2375 2161 2157 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00244 2154 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00243 2375 2161 2158 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00242 2155 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00241 2375 2161 2159 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00240 2375 2161 2160 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00239 2156 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00238 2285 2253 2250 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00237 2375 2285 2327 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00236 2247 2251 2285 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00235 2285 2270 2249 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00234 2285 2252 2248 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00233 2257 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00232 2255 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00231 2254 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00230 2256 67 2372 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00229 544 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00228 545 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00227 2375 530 534 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00226 2375 530 535 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00225 269 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00224 270 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00223 2375 263 273 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00222 2375 263 274 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00221 2375 66 68 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00220 2375 66 69 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00219 265 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00218 266 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00217 546 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00216 2375 530 532 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00215 271 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00214 2375 263 275 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00213 267 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00212 2375 66 70 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00211 547 531 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00210 2375 530 533 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00209 272 264 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00208 2375 263 276 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00207 268 262 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00206 2375 66 71 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00205 738 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00204 739 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00203 2375 736 742 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00202 2375 736 743 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00201 537 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00200 536 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00199 2375 529 540 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00198 2375 529 541 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00197 2375 529 542 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00196 538 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00195 2375 736 744 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00194 740 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00193 2375 529 543 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00192 539 528 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00191 2375 736 745 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00190 741 737 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00189 2375 735 746 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00188 2375 735 747 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00187 1007 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00186 1008 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00185 2375 735 748 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00184 2375 735 749 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00183 1009 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00182 1010 983 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00181 2375 1002 1003 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00180 2375 1002 1004 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00179 2375 1002 1005 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00178 2375 1002 1006 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00177 1015 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00176 1016 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00175 1017 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00174 1018 1001 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00173 1220 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00172 2375 1000 1011 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00171 1221 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00170 2375 1000 1012 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00169 1222 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00168 2375 1000 1013 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00167 2375 1000 1014 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00166 1223 1210 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00165 1491 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00164 1492 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00163 2375 1477 1483 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00162 2375 1477 1484 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00161 1487 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00160 1488 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00159 2375 1475 1481 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00158 2375 1475 1482 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00157 2375 1209 1214 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00156 2375 1209 1215 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00155 1218 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00154 1219 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00153 1493 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00152 2375 1477 1485 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00151 1489 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00150 2375 1475 1480 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00149 1212 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00148 2375 1209 1216 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00147 1494 1476 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00146 2375 1477 1486 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00145 1490 1478 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00144 2375 1475 1479 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00143 1213 1211 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00142 2375 1209 1217 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00141 1957 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00140 1958 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00139 2375 1685 1696 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00138 2375 1685 1697 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00137 1689 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00136 1688 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00135 2375 1687 1692 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00134 2375 1687 1693 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00133 2375 1687 1694 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00132 1690 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00131 2375 1685 1698 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00130 1959 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00129 2375 1687 1695 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00128 1691 1686 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00127 2375 1685 1699 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00126 1960 1933 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00125 2375 1952 1953 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00124 2375 1952 1954 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00123 1965 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00122 1966 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00121 2375 1952 1955 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00120 2375 1952 1956 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00119 1967 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00118 1968 1951 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00117 2375 1950 1961 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00116 2375 1950 1962 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00115 2375 1950 1963 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00114 2375 1950 1964 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00113 2168 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00112 2169 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00111 2170 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00110 2171 2162 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00109 2172 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00108 2375 2161 2164 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00107 2173 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00106 2375 2161 2165 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00105 2174 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00104 2375 2161 2166 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00103 2375 2161 2167 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00102 2175 2163 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00101 2287 2253 2257 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00100 2375 2287 2328 2375 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00099 2254 2251 2287 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00098 2287 2270 2256 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00097 2287 2252 2255 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00096 2375 2342 2343 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00095 2343 2342 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00094 2343 2342 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00093 2375 2346 2349 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00092 2349 2346 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00091 2349 2346 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00090 2375 2345 2348 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00089 2348 2345 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00088 2348 2345 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00087 2375 2344 2347 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00086 2347 2344 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00085 2347 2344 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00084 2375 2352 2355 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00083 2355 2352 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00082 2355 2352 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00081 2375 2351 2354 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00080 2354 2351 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00079 2354 2351 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00078 2375 2350 2353 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00077 2353 2350 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00076 2353 2350 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00075 2375 2356 2357 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00074 2357 2356 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00073 2357 2356 2375 2375 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00072 2375 2294 2295 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00071 2295 2329 2296 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00070 2296 2330 2293 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00069 2293 2292 2375 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00068 2334 2296 2375 2375 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00067 2359 2358 2375 2375 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00066 2375 2358 2359 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00065 2375 2334 2358 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00064 2359 2358 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00063 2375 2298 2301 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00062 2301 2329 2300 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00061 2300 2330 2299 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00060 2299 2297 2375 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00059 2335 2300 2375 2375 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00058 2361 2360 2375 2375 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00057 2375 2360 2361 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00056 2375 2335 2360 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00055 2361 2360 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00054 2375 2305 2304 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00053 2304 2329 2306 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00052 2306 2330 2303 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00051 2303 2302 2375 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00050 2336 2306 2375 2375 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00049 2363 2362 2375 2375 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00048 2375 2362 2363 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00047 2375 2336 2362 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00046 2363 2362 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00045 2375 2309 2312 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00044 2312 2329 2313 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00043 2313 2330 2311 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00042 2311 2307 2375 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00041 2337 2313 2375 2375 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00040 2365 2364 2375 2375 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00039 2375 2364 2365 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00038 2375 2337 2364 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00037 2365 2364 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00036 2375 2314 2315 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00035 2315 2329 2316 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00034 2316 2330 2310 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00033 2310 2308 2375 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00032 2338 2316 2375 2375 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00031 2367 2366 2375 2375 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00030 2375 2366 2367 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00029 2375 2338 2366 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00028 2367 2366 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00027 2375 2318 2320 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00026 2320 2329 2322 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00025 2322 2330 2319 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00024 2319 2317 2375 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00023 2339 2322 2375 2375 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00022 2369 2368 2375 2375 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00021 2375 2368 2369 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00020 2375 2339 2368 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00019 2369 2368 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00018 2375 2325 2323 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00017 2323 2329 2326 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00016 2326 2330 2324 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00015 2324 2321 2375 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00014 2340 2326 2375 2375 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00013 2371 2370 2375 2375 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00012 2375 2370 2371 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 2375 2340 2370 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00010 2371 2370 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 2375 2328 2333 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00008 2333 2329 2332 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00007 2332 2330 2331 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00006 2331 2327 2375 2375 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00005 2341 2332 2375 2375 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00004 2374 2373 2375 2375 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00003 2375 2373 2374 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 2375 2341 2373 2375 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00001 2374 2373 2375 2375 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
.ends r256x8_6

