
.subckt cpu2901 zero y_3 y_2 y_1 y_0 vssi vsse vddi vdde test signe scout scin 
+ r3 r0 q3 q0 ovr np noe ng i_8 i_7 i_6 i_5 i_4 i_3 i_2 i_1 i_0 fonc d_3 d_2 
+ d_1 d_0 cout cke cin b_3 b_2 b_1 b_0 a_3 a_2 a_1 a_0 
M1 vdde mbk_sig55 signe vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M2 signe mbk_sig55 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M3 vdde mbk_sig55 signe vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M4 signe mbk_sig55 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M5 vdde mbk_sig55 signe vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M6 signe mbk_sig55 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M7 vdde mbk_sig55 signe vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M8 signe mbk_sig55 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M9 vdde mbk_sig55 signe vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M10 signe mbk_sig55 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M11 vdde mbk_sig55 signe vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M12 signe mbk_sig55 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M13 vdde mbk_sig55 signe vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M14 signe mbk_sig55 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M15 vdde mbk_sig55 signe vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M16 signe mbk_sig55 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M17 vdde mbk_sig55 signe vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M18 signe mbk_sig55 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M19 vdde mbk_sig55 signe vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M20 signe mbk_sig55 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M21 vdde mbk_sig55 signe vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M22 signe mbk_sig55 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M23 vdde mbk_sig55 signe vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M24 signe mbk_sig55 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M25 vddi mbk_sig178 mbk_sig55 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M26 mbk_sig55 mbk_sig178 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M27 mbk_sig55 mbk_sig178 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M28 vddi mbk_sig179 mbk_sig178 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M29 vddi mbk_sig178 mbk_sig55 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M30 mbk_sig179 signec vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M31 vdde mbk_sig467 ovr vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M32 ovr mbk_sig467 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M33 vdde mbk_sig467 ovr vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M34 ovr mbk_sig467 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M35 vdde mbk_sig467 ovr vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M36 ovr mbk_sig467 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M37 vdde mbk_sig467 ovr vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M38 ovr mbk_sig467 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M39 vdde mbk_sig467 ovr vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M40 ovr mbk_sig467 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M41 vdde mbk_sig467 ovr vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M42 ovr mbk_sig467 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M43 vdde mbk_sig467 ovr vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M44 ovr mbk_sig467 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M45 vdde mbk_sig467 ovr vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M46 ovr mbk_sig467 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M47 vdde mbk_sig467 ovr vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M48 ovr mbk_sig467 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M49 vdde mbk_sig467 ovr vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M50 ovr mbk_sig467 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M51 vdde mbk_sig467 ovr vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M52 ovr mbk_sig467 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M53 vdde mbk_sig467 ovr vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M54 ovr mbk_sig467 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M55 vddi mbk_sig478 mbk_sig467 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M56 mbk_sig467 mbk_sig478 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M57 mbk_sig467 mbk_sig478 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M58 vddi mbk_sig479 mbk_sig478 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M59 vddi mbk_sig478 mbk_sig467 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M60 mbk_sig479 ovrc vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P PS=22.32U 
+ PD=22.32U 
M61 vdde mbk_sig682 cout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M62 cout mbk_sig682 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M63 vdde mbk_sig682 cout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M64 cout mbk_sig682 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M65 vdde mbk_sig682 cout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M66 cout mbk_sig682 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M67 vdde mbk_sig682 cout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M68 cout mbk_sig682 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M69 vdde mbk_sig682 cout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M70 cout mbk_sig682 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M71 vdde mbk_sig682 cout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M72 cout mbk_sig682 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M73 vdde mbk_sig682 cout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M74 cout mbk_sig682 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M75 vdde mbk_sig682 cout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M76 cout mbk_sig682 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M77 vdde mbk_sig682 cout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M78 cout mbk_sig682 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M79 vdde mbk_sig682 cout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M80 cout mbk_sig682 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M81 vdde mbk_sig682 cout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M82 cout mbk_sig682 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M83 vdde mbk_sig682 cout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M84 cout mbk_sig682 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M85 vddi mbk_sig687 mbk_sig682 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M86 mbk_sig682 mbk_sig687 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M87 mbk_sig682 mbk_sig687 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M88 vddi mbk_sig686 mbk_sig687 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M89 vddi mbk_sig687 mbk_sig682 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M90 mbk_sig686 coutc vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M91 vdde mbk_sig871 zero vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M92 zero mbk_sig871 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M93 vdde mbk_sig871 zero vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M94 zero mbk_sig871 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M95 vdde mbk_sig871 zero vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M96 zero mbk_sig871 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M97 vdde mbk_sig871 zero vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M98 zero mbk_sig871 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M99 vdde mbk_sig871 zero vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M100 zero mbk_sig871 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M101 vdde mbk_sig871 zero vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M102 zero mbk_sig871 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M103 vdde mbk_sig871 zero vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M104 zero mbk_sig871 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M105 vdde mbk_sig871 zero vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M106 zero mbk_sig871 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M107 vdde mbk_sig871 zero vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M108 zero mbk_sig871 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M109 vdde mbk_sig871 zero vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M110 zero mbk_sig871 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M111 vdde mbk_sig871 zero vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M112 zero mbk_sig871 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M113 vdde mbk_sig871 zero vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M114 zero mbk_sig871 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M115 vddi mbk_sig878 mbk_sig871 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M116 mbk_sig871 mbk_sig878 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M117 mbk_sig871 mbk_sig878 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M118 vddi mbk_sig879 mbk_sig878 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M119 vddi mbk_sig878 mbk_sig871 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M120 mbk_sig879 zeroc vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M121 fonc vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M122 vdde vdde fonc vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M123 fonc vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M124 vdde vdde fonc vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M125 vddi fonc mbk_sig1066 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M126 fonci mbk_sig1066 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M127 vddi mbk_sig1066 fonci vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M128 test vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M129 vdde vdde test vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M130 test vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M131 vdde vdde test vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M132 vddi test mbk_sig1271 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M133 testi mbk_sig1271 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M134 vddi mbk_sig1271 testi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M135 scin vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M136 vdde vdde scin vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M137 scin vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M138 vdde vdde scin vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M139 vddi scin mbk_sig1466 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M140 scini mbk_sig1466 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M141 vddi mbk_sig1466 scini vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M142 q0 mbk_sig1638 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M143 vdde mbk_sig1638 q0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M144 q0 mbk_sig1638 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M145 vdde mbk_sig1638 q0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M146 vdde mbk_sig1638 q0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M147 q0 mbk_sig1638 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M148 vdde mbk_sig1638 q0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M149 q0 mbk_sig1638 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M150 vdde mbk_sig1638 q0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M151 q0 mbk_sig1638 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M152 vdde mbk_sig1638 q0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M153 q0 mbk_sig1638 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M154 vdde mbk_sig1638 q0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M155 q0 mbk_sig1638 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M156 vdde mbk_sig1638 q0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M157 q0 mbk_sig1638 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M158 vdde mbk_sig1638 q0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M159 q0 mbk_sig1638 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M160 vdde mbk_sig1638 q0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M161 q0 mbk_sig1638 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M162 vdde mbk_sig1638 q0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M163 q0 mbk_sig1638 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M164 vdde mbk_sig1638 q0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M165 q0 mbk_sig1638 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M166 mbk_sig1652 decaldc vddi vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
M167 vddi mbk_sig1652 mbk_sig1653 vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
M168 q0i mbk_sig1636 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M169 vddi q0 mbk_sig1636 vddi TP L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M170 vddi vssi q0 vddi TP L=7.2U W=0.54U AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
+ 
M171 vddi mbk_sig1653 mbk_sig1638 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M172 mbk_sig1647 f0c vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M173 vddi mbk_sig1636 q0i vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M174 mbk_sig1638 mbk_sig1653 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M175 vddi mbk_sig1653 mbk_sig1638 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M176 mbk_sig1638 mbk_sig1653 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M177 vddi mbk_sig1647 mbk_sig1646 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M178 mbk_sig1638 mbk_sig1646 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M179 vddi mbk_sig1646 mbk_sig1638 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M180 vddi mbk_sig1646 mbk_sig1638 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M181 mbk_sig1638 mbk_sig1652 mbk_sig1639 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M182 mbk_sig1639 mbk_sig1652 mbk_sig1638 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M183 mbk_sig1638 mbk_sig1646 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M184 mbk_sig1638 mbk_sig1652 mbk_sig1639 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M185 mbk_sig1639 mbk_sig1652 mbk_sig1638 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M186 q3 mbk_sig1817 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M187 vdde mbk_sig1817 q3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M188 q3 mbk_sig1817 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M189 vdde mbk_sig1817 q3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M190 vdde mbk_sig1817 q3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M191 q3 mbk_sig1817 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M192 vdde mbk_sig1817 q3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M193 q3 mbk_sig1817 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M194 vdde mbk_sig1817 q3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M195 q3 mbk_sig1817 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M196 vdde mbk_sig1817 q3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M197 q3 mbk_sig1817 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M198 vdde mbk_sig1817 q3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M199 q3 mbk_sig1817 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M200 vdde mbk_sig1817 q3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M201 q3 mbk_sig1817 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M202 vdde mbk_sig1817 q3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M203 q3 mbk_sig1817 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M204 vdde mbk_sig1817 q3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M205 q3 mbk_sig1817 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M206 vdde mbk_sig1817 q3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M207 q3 mbk_sig1817 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M208 vdde mbk_sig1817 q3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M209 q3 mbk_sig1817 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M210 mbk_sig1835 decalgc vddi vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
M211 vddi mbk_sig1835 mbk_sig1836 vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
M212 q3i mbk_sig1815 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M213 vddi q3 mbk_sig1815 vddi TP L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M214 vddi vssi q3 vddi TP L=7.2U W=0.54U AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
+ 
M215 vddi mbk_sig1836 mbk_sig1817 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M216 mbk_sig1827 f3c vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M217 vddi mbk_sig1815 q3i vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M218 mbk_sig1817 mbk_sig1836 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M219 vddi mbk_sig1836 mbk_sig1817 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M220 mbk_sig1817 mbk_sig1836 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M221 vddi mbk_sig1827 mbk_sig1826 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M222 mbk_sig1817 mbk_sig1826 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M223 vddi mbk_sig1826 mbk_sig1817 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M224 vddi mbk_sig1826 mbk_sig1817 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M225 mbk_sig1817 mbk_sig1835 mbk_sig1818 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M226 mbk_sig1818 mbk_sig1835 mbk_sig1817 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M227 mbk_sig1817 mbk_sig1826 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M228 mbk_sig1817 mbk_sig1835 mbk_sig1818 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M229 mbk_sig1818 mbk_sig1835 mbk_sig1817 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M230 cin vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M231 vdde vdde cin vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M232 cin vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M233 vdde vdde cin vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M234 vddi cin mbk_sig44 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M235 cini mbk_sig44 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M236 vddi mbk_sig44 cini vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M237 vdde mbk_sig57 np vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M238 np mbk_sig57 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M239 vdde mbk_sig57 np vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M240 np mbk_sig57 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M241 vdde mbk_sig57 np vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M242 np mbk_sig57 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M243 vdde mbk_sig57 np vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M244 np mbk_sig57 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M245 vdde mbk_sig57 np vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M246 np mbk_sig57 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M247 vdde mbk_sig57 np vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M248 np mbk_sig57 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M249 vdde mbk_sig57 np vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M250 np mbk_sig57 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M251 vdde mbk_sig57 np vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M252 np mbk_sig57 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M253 vdde mbk_sig57 np vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M254 np mbk_sig57 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M255 vdde mbk_sig57 np vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M256 np mbk_sig57 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M257 vdde mbk_sig57 np vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M258 np mbk_sig57 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M259 vdde mbk_sig57 np vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M260 np mbk_sig57 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M261 vddi mbk_sig265 mbk_sig57 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M262 mbk_sig57 mbk_sig265 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M263 mbk_sig57 mbk_sig265 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M264 vddi mbk_sig180 mbk_sig265 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M265 vddi mbk_sig265 mbk_sig57 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M266 mbk_sig180 npc vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P PS=22.32U 
+ PD=22.32U 
M267 vdde mbk_sig469 ng vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M268 ng mbk_sig469 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M269 vdde mbk_sig469 ng vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M270 ng mbk_sig469 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M271 vdde mbk_sig469 ng vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M272 ng mbk_sig469 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M273 vdde mbk_sig469 ng vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M274 ng mbk_sig469 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M275 vdde mbk_sig469 ng vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M276 ng mbk_sig469 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M277 vdde mbk_sig469 ng vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M278 ng mbk_sig469 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M279 vdde mbk_sig469 ng vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M280 ng mbk_sig469 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M281 vdde mbk_sig469 ng vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M282 ng mbk_sig469 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M283 vdde mbk_sig469 ng vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M284 ng mbk_sig469 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M285 vdde mbk_sig469 ng vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M286 ng mbk_sig469 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M287 vdde mbk_sig469 ng vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M288 ng mbk_sig469 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M289 vdde mbk_sig469 ng vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M290 ng mbk_sig469 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M291 vddi mbk_sig480 mbk_sig469 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M292 mbk_sig469 mbk_sig480 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M293 mbk_sig469 mbk_sig480 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M294 vddi mbk_sig481 mbk_sig480 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M295 vddi mbk_sig480 mbk_sig469 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M296 mbk_sig481 ngc vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P PS=22.32U 
+ PD=22.32U 
M297 r0 mbk_sig670 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M298 vdde mbk_sig670 r0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M299 r0 mbk_sig670 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M300 vdde mbk_sig670 r0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M301 vdde mbk_sig670 r0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M302 r0 mbk_sig670 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M303 vdde mbk_sig670 r0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M304 r0 mbk_sig670 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M305 vdde mbk_sig670 r0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M306 r0 mbk_sig670 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M307 vdde mbk_sig670 r0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M308 r0 mbk_sig670 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M309 vdde mbk_sig670 r0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M310 r0 mbk_sig670 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M311 vdde mbk_sig670 r0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M312 r0 mbk_sig670 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M313 vdde mbk_sig670 r0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M314 r0 mbk_sig670 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M315 vdde mbk_sig670 r0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M316 r0 mbk_sig670 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M317 vdde mbk_sig670 r0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M318 r0 mbk_sig670 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M319 vdde mbk_sig670 r0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M320 r0 mbk_sig670 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M321 mbk_sig690 decaldrc vddi vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
M322 vddi mbk_sig690 mbk_sig689 vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
M323 r0i mbk_sig671 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P PS=22.32U 
+ PD=22.32U 
M324 vddi r0 mbk_sig671 vddi TP L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M325 vddi vssi r0 vddi TP L=7.2U W=0.54U AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
+ 
M326 vddi mbk_sig689 mbk_sig670 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M327 mbk_sig683 s0c vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P PS=22.32U 
+ PD=22.32U 
M328 vddi mbk_sig671 r0i vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P PS=22.32U 
+ PD=22.32U 
M329 mbk_sig670 mbk_sig689 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M330 vddi mbk_sig689 mbk_sig670 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M331 mbk_sig670 mbk_sig689 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M332 vddi mbk_sig683 mbk_sig688 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M333 mbk_sig670 mbk_sig688 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M334 vddi mbk_sig688 mbk_sig670 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M335 vddi mbk_sig688 mbk_sig670 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M336 mbk_sig670 mbk_sig690 mbk_sig669 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M337 mbk_sig669 mbk_sig690 mbk_sig670 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M338 mbk_sig670 mbk_sig688 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M339 mbk_sig670 mbk_sig690 mbk_sig669 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M340 mbk_sig669 mbk_sig690 mbk_sig670 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M341 r3 mbk_sig874 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M342 vdde mbk_sig874 r3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M343 r3 mbk_sig874 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M344 vdde mbk_sig874 r3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M345 vdde mbk_sig874 r3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M346 r3 mbk_sig874 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M347 vdde mbk_sig874 r3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M348 r3 mbk_sig874 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M349 vdde mbk_sig874 r3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M350 r3 mbk_sig874 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M351 vdde mbk_sig874 r3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M352 r3 mbk_sig874 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M353 vdde mbk_sig874 r3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M354 r3 mbk_sig874 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M355 vdde mbk_sig874 r3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M356 r3 mbk_sig874 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M357 vdde mbk_sig874 r3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M358 r3 mbk_sig874 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M359 vdde mbk_sig874 r3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M360 r3 mbk_sig874 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M361 vdde mbk_sig874 r3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M362 r3 mbk_sig874 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M363 vdde mbk_sig874 r3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M364 r3 mbk_sig874 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M365 mbk_sig885 decalgrc vddi vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
M366 vddi mbk_sig885 mbk_sig884 vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
M367 r3i mbk_sig876 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P PS=22.32U 
+ PD=22.32U 
M368 vddi r3 mbk_sig876 vddi TP L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M369 vddi vssi r3 vddi TP L=7.2U W=0.54U AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
+ 
M370 vddi mbk_sig884 mbk_sig874 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M371 mbk_sig881 s3c vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P PS=22.32U 
+ PD=22.32U 
M372 vddi mbk_sig876 r3i vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P PS=22.32U 
+ PD=22.32U 
M373 mbk_sig874 mbk_sig884 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M374 vddi mbk_sig884 mbk_sig874 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M375 mbk_sig874 mbk_sig884 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M376 vddi mbk_sig881 mbk_sig880 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M377 mbk_sig874 mbk_sig880 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M378 vddi mbk_sig880 mbk_sig874 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M379 vddi mbk_sig880 mbk_sig874 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M380 mbk_sig874 mbk_sig885 mbk_sig873 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M381 mbk_sig873 mbk_sig885 mbk_sig874 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M382 mbk_sig874 mbk_sig880 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M383 mbk_sig874 mbk_sig885 mbk_sig873 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M384 mbk_sig873 mbk_sig885 mbk_sig874 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M385 y_0 mbk_sig1076 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M386 vdde mbk_sig1076 y_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M387 y_0 mbk_sig1076 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M388 vdde mbk_sig1076 y_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M389 vdde mbk_sig1076 y_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M390 y_0 mbk_sig1076 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M391 vdde mbk_sig1076 y_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M392 y_0 mbk_sig1076 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M393 vdde mbk_sig1076 y_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M394 y_0 mbk_sig1076 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M395 vdde mbk_sig1076 y_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M396 y_0 mbk_sig1076 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M397 vdde mbk_sig1076 y_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M398 y_0 mbk_sig1076 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M399 vdde mbk_sig1076 y_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M400 y_0 mbk_sig1076 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M401 vdde mbk_sig1076 y_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M402 y_0 mbk_sig1076 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M403 vdde mbk_sig1076 y_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M404 y_0 mbk_sig1076 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M405 vdde mbk_sig1076 y_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M406 y_0 mbk_sig1076 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M407 vdde mbk_sig1076 y_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M408 y_0 mbk_sig1076 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M409 mbk_sig1076 mbk_sig1224 mbk_sig1075 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M410 mbk_sig1075 mbk_sig1224 mbk_sig1076 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M411 mbk_sig1076 mbk_sig1224 mbk_sig1075 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M412 mbk_sig1075 mbk_sig1224 mbk_sig1076 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M413 mbk_sig1076 mbk_sig1084 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M414 vddi mbk_sig1084 mbk_sig1076 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M415 vddi mbk_sig1085 mbk_sig1084 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M416 mbk_sig1076 mbk_sig1084 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M417 vddi mbk_sig1084 mbk_sig1076 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M418 mbk_sig1076 mbk_sig1223 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M419 vddi mbk_sig1223 mbk_sig1076 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M420 mbk_sig1076 mbk_sig1223 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M421 vddi mbk_sig1223 mbk_sig1076 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M422 mbk_sig1085 yc_0 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M423 mbk_sig1224 oec vddi vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
M424 vddi mbk_sig1224 mbk_sig1223 vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
M425 vddi vssi y_0 vddi TP L=7.2U W=0.54U AS=0.1944P AD=0.1944P PS=1.8U 
+ PD=1.8U 
M426 y_1 mbk_sig1248 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M427 vdde mbk_sig1248 y_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M428 y_1 mbk_sig1248 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M429 vdde mbk_sig1248 y_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M430 vdde mbk_sig1248 y_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M431 y_1 mbk_sig1248 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M432 vdde mbk_sig1248 y_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M433 y_1 mbk_sig1248 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M434 vdde mbk_sig1248 y_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M435 y_1 mbk_sig1248 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M436 vdde mbk_sig1248 y_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M437 y_1 mbk_sig1248 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M438 vdde mbk_sig1248 y_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M439 y_1 mbk_sig1248 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M440 vdde mbk_sig1248 y_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M441 y_1 mbk_sig1248 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M442 vdde mbk_sig1248 y_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M443 y_1 mbk_sig1248 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M444 vdde mbk_sig1248 y_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M445 y_1 mbk_sig1248 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M446 vdde mbk_sig1248 y_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M447 y_1 mbk_sig1248 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M448 vdde mbk_sig1248 y_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M449 y_1 mbk_sig1248 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M450 mbk_sig1248 mbk_sig1261 mbk_sig1247 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M451 mbk_sig1247 mbk_sig1261 mbk_sig1248 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M452 mbk_sig1248 mbk_sig1261 mbk_sig1247 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M453 mbk_sig1247 mbk_sig1261 mbk_sig1248 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M454 mbk_sig1248 mbk_sig1251 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M455 vddi mbk_sig1251 mbk_sig1248 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M456 vddi mbk_sig1250 mbk_sig1251 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M457 mbk_sig1248 mbk_sig1251 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M458 vddi mbk_sig1251 mbk_sig1248 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M459 mbk_sig1248 mbk_sig1260 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M460 vddi mbk_sig1260 mbk_sig1248 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M461 mbk_sig1248 mbk_sig1260 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M462 vddi mbk_sig1260 mbk_sig1248 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M463 mbk_sig1250 yc_1 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M464 mbk_sig1261 oec vddi vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
M465 vddi mbk_sig1261 mbk_sig1260 vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
M466 vddi vssi y_1 vddi TP L=7.2U W=0.54U AS=0.1944P AD=0.1944P PS=1.8U 
+ PD=1.8U 
M467 y_2 mbk_sig1449 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M468 vdde mbk_sig1449 y_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M469 y_2 mbk_sig1449 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M470 vdde mbk_sig1449 y_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M471 vdde mbk_sig1449 y_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M472 y_2 mbk_sig1449 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M473 vdde mbk_sig1449 y_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M474 y_2 mbk_sig1449 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M475 vdde mbk_sig1449 y_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M476 y_2 mbk_sig1449 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M477 vdde mbk_sig1449 y_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M478 y_2 mbk_sig1449 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M479 vdde mbk_sig1449 y_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M480 y_2 mbk_sig1449 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M481 vdde mbk_sig1449 y_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M482 y_2 mbk_sig1449 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M483 vdde mbk_sig1449 y_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M484 y_2 mbk_sig1449 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M485 vdde mbk_sig1449 y_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M486 y_2 mbk_sig1449 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M487 vdde mbk_sig1449 y_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M488 y_2 mbk_sig1449 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M489 vdde mbk_sig1449 y_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M490 y_2 mbk_sig1449 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M491 mbk_sig1449 mbk_sig1459 mbk_sig1448 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M492 mbk_sig1448 mbk_sig1459 mbk_sig1449 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M493 mbk_sig1449 mbk_sig1459 mbk_sig1448 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M494 mbk_sig1448 mbk_sig1459 mbk_sig1449 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M495 mbk_sig1449 mbk_sig1454 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M496 vddi mbk_sig1454 mbk_sig1449 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M497 vddi mbk_sig1450 mbk_sig1454 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M498 mbk_sig1449 mbk_sig1454 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M499 vddi mbk_sig1454 mbk_sig1449 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M500 mbk_sig1449 mbk_sig1458 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M501 vddi mbk_sig1458 mbk_sig1449 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M502 mbk_sig1449 mbk_sig1458 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M503 vddi mbk_sig1458 mbk_sig1449 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M504 mbk_sig1450 yc_2 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M505 mbk_sig1459 oec vddi vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
M506 vddi mbk_sig1459 mbk_sig1458 vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
M507 vddi vssi y_2 vddi TP L=7.2U W=0.54U AS=0.1944P AD=0.1944P PS=1.8U 
+ PD=1.8U 
M508 y_3 mbk_sig1633 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M509 vdde mbk_sig1633 y_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M510 y_3 mbk_sig1633 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M511 vdde mbk_sig1633 y_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M512 vdde mbk_sig1633 y_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M513 y_3 mbk_sig1633 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M514 vdde mbk_sig1633 y_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M515 y_3 mbk_sig1633 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M516 vdde mbk_sig1633 y_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M517 y_3 mbk_sig1633 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M518 vdde mbk_sig1633 y_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M519 y_3 mbk_sig1633 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M520 vdde mbk_sig1633 y_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M521 y_3 mbk_sig1633 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M522 vdde mbk_sig1633 y_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M523 y_3 mbk_sig1633 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M524 vdde mbk_sig1633 y_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M525 y_3 mbk_sig1633 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M526 vdde mbk_sig1633 y_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M527 y_3 mbk_sig1633 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M528 vdde mbk_sig1633 y_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M529 y_3 mbk_sig1633 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M530 vdde mbk_sig1633 y_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M531 y_3 mbk_sig1633 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M532 mbk_sig1633 mbk_sig1641 mbk_sig1632 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M533 mbk_sig1632 mbk_sig1641 mbk_sig1633 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M534 mbk_sig1633 mbk_sig1641 mbk_sig1632 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M535 mbk_sig1632 mbk_sig1641 mbk_sig1633 vddi TP L=0.18U W=10.62U AS=3.8232P 
+ AD=3.8232P PS=21.96U PD=21.96U 
M536 mbk_sig1633 mbk_sig1634 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M537 vddi mbk_sig1634 mbk_sig1633 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M538 vddi mbk_sig1635 mbk_sig1634 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M539 mbk_sig1633 mbk_sig1634 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M540 vddi mbk_sig1634 mbk_sig1633 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M541 mbk_sig1633 mbk_sig1640 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M542 vddi mbk_sig1640 mbk_sig1633 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M543 mbk_sig1633 mbk_sig1640 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M544 vddi mbk_sig1640 mbk_sig1633 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M545 mbk_sig1635 yc_3 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M546 mbk_sig1641 oec vddi vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
M547 vddi mbk_sig1641 mbk_sig1640 vddi TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
M548 vddi vssi y_3 vddi TP L=7.2U W=0.54U AS=0.1944P AD=0.1944P PS=1.8U 
+ PD=1.8U 
M549 noe vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M550 vdde vdde noe vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M551 noe vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M552 vdde vdde noe vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M553 vddi noe mbk_sig1975 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M554 noei mbk_sig1975 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M555 vddi mbk_sig1975 noei vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M556 vdde mbk_sig13 scout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M557 scout mbk_sig13 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M558 vdde mbk_sig13 scout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M559 scout mbk_sig13 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M560 vdde mbk_sig13 scout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M561 scout mbk_sig13 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M562 vdde mbk_sig13 scout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M563 scout mbk_sig13 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M564 vdde mbk_sig13 scout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M565 scout mbk_sig13 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M566 vdde mbk_sig13 scout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M567 scout mbk_sig13 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M568 vdde mbk_sig13 scout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M569 scout mbk_sig13 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M570 vdde mbk_sig13 scout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M571 scout mbk_sig13 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M572 vdde mbk_sig13 scout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M573 scout mbk_sig13 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M574 vdde mbk_sig13 scout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M575 scout mbk_sig13 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M576 vdde mbk_sig13 scout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M577 scout mbk_sig13 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M578 vdde mbk_sig13 scout vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M579 scout mbk_sig13 vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P 
+ PS=29.52U PD=29.52U 
M580 vddi mbk_sig16 mbk_sig13 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M581 mbk_sig13 mbk_sig16 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M582 mbk_sig13 mbk_sig16 vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M583 vddi mbk_sig17 mbk_sig16 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M584 vddi mbk_sig16 mbk_sig13 vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M585 mbk_sig17 scoutc vddi vddi TP L=0.18U W=10.8U AS=3.888P AD=3.888P 
+ PS=22.32U PD=22.32U 
M586 i_8 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M587 vdde vdde i_8 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M588 i_8 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M589 vdde vdde i_8 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M590 vddi i_8 mbk_sig20 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M591 ii_8 mbk_sig20 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M592 vddi mbk_sig20 ii_8 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M593 i_7 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M594 vdde vdde i_7 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M595 i_7 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M596 vdde vdde i_7 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M597 vddi i_7 mbk_sig22 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M598 ii_7 mbk_sig22 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M599 vddi mbk_sig22 ii_7 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M600 i_6 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M601 vdde vdde i_6 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M602 i_6 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M603 vdde vdde i_6 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M604 vddi i_6 mbk_sig24 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M605 ii_6 mbk_sig24 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M606 vddi mbk_sig24 ii_6 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M607 cko mbk_sig40 vddi vddi TP L=0.18U W=6.12U AS=2.2032P AD=2.2032P 
+ PS=12.96U PD=12.96U 
M608 vddi mbk_sig40 cko vddi TP L=0.18U W=6.12U AS=2.2032P AD=2.2032P 
+ PS=12.96U PD=12.96U 
M609 cko mbk_sig40 vddi vddi TP L=0.18U W=6.12U AS=2.2032P AD=2.2032P 
+ PS=12.96U PD=12.96U 
M610 vddi mbk_sig40 cko vddi TP L=0.18U W=6.12U AS=2.2032P AD=2.2032P 
+ PS=12.96U PD=12.96U 
M611 cko mbk_sig40 vddi vddi TP L=0.18U W=6.12U AS=2.2032P AD=2.2032P 
+ PS=12.96U PD=12.96U 
M612 mbk_sig40 ck_log_log_ck vddi vddi TP L=0.18U W=7.2U AS=2.592P AD=2.592P 
+ PS=15.12U PD=15.12U 
M613 i_5 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M614 vdde vdde i_5 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M615 i_5 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M616 vdde vdde i_5 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M617 vddi i_5 mbk_sig26 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M618 ii_5 mbk_sig26 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M619 vddi mbk_sig26 ii_5 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M620 i_4 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M621 vdde vdde i_4 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M622 i_4 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M623 vdde vdde i_4 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M624 vddi i_4 mbk_sig28 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M625 ii_4 mbk_sig28 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M626 vddi mbk_sig28 ii_4 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M627 i_3 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M628 vdde vdde i_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M629 i_3 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M630 vdde vdde i_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M631 vddi i_3 mbk_sig30 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M632 ii_3 mbk_sig30 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M633 vddi mbk_sig30 ii_3 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M634 i_2 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M635 vdde vdde i_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M636 i_2 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M637 vdde vdde i_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M638 vddi i_2 mbk_sig32 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M639 ii_2 mbk_sig32 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M640 vddi mbk_sig32 ii_2 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M641 i_1 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M642 vdde vdde i_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M643 i_1 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M644 vdde vdde i_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M645 vddi i_1 mbk_sig34 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M646 ii_1 mbk_sig34 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M647 vddi mbk_sig34 ii_1 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M648 i_0 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M649 vdde vdde i_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M650 i_0 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M651 vdde vdde i_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M652 vddi i_0 mbk_sig36 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M653 ii_0 mbk_sig36 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M654 vddi mbk_sig36 ii_0 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M655 vdde vdde cke vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M656 cke vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M657 vdde vdde cke vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M658 cke vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M659 ck_log_log_ck mbk_sig38 vddi vddi TP L=0.18U W=10.26U AS=3.6936P 
+ AD=3.6936P PS=21.24U PD=21.24U 
M660 vddi mbk_sig38 ck_log_log_ck vddi TP L=0.18U W=10.26U AS=3.6936P 
+ AD=3.6936P PS=21.24U PD=21.24U 
M661 ck_log_log_ck mbk_sig38 vddi vddi TP L=0.18U W=10.26U AS=3.6936P 
+ AD=3.6936P PS=21.24U PD=21.24U 
M662 ck_log_log_ck mbk_sig38 vddi vddi TP L=0.18U W=10.26U AS=3.6936P 
+ AD=3.6936P PS=21.24U PD=21.24U 
M663 vddi mbk_sig38 ck_log_log_ck vddi TP L=0.18U W=10.26U AS=3.6936P 
+ AD=3.6936P PS=21.24U PD=21.24U 
M664 ck_log_log_ck mbk_sig38 vddi vddi TP L=0.18U W=10.26U AS=3.6936P 
+ AD=3.6936P PS=21.24U PD=21.24U 
M665 vddi mbk_sig38 ck_log_log_ck vddi TP L=0.18U W=10.26U AS=3.6936P 
+ AD=3.6936P PS=21.24U PD=21.24U 
M666 vddi mbk_sig38 ck_log_log_ck vddi TP L=0.18U W=10.26U AS=3.6936P 
+ AD=3.6936P PS=21.24U PD=21.24U 
M667 vddi cke mbk_sig38 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M668 mbk_sig38 cke vddi vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M669 vddi cke mbk_sig38 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M670 mbk_sig38 cke vddi vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M671 a_3 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M672 vdde vdde a_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M673 a_3 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M674 vdde vdde a_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M675 vddi a_3 mbk_sig1976 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M676 heart_a_3 mbk_sig1976 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M677 vddi mbk_sig1976 heart_a_3 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M678 a_2 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M679 vdde vdde a_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M680 a_2 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M681 vdde vdde a_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M682 vddi a_2 mbk_sig1977 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M683 heart_a_2 mbk_sig1977 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M684 vddi mbk_sig1977 heart_a_2 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M685 a_1 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M686 vdde vdde a_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M687 a_1 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M688 vdde vdde a_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M689 vddi a_1 mbk_sig1978 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M690 heart_a_1 mbk_sig1978 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M691 vddi mbk_sig1978 heart_a_1 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M692 a_0 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M693 vdde vdde a_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M694 a_0 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M695 vdde vdde a_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M696 vddi a_0 mbk_sig1979 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M697 heart_a_0 mbk_sig1979 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M698 vddi mbk_sig1979 heart_a_0 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M699 b_3 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M700 vdde vdde b_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M701 b_3 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M702 vdde vdde b_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M703 vddi b_3 mbk_sig1980 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M704 heart_b_3 mbk_sig1980 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M705 vddi mbk_sig1980 heart_b_3 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M706 b_2 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M707 vdde vdde b_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M708 b_2 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M709 vdde vdde b_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M710 vddi b_2 mbk_sig1981 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M711 heart_b_2 mbk_sig1981 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M712 vddi mbk_sig1981 heart_b_2 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M713 b_1 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M714 vdde vdde b_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M715 b_1 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M716 vdde vdde b_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M717 vddi b_1 mbk_sig1982 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M718 heart_b_1 mbk_sig1982 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M719 vddi mbk_sig1982 heart_b_1 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M720 b_0 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M721 vdde vdde b_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M722 b_0 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M723 vdde vdde b_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M724 vddi b_0 mbk_sig1983 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M725 heart_b_0 mbk_sig1983 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M726 vddi mbk_sig1983 heart_b_0 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M727 d_3 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M728 vdde vdde d_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M729 d_3 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M730 vdde vdde d_3 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M731 vddi d_3 mbk_sig1984 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M732 heart_d_3 mbk_sig1984 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M733 vddi mbk_sig1984 heart_d_3 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M734 d_2 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M735 vdde vdde d_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M736 d_2 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M737 vdde vdde d_2 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M738 vddi d_2 mbk_sig1985 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M739 heart_d_2 mbk_sig1985 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M740 vddi mbk_sig1985 heart_d_2 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M741 d_1 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M742 vdde vdde d_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M743 d_1 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M744 vdde vdde d_1 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M745 vddi d_1 mbk_sig1986 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M746 heart_d_1 mbk_sig1986 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M747 vddi mbk_sig1986 heart_d_1 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M748 d_0 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M749 vdde vdde d_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M750 d_0 vdde vdde vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M751 vdde vdde d_0 vddi TP L=0.18U W=14.4U AS=5.184P AD=5.184P PS=29.52U 
+ PD=29.52U 
M752 vddi d_0 mbk_sig1987 vddi TP L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M753 heart_d_0 mbk_sig1987 vddi vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M754 vddi mbk_sig1987 heart_d_0 vddi TP L=0.18U W=10.26U AS=3.6936P AD=3.6936P 
+ PS=21.24U PD=21.24U 
M755 mbk_sig1972 heart_block3_pb1 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M756 heart_block3_no31 heart_block3_n3 mbk_sig1972 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M757 mbk_sig1971 heart_block3_no21 mbk_sig1967 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M758 vddi heart_block3_no31 mbk_sig1971 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M759 vddi heart_block3_no31 mbk_sig1970 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M760 mbk_sig1970 heart_block3_no21 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M761 heart_block3_x21 mbk_sig1967 mbk_sig1970 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M762 mbk_sig1968 heart_block3_gb1 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M763 heart_block3_no21 heart_block3_n2 mbk_sig1968 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M764 mbk_sig1966 heart_block4_a29s vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M765 mbk_sig1965 heart_block4_a213s mbk_sig1966 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M766 vddi mbk_sig1965 heart_block4_insh1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M767 mbk_sig1962 heart_block3_x21 mbk_sig1961 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M768 vddi heart_block3_no41 mbk_sig1962 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M769 vddi heart_block3_no41 mbk_sig1964 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M770 mbk_sig1964 heart_block3_x21 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M771 heart_block3_fb1 mbk_sig1961 mbk_sig1964 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M772 heart_block3_na0_csb heart_block3_fb1 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M773 vddi heart_block3_fb0 heart_block3_na0_csb vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M774 vddi heart_block4_decalga mbk_sig1959 vddi TP L=0.18U W=2.7U AS=0.972P 
+ AD=0.972P PS=6.12U PD=6.12U 
M775 vddi mbk_sig1959 decalgc vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M776 decalgc mbk_sig1959 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M777 vddi mbk_sig1958 heart_block4_a221s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M778 vddi heart_block4_insh1 mbk_sig1958 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M779 mbk_sig1958 heart_block4_decalga vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M780 vddi mbk_sig1955 heart_block4_a29s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M781 vddi heart_block2_a26ms_i0 mbk_sig1955 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M782 mbk_sig1955 heart_block4_selalu vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M783 vddi heart_block3_fb1 heart_block2_a26ms_i0 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M784 vddi mbk_sig1953 heart_block4_a28s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M785 vddi heart_block2_a27ms_i0 mbk_sig1953 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M786 mbk_sig1953 heart_block4_selalu vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M787 vddi mbk_sig1952 heart_block4_a212s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M788 vddi heart_q_2 mbk_sig1952 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M789 mbk_sig1952 ii_8 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M790 vddi mbk_sig1949 heart_block4_a219s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M791 vddi heart_block4_insh3 mbk_sig1949 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M792 mbk_sig1949 heart_block4_decalda vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M793 mbk_sig1948 heart_block4_a220s mbk_sig1947 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M794 mbk_sig1946 heart_block4_a221s mbk_sig1948 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M795 vddi mbk_sig1946 heart_block4_shacc2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M796 mbk_sig1947 heart_block4_a219s vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M797 vddi mbk_sig1945 heart_block4_a220s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M798 vddi heart_block4_insh2 mbk_sig1945 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M799 mbk_sig1945 heart_block4_decaln vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M800 mbk_sig1944 heart_block4_a28s vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M801 mbk_sig1942 heart_block4_a212s mbk_sig1944 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M802 vddi mbk_sig1942 heart_block4_insh2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M803 vddi mbk_sig1940 heart_block4_a223s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M804 vddi heart_block4_insh1 mbk_sig1940 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M805 mbk_sig1940 heart_block4_decaln vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M806 vddi mbk_sig1939 heart_block4_a227s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M807 vddi q0i mbk_sig1939 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M808 mbk_sig1939 heart_block4_decalga vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M809 vddi ii_8 heart_block4_decaln vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M810 vddi mbk_sig1936 heart_block4_a217s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M811 vddi heart_block4_insh3 mbk_sig1936 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M812 mbk_sig1936 heart_block4_decaln vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M813 vddi mbk_sig1935 f3c vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M814 vddi heart_block4_decalga mbk_sig1935 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M815 mbk_sig1935 heart_block4_insh3 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M816 vddi mbk_sig1933 heart_block4_a225s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M817 vddi heart_block4_insh1 mbk_sig1933 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M818 mbk_sig1933 heart_block4_decalda vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M819 mbk_sig1929 mbk_sig1925 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M820 vddi heart_block5_m_1_2_dff_m mbk_sig1925 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M821 mbk_sig1930 heart_block5_ck1 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M822 heart_block5_m_1_2_dff_s mbk_sig1931 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M823 vddi heart_block5_m_1_2_dff_s mbk_sig1931 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M824 heart_block5_s21 heart_block5_m_1_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M825 heart_block5_m_1_2_dff_m mbk_sig1925 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M826 mbk_sig1927 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M827 vddi heart_b_1 heart_block5_nb1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M828 mbk_sig1924 heart_block4_a226s mbk_sig1923 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M829 mbk_sig1922 heart_block4_a227s mbk_sig1924 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M830 vddi mbk_sig1922 heart_block4_shacc0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M831 mbk_sig1923 heart_block4_a225s vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M832 vddi mbk_sig1921 heart_block4_a224s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M833 vddi heart_block4_insh0 mbk_sig1921 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M834 mbk_sig1921 heart_block4_decalga vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M835 vddi mbk_sig1919 heart_block5_b16 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M836 vddi heart_b_1 mbk_sig1919 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M837 mbk_sig1919 heart_b_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M838 vddi heart_b_3 mbk_sig1919 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M839 mbk_sig1919 heart_b_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M840 vddi mbk_sig1914 heart_block5_b14 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M841 vddi heart_block5_nb1 mbk_sig1914 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M842 mbk_sig1914 heart_b_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M843 vddi heart_b_3 mbk_sig1914 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M844 mbk_sig1914 heart_b_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M845 vddi mbk_sig1911 heart_block4_a226s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M846 vddi heart_block4_insh0 mbk_sig1911 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M847 mbk_sig1911 heart_block4_decaln vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M848 vddi mbk_sig1909 heart_block5_b8 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M849 vddi heart_b_1 mbk_sig1909 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M850 mbk_sig1909 heart_b_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M851 vddi heart_block5_nb3 mbk_sig1909 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M852 mbk_sig1909 heart_b_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M853 vddi mbk_sig1905 heart_block5_b15 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M854 vddi heart_b_1 mbk_sig1905 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M855 mbk_sig1905 heart_b_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M856 vddi heart_b_3 mbk_sig1905 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M857 mbk_sig1905 heart_block5_nb0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M858 vddi mbk_sig1900 heart_block5_b13 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M859 vddi heart_block5_nb1 mbk_sig1900 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M860 mbk_sig1900 heart_b_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M861 vddi heart_b_3 mbk_sig1900 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M862 mbk_sig1900 heart_block5_nb0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M863 vddi mbk_sig1894 heart_block5_b5 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M864 vddi heart_block5_nb1 mbk_sig1894 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M865 mbk_sig1894 heart_b_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M866 vddi heart_block5_nb3 mbk_sig1894 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M867 mbk_sig1894 heart_block5_nb0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M868 vddi mbk_sig1890 heart_block5_b1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M869 vddi heart_block5_nb1 mbk_sig1890 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M870 mbk_sig1890 heart_block5_nb2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M871 vddi heart_block5_nb3 mbk_sig1890 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M872 mbk_sig1890 heart_block5_nb0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M873 heart_block5_b18s heart_block5_s18 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M874 vddi heart_block5_b8 heart_block5_b18s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M875 mbk_sig1887 mbk_sig1883 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M876 vddi heart_block5_m_8_1_dff_m mbk_sig1883 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M877 mbk_sig1885 heart_block5_ck8 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M878 heart_block5_m_8_1_dff_s mbk_sig1888 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M879 vddi heart_block5_m_8_1_dff_s mbk_sig1888 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M880 heart_block5_s18 heart_block5_m_8_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M881 heart_block5_m_8_1_dff_m mbk_sig1883 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M882 mbk_sig1881 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M883 heart_block5_a18s heart_block5_s18 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M884 vddi heart_block5_a8 heart_block5_a18s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M885 vddi mbk_sig1880 heart_block5_b10 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M886 vddi heart_block5_nb1 mbk_sig1880 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M887 mbk_sig1880 heart_block5_nb2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M888 vddi heart_b_3 mbk_sig1880 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M889 mbk_sig1880 heart_b_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M890 vddi mbk_sig1876 heart_block5_ck5 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M891 vddi heart_block5_enable mbk_sig1876 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M892 mbk_sig1876 heart_block5_b5 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M893 vddi mbk_sig1874 heart_block5_ck8 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M894 vddi heart_block5_enable mbk_sig1874 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M895 mbk_sig1874 heart_block5_b8 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M896 mbk_sig1870 mbk_sig1866 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M897 vddi heart_block5_m_8_2_dff_m mbk_sig1866 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M898 mbk_sig1872 heart_block5_ck8 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M899 heart_block5_m_8_2_dff_s mbk_sig1871 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M900 vddi heart_block5_m_8_2_dff_s mbk_sig1871 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M901 heart_block5_s28 heart_block5_m_8_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M902 heart_block5_m_8_2_dff_m mbk_sig1866 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M903 mbk_sig1868 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M904 heart_block5_b38s heart_block5_s38 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M905 vddi heart_block5_b8 heart_block5_b38s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M906 mbk_sig1862 mbk_sig1857 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M907 vddi heart_block5_m_5_1_dff_m mbk_sig1857 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M908 mbk_sig1863 heart_block5_ck5 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M909 heart_block5_m_5_1_dff_s mbk_sig1865 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M910 vddi heart_block5_m_5_1_dff_s mbk_sig1865 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M911 heart_block5_s15 heart_block5_m_5_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M912 heart_block5_m_5_1_dff_m mbk_sig1857 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M913 mbk_sig1860 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M914 heart_block5_b04s heart_block5_s04 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M915 vddi heart_block5_b4 heart_block5_b04s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M916 mbk_sig1852 mbk_sig1854 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M917 vddi heart_block5_m_4_0_dff_m mbk_sig1854 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M918 mbk_sig1853 heart_block5_ck4 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M919 heart_block5_m_4_0_dff_s mbk_sig1856 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M920 vddi heart_block5_m_4_0_dff_s mbk_sig1856 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M921 heart_block5_s04 heart_block5_m_4_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M922 heart_block5_m_4_0_dff_m mbk_sig1854 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M923 mbk_sig1851 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M924 vddi heart_b_0 heart_block5_nb0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M925 mbk_sig1848 mbk_sig1844 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M926 vddi heart_block5_m_8_3_dff_m mbk_sig1844 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M927 mbk_sig1846 heart_block5_ck8 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M928 heart_block5_m_8_3_dff_s mbk_sig1849 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M929 vddi heart_block5_m_8_3_dff_s mbk_sig1849 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M930 heart_block5_s38 heart_block5_m_8_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M931 heart_block5_m_8_3_dff_m mbk_sig1844 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M932 mbk_sig1843 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M933 heart_block5_a33s heart_block5_s33 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M934 vddi heart_block5_a3 heart_block5_a33s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M935 vddi mbk_sig1841 heart_block5_ck2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M936 vddi heart_block5_enable mbk_sig1841 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M937 mbk_sig1841 heart_block5_b2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M938 vddi mbk_sig1838 heart_block5_ck3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M939 vddi heart_block5_enable mbk_sig1838 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M940 mbk_sig1838 heart_block5_b3 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M941 heart_block5_b33s heart_block5_s33 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M942 vddi heart_block5_b3 heart_block5_b33s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M943 vddi heart_block3_pb1 heart_block3_not1 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M944 heart_block3_na21 heart_block3_cout0 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M945 vddi heart_block3_not1 heart_block3_na21 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M946 heart_block3_nn3 heart_block3_ni5 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M947 vddi ii_4 heart_block3_nn3 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M948 heart_block3_nn3 ii_3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M949 heart_block3_cout0 heart_block3_na20 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M950 vddi heart_block3_gb0 heart_block3_cout0 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M951 mbk_sig1811 heart_block3_cout0 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M952 heart_block3_no41 heart_block3_n4 mbk_sig1811 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M953 mbk_sig1810 heart_block3_ni5 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M954 heart_block3_n2 ii_4 mbk_sig1810 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M955 heart_block3_flag1 ii_3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M956 vddi ii_4 heart_block3_flag1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M957 heart_block3_n4 heart_block3_nn3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M958 vddi heart_block3_ni5 heart_block3_n4 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M959 heart_block3_cout1 heart_block3_na21 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M960 vddi heart_block3_gb1 heart_block3_cout1 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M961 vddi mbk_sig1779 heart_block4_a213s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M962 vddi heart_q_1 mbk_sig1779 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M963 mbk_sig1779 ii_8 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M964 heart_block3_na1_csb heart_block3_signea vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M965 vddi heart_block3_fb2 heart_block3_na1_csb vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M966 mbk_sig1808 heart_block3_na1_csb vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M967 zeroc heart_block3_na0_csb mbk_sig1808 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M968 mbk_sig1806 heart_block3_x22 mbk_sig1805 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M969 vddi heart_block3_no42 mbk_sig1806 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M970 vddi heart_block3_no42 mbk_sig1807 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M971 mbk_sig1807 heart_block3_x22 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M972 heart_block3_fb2 mbk_sig1805 mbk_sig1807 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M973 vddi mbk_sig1774 heart_block5_a26sh vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M974 vddi heart_block2_a26ms_i0 mbk_sig1774 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M975 mbk_sig1774 heart_block5_decalgra vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M976 mbk_sig1803 heart_block3_cout1 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M977 heart_block3_no42 heart_block3_n4 mbk_sig1803 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M978 vddi mbk_sig1773 heart_block3_flag vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M979 vddi heart_block3_ni5 mbk_sig1773 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M980 mbk_sig1773 heart_block3_flag1 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M981 mbk_sig1801 mbk_sig1765 mbk_sig1764 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M982 mbk_sig1764 heart_block4_shacc1 mbk_sig1801 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M983 mbk_sig1765 heart_block4_test_mode vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M984 mbk_sig1801 heart_q_0 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M985 vddi heart_block4_test_mode mbk_sig1801 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M986 heart_q_1 heart_block4_m1_dff_s vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M987 vddi heart_block4_m1_dff_s mbk_sig1772 vddi TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M988 heart_block4_m1_dff_s mbk_sig1772 vddi vddi TP L=0.72U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
M989 mbk_sig1770 mbk_sig1769 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M990 vddi heart_block4_m1_dff_m mbk_sig1769 vddi TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M991 heart_block4_m1_dff_m mbk_sig1769 vddi vddi TP L=0.72U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
M992 mbk_sig1768 heart_block4_ckin vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M993 mbk_sig1800 heart_block4_a223s mbk_sig1799 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M994 mbk_sig1762 heart_block4_a224s mbk_sig1800 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M995 vddi mbk_sig1762 heart_block4_shacc1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M996 mbk_sig1799 heart_block4_a222s vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M997 vddi mbk_sig1757 heart_block4_a222s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M998 vddi heart_block4_insh2 mbk_sig1757 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M999 mbk_sig1757 heart_block4_decalda vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1000 mbk_sig1797 heart_block5_a27sh mbk_sig1796 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1001 mbk_sig1756 heart_block5_a28sh mbk_sig1797 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1002 vddi mbk_sig1756 heart_block5_shram2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1003 mbk_sig1796 heart_block5_a26sh vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M1004 vddi mbk_sig1754 heart_block4_a27s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1005 vddi heart_block2_a28ms_i0 mbk_sig1754 vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1006 mbk_sig1754 heart_block4_selalu vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1007 mbk_sig1795 heart_block4_a27s vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M1008 mbk_sig1752 heart_block4_a211s mbk_sig1795 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1009 vddi mbk_sig1752 heart_block4_insh3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1010 vddi heart_b_3 heart_block5_nb3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1011 vddi mbk_sig1751 heart_block4_decalda vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1012 vddi ii_8 mbk_sig1751 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1013 mbk_sig1751 heart_block4_ni7 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1014 mbk_sig1748 mbk_sig1746 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1015 vddi heart_block5_m_1_1_dff_m mbk_sig1746 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1016 mbk_sig1749 heart_block5_ck1 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1017 heart_block5_m_1_1_dff_s mbk_sig1750 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1018 vddi heart_block5_m_1_1_dff_s mbk_sig1750 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1019 heart_block5_s11 heart_block5_m_1_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1020 heart_block5_m_1_1_dff_m mbk_sig1746 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1021 mbk_sig1745 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1022 vddi heart_b_2 heart_block5_nb2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1023 vddi mbk_sig1743 f0c vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1024 vddi heart_block4_decalda mbk_sig1743 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1025 mbk_sig1743 heart_block4_insh0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1026 vddi mbk_sig1739 heart_block5_b6 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1027 vddi heart_block5_nb1 mbk_sig1739 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1028 mbk_sig1739 heart_b_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1029 vddi heart_block5_nb3 mbk_sig1739 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1030 mbk_sig1739 heart_b_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1031 heart_block5_b27s heart_block5_s27 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1032 vddi heart_block5_b7 heart_block5_b27s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1033 vddi mbk_sig1735 heart_block5_b7 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1034 vddi heart_b_1 mbk_sig1735 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1035 mbk_sig1735 heart_b_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1036 vddi heart_block5_nb3 mbk_sig1735 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1037 mbk_sig1735 heart_block5_nb0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1038 heart_block5_b11s heart_block5_s11 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1039 vddi heart_block5_b1 heart_block5_b11s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1040 vddi mbk_sig1728 heart_block5_b4 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1041 vddi heart_b_1 mbk_sig1728 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1042 mbk_sig1728 heart_block5_nb2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1043 vddi heart_block5_nb3 mbk_sig1728 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1044 mbk_sig1728 heart_b_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1045 vddi mbk_sig1724 heart_block5_ob431s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1046 vddi heart_block5_b16s mbk_sig1724 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1047 mbk_sig1724 heart_block5_b17s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1048 vddi heart_block5_b18s mbk_sig1724 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1049 mbk_sig1724 heart_block5_b15s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1050 vddi mbk_sig1721 heart_block5_b2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1051 vddi heart_block5_nb1 mbk_sig1721 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1052 mbk_sig1721 heart_block5_nb2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1053 vddi heart_block5_nb3 mbk_sig1721 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1054 mbk_sig1721 heart_b_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1055 mbk_sig1716 mbk_sig1714 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1056 vddi heart_block5_m_1_0_dff_m mbk_sig1714 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1057 mbk_sig1717 heart_block5_ck1 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1058 heart_block5_m_1_0_dff_s mbk_sig1718 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1059 vddi heart_block5_m_1_0_dff_s mbk_sig1718 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1060 heart_block5_s01 heart_block5_m_1_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1061 heart_block5_m_1_0_dff_m mbk_sig1714 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1062 mbk_sig1713 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1063 heart_block5_b25s heart_block5_s25 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1064 vddi heart_block5_b5 heart_block5_b25s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1065 heart_block5_b17s heart_block5_s17 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1066 vddi heart_block5_b7 heart_block5_b17s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1067 vddi mbk_sig1704 heart_block5_b12 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1068 vddi heart_b_1 mbk_sig1704 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1069 mbk_sig1704 heart_block5_nb2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1070 vddi heart_b_3 mbk_sig1704 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1071 mbk_sig1704 heart_b_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1072 heart_block5_b24s heart_block5_s24 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1073 vddi heart_block5_b4 heart_block5_b24s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1074 heart_block5_a17s heart_block5_s17 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1075 vddi heart_block5_a7 heart_block5_a17s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1076 vddi mbk_sig1698 heart_block5_b3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1077 vddi heart_b_1 mbk_sig1698 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1078 mbk_sig1698 heart_block5_nb2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1079 vddi heart_block5_nb3 mbk_sig1698 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1080 mbk_sig1698 heart_block5_nb0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1081 mbk_sig1694 mbk_sig1692 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1082 vddi heart_block5_m_5_2_dff_m mbk_sig1692 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1083 mbk_sig1695 heart_block5_ck5 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1084 heart_block5_m_5_2_dff_s mbk_sig1696 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1085 vddi heart_block5_m_5_2_dff_s mbk_sig1696 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1086 heart_block5_s25 heart_block5_m_5_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1087 heart_block5_m_5_2_dff_m mbk_sig1692 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1088 mbk_sig1691 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1089 heart_block5_a28s heart_block5_s28 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1090 vddi heart_block5_a8 heart_block5_a28s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1091 heart_block5_a38s heart_block5_s38 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1092 vddi heart_block5_a8 heart_block5_a38s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1093 mbk_sig1685 mbk_sig1683 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1094 vddi heart_block5_m_4_2_dff_m mbk_sig1683 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1095 mbk_sig1680 heart_block5_ck4 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1096 heart_block5_m_4_2_dff_s mbk_sig1686 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1097 vddi heart_block5_m_4_2_dff_s mbk_sig1686 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1098 heart_block5_s24 heart_block5_m_4_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1099 heart_block5_m_4_2_dff_m mbk_sig1683 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1100 mbk_sig1682 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1101 vddi mbk_sig1679 heart_block5_ck1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1102 vddi heart_block5_enable mbk_sig1679 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1103 mbk_sig1679 heart_block5_b1 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1104 heart_block5_a04s heart_block5_s04 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1105 vddi heart_block5_a4 heart_block5_a04s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1106 heart_block5_b31s heart_block5_s31 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1107 vddi heart_block5_b1 heart_block5_b31s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1108 mbk_sig1671 mbk_sig1673 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1109 vddi heart_block5_m_1_3_dff_m mbk_sig1673 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1110 mbk_sig1672 heart_block5_ck1 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1111 heart_block5_m_1_3_dff_s mbk_sig1675 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1112 vddi heart_block5_m_1_3_dff_s mbk_sig1675 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1113 heart_block5_s31 heart_block5_m_1_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1114 heart_block5_m_1_3_dff_m mbk_sig1673 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1115 mbk_sig1666 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1116 vddi mbk_sig1664 heart_block5_ob443s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1117 vddi heart_block5_b32s mbk_sig1664 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1118 mbk_sig1664 heart_block5_b33s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1119 vddi heart_block5_b34s mbk_sig1664 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1120 mbk_sig1664 heart_block5_b31s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1121 mbk_sig1658 mbk_sig1656 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1122 vddi heart_block5_m_3_3_dff_m mbk_sig1656 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1123 mbk_sig1659 heart_block5_ck3 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1124 heart_block5_m_3_3_dff_s mbk_sig1660 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1125 vddi heart_block5_m_3_3_dff_s mbk_sig1660 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1126 heart_block5_s33 heart_block5_m_3_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1127 heart_block5_m_3_3_dff_m mbk_sig1656 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1128 mbk_sig1655 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1129 vddi heart_block3_nn3 heart_block3_n3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1130 mbk_sig1627 heart_block3_x23 mbk_sig1626 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1131 vddi heart_block3_no43 mbk_sig1627 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1132 vddi heart_block3_no43 mbk_sig1629 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1133 mbk_sig1629 heart_block3_x23 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1134 heart_block3_signea mbk_sig1626 mbk_sig1629 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1135 mbk_sig1624 heart_block3_no23 mbk_sig1623 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1136 vddi heart_block3_no33 mbk_sig1624 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1137 vddi heart_block3_no33 mbk_sig1625 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1138 mbk_sig1625 heart_block3_no23 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1139 heart_block3_x23 mbk_sig1623 mbk_sig1625 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1140 heart_block3_na20 cini vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1141 vddi heart_block3_not0 heart_block3_na20 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1142 mbk_sig1619 heart_block3_gb3 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1143 heart_block3_no23 heart_block3_n2 mbk_sig1619 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1144 mbk_sig1618 cini vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1145 heart_block3_no40 heart_block3_n4 mbk_sig1618 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1146 mbk_sig1615 heart_block3_x20 mbk_sig1614 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1147 vddi heart_block3_no40 mbk_sig1615 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1148 vddi heart_block3_no40 mbk_sig1617 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1149 mbk_sig1617 heart_block3_x20 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1150 heart_block3_fb0 mbk_sig1614 mbk_sig1617 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1151 vddi heart_block3_signea heart_block2_a28ms_i0 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1152 vddi heart_block3_signea signec vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1153 mbk_sig1605 mbk_sig1602 mbk_sig1603 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1154 mbk_sig1603 heart_block4_shacc2 mbk_sig1605 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1155 mbk_sig1602 heart_block4_test_mode vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1156 mbk_sig1605 heart_q_1 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1157 vddi heart_block4_test_mode mbk_sig1605 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1158 heart_q_2 heart_block4_m2_dff_s vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1159 vddi heart_block4_m2_dff_s mbk_sig1612 vddi TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M1160 heart_block4_m2_dff_s mbk_sig1612 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1161 mbk_sig1610 mbk_sig1609 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1162 vddi heart_block4_m2_dff_m mbk_sig1609 vddi TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M1163 heart_block4_m2_dff_m mbk_sig1609 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1164 mbk_sig1608 heart_block4_ckin vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1165 vddi mbk_sig1597 heart_block5_a27sh vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1166 vddi heart_block2_a27ms_i0 mbk_sig1597 vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1167 mbk_sig1597 heart_block5_decalnr vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1168 vddi heart_block3_fb0 heart_block2_a25ms_i0 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1169 vddi heart_block3_fb2 heart_block2_a27ms_i0 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1170 mbk_sig1594 mbk_sig1590 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1171 vddi heart_block5_m_3_2_dff_m mbk_sig1590 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1172 mbk_sig1592 heart_block5_ck3 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1173 heart_block5_m_3_2_dff_s mbk_sig1595 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1174 vddi heart_block5_m_3_2_dff_s mbk_sig1595 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1175 heart_block5_s23 heart_block5_m_3_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1176 heart_block5_m_3_2_dff_m mbk_sig1590 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1177 mbk_sig1587 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1178 vddi mbk_sig1588 heart_block4_a210s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1179 vddi heart_block2_a25ms_i0 mbk_sig1588 vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1180 mbk_sig1588 heart_block4_selalu vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1181 vddi mbk_sig1586 s3c vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1182 vddi heart_block5_decalgra mbk_sig1586 vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1183 mbk_sig1586 heart_block2_a28ms_i0 vddi vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1184 vddi mbk_sig1584 heart_block5_a28sh vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1185 vddi heart_block2_a28ms_i0 mbk_sig1584 vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1186 mbk_sig1584 heart_block5_decaldra vddi vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1187 vddi mbk_sig1580 heart_block4_a216s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1188 vddi q3i mbk_sig1580 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1189 mbk_sig1580 heart_block4_decalda vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1190 mbk_sig1577 mbk_sig1573 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1191 vddi heart_block5_m_6_3_dff_m mbk_sig1573 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1192 mbk_sig1578 heart_block5_ck6 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1193 heart_block5_m_6_3_dff_s mbk_sig1579 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1194 vddi heart_block5_m_6_3_dff_s mbk_sig1579 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1195 heart_block5_s36 heart_block5_m_6_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1196 heart_block5_m_6_3_dff_m mbk_sig1573 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1197 mbk_sig1575 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1198 vddi mbk_sig1572 heart_block4_a211s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1199 vddi heart_q_3 mbk_sig1572 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1200 mbk_sig1572 ii_8 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1201 vddi heart_block4_decalda mbk_sig1567 vddi TP L=0.18U W=2.7U AS=0.972P 
+ AD=0.972P PS=6.12U PD=6.12U 
M1202 vddi mbk_sig1567 decaldc vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1203 decaldc mbk_sig1567 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1204 heart_block5_b21s heart_block5_s21 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1205 vddi heart_block5_b1 heart_block5_b21s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1206 heart_block5_b23s heart_block5_s23 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1207 vddi heart_block5_b3 heart_block5_b23s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1208 heart_block5_a21s heart_block5_s21 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1209 vddi heart_block5_a1 heart_block5_a21s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1210 heart_block5_b26s heart_block5_s26 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1211 vddi heart_block5_b6 heart_block5_b26s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1212 vddi mbk_sig1558 heart_block5_ob432s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1213 vddi heart_block5_b26s mbk_sig1558 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1214 mbk_sig1558 heart_block5_b27s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1215 vddi heart_block5_b28s mbk_sig1558 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1216 mbk_sig1558 heart_block5_b25s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1217 vddi mbk_sig1554 heart_block5_ck7 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1218 vddi heart_block5_enable mbk_sig1554 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1219 mbk_sig1554 heart_block5_b7 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1220 vddi mbk_sig1549 heart_block5_ob442s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1221 vddi heart_block5_b22s mbk_sig1549 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1222 mbk_sig1549 heart_block5_b23s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1223 vddi heart_block5_b24s mbk_sig1549 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1224 mbk_sig1549 heart_block5_b21s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1225 vddi mbk_sig1546 heart_block5_b11 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1226 vddi heart_b_1 mbk_sig1546 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1227 mbk_sig1546 heart_block5_nb2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1228 vddi heart_b_3 mbk_sig1546 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1229 mbk_sig1546 heart_block5_nb0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1230 heart_block5_b15s heart_block5_s15 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1231 vddi heart_block5_b5 heart_block5_b15s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1232 mbk_sig1540 mbk_sig1536 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1233 vddi heart_block5_m_7_1_dff_m mbk_sig1536 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1234 mbk_sig1538 heart_block5_ck7 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1235 heart_block5_m_7_1_dff_s mbk_sig1542 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1236 vddi heart_block5_m_7_1_dff_s mbk_sig1542 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1237 heart_block5_s17 heart_block5_m_7_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1238 heart_block5_m_7_1_dff_m mbk_sig1536 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1239 mbk_sig1534 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1240 mbk_sig1532 mbk_sig1526 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1241 vddi heart_block5_m_8_0_dff_m mbk_sig1526 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1242 mbk_sig1533 heart_block5_ck8 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1243 heart_block5_m_8_0_dff_s mbk_sig1535 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1244 vddi heart_block5_m_8_0_dff_s mbk_sig1535 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1245 heart_block5_s08 heart_block5_m_8_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1246 heart_block5_m_8_0_dff_m mbk_sig1526 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1247 mbk_sig1529 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1248 heart_block5_b22s heart_block5_s22 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1249 vddi heart_block5_b2 heart_block5_b22s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1250 heart_block5_a15s heart_block5_s15 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1251 vddi heart_block5_a5 heart_block5_a15s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1252 vddi mbk_sig1521 heart_block5_oa431s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1253 vddi heart_block5_a16s mbk_sig1521 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1254 mbk_sig1521 heart_block5_a17s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1255 vddi heart_block5_a18s mbk_sig1521 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1256 mbk_sig1521 heart_block5_a15s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1257 heart_block5_b01s heart_block5_s01 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1258 vddi heart_block5_b1 heart_block5_b01s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1259 vddi mbk_sig1514 heart_block5_ck4 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1260 vddi heart_block5_enable mbk_sig1514 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1261 mbk_sig1514 heart_block5_b4 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1262 heart_block5_a24s heart_block5_s24 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1263 vddi heart_block5_a4 heart_block5_a24s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1264 heart_block5_b28s heart_block5_s28 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1265 vddi heart_block5_b8 heart_block5_b28s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1266 vddi mbk_sig1506 heart_block5_ob441s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1267 vddi heart_block5_b12s mbk_sig1506 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1268 mbk_sig1506 heart_block5_b13s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1269 vddi heart_block5_b14s mbk_sig1506 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1270 mbk_sig1506 heart_block5_b11s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1271 heart_block5_a14s heart_block5_s14 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1272 vddi heart_block5_a4 heart_block5_a14s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1273 heart_block5_b14s heart_block5_s14 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1274 vddi heart_block5_b4 heart_block5_b14s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1275 heart_block5_a31s heart_block5_s31 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1276 vddi heart_block5_a1 heart_block5_a31s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1277 mbk_sig1496 mbk_sig1498 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1278 vddi heart_block5_m_4_1_dff_m mbk_sig1498 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1279 mbk_sig1497 heart_block5_ck4 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1280 heart_block5_m_4_1_dff_s mbk_sig1501 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1281 vddi heart_block5_m_4_1_dff_s mbk_sig1501 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1282 heart_block5_s14 heart_block5_m_4_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1283 heart_block5_m_4_1_dff_m mbk_sig1498 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1284 mbk_sig1493 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1285 vddi mbk_sig1491 heart_block5_oa443s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1286 vddi heart_block5_a32s mbk_sig1491 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1287 mbk_sig1491 heart_block5_a33s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1288 vddi heart_block5_a34s mbk_sig1491 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1289 mbk_sig1491 heart_block5_a31s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1290 mbk_sig1486 mbk_sig1481 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1291 vddi heart_block5_m_4_3_dff_m mbk_sig1481 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1292 mbk_sig1488 heart_block5_ck4 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1293 heart_block5_m_4_3_dff_s mbk_sig1487 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1294 vddi heart_block5_m_4_3_dff_s mbk_sig1487 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1295 heart_block5_s34 heart_block5_m_4_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1296 heart_block5_m_4_3_dff_m mbk_sig1481 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1297 mbk_sig1483 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1298 heart_block5_b34s heart_block5_s34 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1299 vddi heart_block5_b4 heart_block5_b34s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1300 heart_block5_b32s heart_block5_s32 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1301 vddi heart_block5_b2 heart_block5_b32s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1302 heart_block5_a32s heart_block5_s32 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1303 vddi heart_block5_a2 heart_block5_a32s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1304 heart_block5_b12s heart_block5_s12 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1305 vddi heart_block5_b2 heart_block5_b12s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1306 heart_block5_a03s heart_block5_s03 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1307 vddi heart_block5_a3 heart_block5_a03s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1308 heart_block3_cout2 heart_block3_na22 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1309 vddi heart_block3_gb2 heart_block3_cout2 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1310 heart_block3_na22 heart_block3_cout1 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1311 vddi heart_block3_not2 heart_block3_na22 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1312 mbk_sig1442 heart_block3_cout2 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1313 heart_block3_no43 heart_block3_n4 mbk_sig1442 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1314 mbk_sig1440 heart_block3_pb3 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1315 heart_block3_no33 heart_block3_n3 mbk_sig1440 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1316 vddi ii_5 heart_block3_ni5 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1317 mbk_sig1434 ii_5 vddi vddi TP L=0.18U W=1.98U AS=0.7128P AD=0.7128P 
+ PS=4.68U PD=4.68U 
M1318 vddi ii_3 mbk_sig1434 vddi TP L=0.18U W=1.98U AS=0.7128P AD=0.7128P 
+ PS=4.68U PD=4.68U 
M1319 mbk_sig1437 ii_5 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1320 heart_block3_nn0 ii_3 mbk_sig1437 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1321 vddi mbk_sig1434 heart_block3_nn0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1322 mbk_sig1430 heart_block3_no20 mbk_sig1429 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1323 vddi heart_block3_no30 mbk_sig1430 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1324 vddi heart_block3_no30 mbk_sig1433 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1325 mbk_sig1433 heart_block3_no20 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1326 heart_block3_x20 mbk_sig1429 mbk_sig1433 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1327 vddi heart_block3_g ngc vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1328 mbk_sig1428 heart_block3_x11 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1329 heart_block3_pb1 heart_block3_x01 mbk_sig1428 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1330 heart_block3_gb1 heart_block3_x11 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1331 vddi heart_block3_x01 heart_block3_gb1 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1332 mbk_sig1426 heart_block4_decaln vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1333 vddi heart_block4_ni7 mbk_sig1426 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1334 mbk_sig1426 heart_block4_ni6 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1335 vddi mbk_sig1426 heart_block4_selalu vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1336 mbk_sig1412 mbk_sig1413 mbk_sig1414 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1337 mbk_sig1414 heart_block4_shacc3 mbk_sig1412 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1338 mbk_sig1413 heart_block4_test_mode vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1339 mbk_sig1412 heart_q_2 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1340 vddi heart_block4_test_mode mbk_sig1412 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1341 heart_q_3 heart_block4_m3_dff_s vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1342 vddi heart_block4_m3_dff_s mbk_sig1421 vddi TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M1343 heart_block4_m3_dff_s mbk_sig1421 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1344 mbk_sig1420 mbk_sig1418 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1345 vddi heart_block4_m3_dff_m mbk_sig1418 vddi TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M1346 heart_block4_m3_dff_m mbk_sig1418 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1347 mbk_sig1417 heart_block4_ckin vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1348 vddi mbk_sig1409 heart_block5_a214sh vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1349 vddi heart_block2_a26ms_i0 mbk_sig1409 vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1350 mbk_sig1409 heart_block5_decaldra vddi vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1351 vddi mbk_sig1407 heart_block5_a29sh vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1352 vddi heart_block2_a25ms_i0 mbk_sig1407 vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1353 mbk_sig1407 heart_block5_decalgra vddi vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1354 mbk_sig1392 mbk_sig1397 mbk_sig1398 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1355 mbk_sig1398 heart_block4_shacc0 mbk_sig1392 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1356 mbk_sig1397 heart_block4_test_mode vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1357 mbk_sig1392 scini vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1358 vddi heart_block4_test_mode mbk_sig1392 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1359 heart_q_0 heart_block4_m0_dff_s vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1360 vddi heart_block4_m0_dff_s mbk_sig1406 vddi TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M1361 heart_block4_m0_dff_s mbk_sig1406 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1362 mbk_sig1404 mbk_sig1403 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1363 vddi heart_block4_m0_dff_m mbk_sig1403 vddi TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M1364 heart_block4_m0_dff_m mbk_sig1403 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1365 mbk_sig1402 heart_block4_ckin vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1366 mbk_sig1394 heart_block4_a217s mbk_sig1393 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1367 mbk_sig1389 heart_block4_a218s mbk_sig1394 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1368 vddi mbk_sig1389 heart_block4_shacc3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1369 mbk_sig1393 heart_block4_a216s vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M1370 vddi noei oec vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
M1371 vddi mbk_sig1387 heart_block4_a218s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1372 vddi heart_block4_insh2 mbk_sig1387 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1373 mbk_sig1387 heart_block4_decalga vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1374 vddi mbk_sig1385 heart_block4_a214s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1375 vddi heart_q_0 mbk_sig1385 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1376 mbk_sig1385 ii_8 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1377 vddi mbk_sig1384 scoutc vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1378 vddi heart_block4_test_mode mbk_sig1384 vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1379 mbk_sig1384 heart_q_3 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1380 mbk_sig1381 heart_block4_a210s vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M1381 mbk_sig1378 heart_block4_a214s mbk_sig1381 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1382 vddi mbk_sig1378 heart_block4_insh0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1383 heart_block5_b16s heart_block5_s16 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1384 vddi heart_block5_b6 heart_block5_b16s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1385 vddi ii_8 heart_block5_decalnr vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1386 heart_block5_a23s heart_block5_s23 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1387 vddi heart_block5_a3 heart_block5_a23s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1388 heart_block5_a36s heart_block5_s36 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1389 vddi heart_block5_a6 heart_block5_a36s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1390 vddi mbk_sig1371 heart_block5_oa442s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1391 vddi heart_block5_a22s mbk_sig1371 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1392 mbk_sig1371 heart_block5_a23s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1393 vddi heart_block5_a24s mbk_sig1371 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1394 mbk_sig1371 heart_block5_a21s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1395 heart_block5_b06s heart_block5_s06 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1396 vddi heart_block5_b6 heart_block5_b06s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1397 vddi mbk_sig1360 heart_block5_b9 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1398 vddi heart_block5_nb1 mbk_sig1360 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1399 mbk_sig1360 heart_block5_nb2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1400 vddi heart_b_3 mbk_sig1360 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1401 mbk_sig1360 heart_block5_nb0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1402 heart_block5_b07s heart_block5_s07 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1403 vddi heart_block5_b7 heart_block5_b07s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1404 vddi mbk_sig1356 heart_block5_oa430s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1405 vddi heart_block5_a06s mbk_sig1356 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1406 mbk_sig1356 heart_block5_a07s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1407 vddi heart_block5_a08s mbk_sig1356 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1408 mbk_sig1356 heart_block5_a05s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1409 vddi mbk_sig1350 heart_block5_ob430s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1410 vddi heart_block5_b06s mbk_sig1350 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1411 mbk_sig1350 heart_block5_b07s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1412 vddi heart_block5_b08s mbk_sig1350 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1413 mbk_sig1350 heart_block5_b05s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1414 heart_block5_b05s heart_block5_s05 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1415 vddi heart_block5_b5 heart_block5_b05s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1416 mbk_sig1347 mbk_sig1343 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1417 vddi heart_block5_m_7_0_dff_m mbk_sig1343 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1418 mbk_sig1345 heart_block5_ck7 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1419 heart_block5_m_7_0_dff_s mbk_sig1348 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1420 vddi heart_block5_m_7_0_dff_s mbk_sig1348 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1421 heart_block5_s07 heart_block5_m_7_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1422 heart_block5_m_7_0_dff_m mbk_sig1343 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1423 mbk_sig1342 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1424 heart_block5_a22s heart_block5_s22 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1425 vddi heart_block5_a2 heart_block5_a22s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1426 heart_block5_a07s heart_block5_s07 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1427 vddi heart_block5_a7 heart_block5_a07s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1428 heart_block5_a11s heart_block5_s11 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1429 vddi heart_block5_a1 heart_block5_a11s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1430 heart_block5_a05s heart_block5_s05 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1431 vddi heart_block5_a5 heart_block5_a05s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1432 vddi mbk_sig1333 heart_block5_oa441s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1433 vddi heart_block5_a12s mbk_sig1333 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1434 mbk_sig1333 heart_block5_a13s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1435 vddi heart_block5_a14s mbk_sig1333 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1436 mbk_sig1333 heart_block5_a11s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1437 heart_block5_a13s heart_block5_s13 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1438 vddi heart_block5_a3 heart_block5_a13s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1439 mbk_sig1326 mbk_sig1325 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1440 vddi heart_block5_m_3_1_dff_m mbk_sig1325 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1441 mbk_sig1328 heart_block5_ck3 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1442 heart_block5_m_3_1_dff_s mbk_sig1330 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1443 vddi heart_block5_m_3_1_dff_s mbk_sig1330 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1444 heart_block5_s13 heart_block5_m_3_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1445 heart_block5_m_3_1_dff_m mbk_sig1325 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1446 mbk_sig1322 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1447 heart_block5_b13s heart_block5_s13 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1448 vddi heart_block5_b3 heart_block5_b13s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1449 heart_block5_a01s heart_block5_s01 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1450 vddi heart_block5_a1 heart_block5_a01s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1451 vddi mbk_sig1317 heart_block5_oa433s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1452 vddi heart_block5_a36s mbk_sig1317 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1453 mbk_sig1317 heart_block5_a37s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1454 vddi heart_block5_a38s mbk_sig1317 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1455 mbk_sig1317 heart_block5_a35s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1456 vddi mbk_sig1312 heart_block5_ob440s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1457 vddi heart_block5_b02s mbk_sig1312 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1458 mbk_sig1312 heart_block5_b03s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1459 vddi heart_block5_b04s mbk_sig1312 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1460 mbk_sig1312 heart_block5_b01s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1461 heart_block5_b02s heart_block5_s02 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1462 vddi heart_block5_b2 heart_block5_b02s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1463 heart_block5_a35s heart_block5_s35 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1464 vddi heart_block5_a5 heart_block5_a35s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1465 heart_block5_b03s heart_block5_s03 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1466 vddi heart_block5_b3 heart_block5_b03s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1467 mbk_sig1300 mbk_sig1296 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1468 vddi heart_block5_m_2_2_dff_m mbk_sig1296 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1469 mbk_sig1302 heart_block5_ck2 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1470 heart_block5_m_2_2_dff_s mbk_sig1301 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1471 vddi heart_block5_m_2_2_dff_s mbk_sig1301 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1472 heart_block5_s22 heart_block5_m_2_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1473 heart_block5_m_2_2_dff_m mbk_sig1296 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1474 mbk_sig1298 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1475 heart_block5_a34s heart_block5_s34 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1476 vddi heart_block5_a4 heart_block5_a34s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1477 vddi mbk_sig1288 heart_block5_oa440s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1478 vddi heart_block5_a02s mbk_sig1288 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1479 mbk_sig1288 heart_block5_a03s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1480 vddi heart_block5_a04s mbk_sig1288 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1481 mbk_sig1288 heart_block5_a01s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1482 mbk_sig1283 mbk_sig1280 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1483 vddi heart_block5_m_3_0_dff_m mbk_sig1280 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1484 mbk_sig1285 heart_block5_ck3 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1485 heart_block5_m_3_0_dff_s mbk_sig1284 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1486 vddi heart_block5_m_3_0_dff_s mbk_sig1284 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1487 heart_block5_s03 heart_block5_m_3_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1488 heart_block5_m_3_0_dff_m mbk_sig1280 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1489 mbk_sig1279 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1490 vddi heart_block3_pb2 heart_block3_not2 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1491 vddi heart_block5_decalgra mbk_sig1220 vddi TP L=0.18U W=2.7U AS=0.972P 
+ AD=0.972P PS=6.12U PD=6.12U 
M1492 vddi mbk_sig1220 decalgrc vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1493 decalgrc mbk_sig1220 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1494 vddi heart_block3_pb0 heart_block3_not0 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1495 mbk_sig1243 heart_block3_pb3 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1496 mbk_sig1242 heart_block3_pb2 mbk_sig1243 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1497 heart_block3_no31_csh heart_block3_gb1 mbk_sig1242 vddi TP L=0.18U 
+ W=4.14U AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1498 mbk_sig1241 heart_block3_ngb3 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1499 mbk_sig1240 heart_block3_no31_csh mbk_sig1241 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1500 heart_block3_no32_csh heart_block3_no2_csh mbk_sig1240 vddi TP L=0.18U 
+ W=4.14U AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1501 vddi heart_block3_gb3 heart_block3_ngb3 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1502 mbk_sig1216 ii_5 vddi vddi TP L=0.18U W=1.98U AS=0.7128P AD=0.7128P 
+ PS=4.68U PD=4.68U 
M1503 vddi ii_4 mbk_sig1216 vddi TP L=0.18U W=1.98U AS=0.7128P AD=0.7128P 
+ PS=4.68U PD=4.68U 
M1504 mbk_sig1239 ii_5 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1505 heart_block3_nn1 ii_4 mbk_sig1239 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1506 vddi mbk_sig1216 heart_block3_nn1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1507 mbk_sig1237 heart_block3_gb2 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1508 heart_block3_no22 heart_block3_n2 mbk_sig1237 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1509 mbk_sig1238 heart_block3_pb2 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1510 heart_block3_no32 heart_block3_n3 mbk_sig1238 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1511 mbk_sig1236 heart_block3_gb0 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1512 heart_block3_no20 heart_block3_n2 mbk_sig1236 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1513 vddi heart_block3_nn0 heart_block3_n0 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1514 mbk_sig1235 heart_block3_pb1 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1515 mbk_sig1234 heart_block3_pb2 mbk_sig1235 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1516 heart_block3_no30_csh heart_block3_pb3 mbk_sig1234 vddi TP L=0.18U 
+ W=4.14U AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1517 mbk_sig1232 heart_block3_no22 mbk_sig1209 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1518 vddi heart_block3_no32 mbk_sig1232 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1519 vddi heart_block3_no32 mbk_sig1233 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1520 mbk_sig1233 heart_block3_no22 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1521 heart_block3_x22 mbk_sig1209 mbk_sig1233 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1522 vddi mbk_sig1208 heart_block5_a213sh vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1523 vddi heart_block2_a25ms_i0 mbk_sig1208 vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1524 mbk_sig1208 heart_block5_decalnr vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1525 mbk_sig1231 heart_block5_a213sh mbk_sig1230 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1526 mbk_sig1205 heart_block5_a214sh mbk_sig1231 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1527 vddi mbk_sig1205 heart_block5_shram0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1528 mbk_sig1230 heart_block5_a212sh vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M1529 vddi mbk_sig1204 heart_block5_a211sh vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1530 vddi heart_block2_a27ms_i0 mbk_sig1204 vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1531 mbk_sig1204 heart_block5_decaldra vddi vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1532 mbk_sig1229 heart_block5_a210sh mbk_sig1228 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1533 mbk_sig1202 heart_block5_a211sh mbk_sig1229 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1534 vddi mbk_sig1202 heart_block5_shram1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1535 mbk_sig1228 heart_block5_a29sh vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M1536 vddi mbk_sig1199 heart_block5_a210sh vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1537 vddi heart_block2_a26ms_i0 mbk_sig1199 vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1538 mbk_sig1199 heart_block5_decalnr vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1539 vddi mbk_sig1197 heart_block5_a212sh vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1540 vddi r0i mbk_sig1197 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1541 mbk_sig1197 heart_block5_decalgra vddi vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1542 vddi mbk_sig1194 heart_block5_a24sh vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1543 vddi heart_block2_a28ms_i0 mbk_sig1194 vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1544 mbk_sig1194 heart_block5_decalnr vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1545 mbk_sig1227 ii_8 vddi vddi TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
M1546 mbk_sig1192 heart_block4_ni7 mbk_sig1227 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1547 vddi mbk_sig1192 heart_block4_o21s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1548 vddi mbk_sig1191 heart_block5_decalgra vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1549 vddi ii_8 mbk_sig1191 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1550 mbk_sig1191 ii_7 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1551 mbk_sig1225 heart_block5_a24sh mbk_sig1226 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1552 mbk_sig1190 heart_block5_a25sh mbk_sig1225 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1553 vddi mbk_sig1190 heart_block5_shram3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1554 mbk_sig1226 heart_block5_a23sh vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M1555 vddi ii_7 heart_block4_ni7 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1556 vddi mbk_sig1186 heart_block5_a23sh vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1557 vddi heart_block2_a27ms_i0 mbk_sig1186 vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1558 mbk_sig1186 heart_block5_decalgra vddi vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1559 heart_block5_b313s heart_block5_s313 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1560 vddi heart_block5_b13 heart_block5_b313s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1561 heart_block5_b36s heart_block5_s36 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1562 vddi heart_block5_b6 heart_block5_b36s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1563 vddi mbk_sig1181 heart_block5_a25sh vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1564 vddi r3i mbk_sig1181 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1565 mbk_sig1181 heart_block5_decaldra vddi vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1566 mbk_sig1176 mbk_sig1178 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1567 vddi heart_block5_m_7_2_dff_m mbk_sig1178 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1568 mbk_sig1177 heart_block5_ck7 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1569 heart_block5_m_7_2_dff_s mbk_sig1180 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1570 vddi heart_block5_m_7_2_dff_s mbk_sig1180 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1571 heart_block5_s27 heart_block5_m_7_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1572 heart_block5_m_7_2_dff_m mbk_sig1178 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1573 mbk_sig1174 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1574 vddi mbk_sig1172 heart_block5_ck6 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1575 vddi heart_block5_enable mbk_sig1172 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1576 mbk_sig1172 heart_block5_b6 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1577 heart_block5_a06s heart_block5_s06 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1578 vddi heart_block5_a6 heart_block5_a06s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1579 mbk_sig1166 mbk_sig1162 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1580 vddi heart_block5_m_6_1_dff_m mbk_sig1162 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1581 mbk_sig1168 heart_block5_ck6 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1582 heart_block5_m_6_1_dff_s mbk_sig1167 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1583 vddi heart_block5_m_6_1_dff_s mbk_sig1167 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1584 heart_block5_s16 heart_block5_m_6_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1585 heart_block5_m_6_1_dff_m mbk_sig1162 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1586 mbk_sig1164 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1587 vddi mbk_sig1159 heart_block5_oa432s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1588 vddi heart_block5_a26s mbk_sig1159 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1589 mbk_sig1159 heart_block5_a27s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1590 vddi heart_block5_a28s mbk_sig1159 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1591 mbk_sig1159 heart_block5_a25s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1592 heart_block5_a26s heart_block5_s26 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1593 vddi heart_block5_a6 heart_block5_a26s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1594 heart_block5_a27s heart_block5_s27 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1595 vddi heart_block5_a7 heart_block5_a27s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1596 heart_block5_a08s heart_block5_s08 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1597 vddi heart_block5_a8 heart_block5_a08s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1598 heart_block5_a16s heart_block5_s16 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1599 vddi heart_block5_a6 heart_block5_a16s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1600 heart_block5_b08s heart_block5_s08 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1601 vddi heart_block5_b8 heart_block5_b08s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1602 mbk_sig1142 mbk_sig1138 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1603 vddi heart_block5_m_5_0_dff_m mbk_sig1138 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1604 mbk_sig1140 heart_block5_ck5 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1605 heart_block5_m_5_0_dff_s mbk_sig1144 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1606 vddi heart_block5_m_5_0_dff_s mbk_sig1144 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1607 heart_block5_s05 heart_block5_m_5_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1608 heart_block5_m_5_0_dff_m mbk_sig1138 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1609 mbk_sig1137 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1610 heart_block5_b35s heart_block5_s35 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1611 vddi heart_block5_b5 heart_block5_b35s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1612 heart_block5_a25s heart_block5_s25 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1613 vddi heart_block5_a5 heart_block5_a25s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1614 mbk_sig1130 mbk_sig1127 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1615 vddi heart_block5_m_11_3_dff_m mbk_sig1127 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1616 mbk_sig1131 heart_block5_ck11 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1617 heart_block5_m_11_3_dff_s mbk_sig1133 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1618 vddi heart_block5_m_11_3_dff_s mbk_sig1133 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1619 heart_block5_s311 heart_block5_m_11_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1620 heart_block5_m_11_3_dff_m mbk_sig1127 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1621 mbk_sig1125 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1622 mbk_sig1122 mbk_sig1118 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1623 vddi heart_block5_m_5_3_dff_m mbk_sig1118 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1624 mbk_sig1124 heart_block5_ck5 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1625 heart_block5_m_5_3_dff_s mbk_sig1123 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1626 vddi heart_block5_m_5_3_dff_s mbk_sig1123 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1627 heart_block5_s35 heart_block5_m_5_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1628 heart_block5_m_5_3_dff_m mbk_sig1118 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1629 mbk_sig1117 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1630 mbk_sig1115 mbk_sig1111 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1631 vddi heart_block5_m_2_0_dff_m mbk_sig1111 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1632 mbk_sig1113 heart_block5_ck2 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1633 heart_block5_m_2_0_dff_s mbk_sig1116 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1634 vddi heart_block5_m_2_0_dff_s mbk_sig1116 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1635 heart_block5_s02 heart_block5_m_2_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1636 heart_block5_m_2_0_dff_m mbk_sig1111 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1637 mbk_sig1110 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1638 mbk_sig1105 mbk_sig1107 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1639 vddi heart_block5_m_2_1_dff_m mbk_sig1107 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1640 mbk_sig1106 heart_block5_ck2 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1641 heart_block5_m_2_1_dff_s mbk_sig1109 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1642 vddi heart_block5_m_2_1_dff_s mbk_sig1109 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1643 heart_block5_s12 heart_block5_m_2_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1644 heart_block5_m_2_1_dff_m mbk_sig1107 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1645 mbk_sig1101 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1646 heart_block5_a12s heart_block5_s12 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1647 vddi heart_block5_a2 heart_block5_a12s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1648 heart_block5_b310s heart_block5_s310 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1649 vddi heart_block5_b10 heart_block5_b310s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1650 vddi mbk_sig1097 heart_block5_ck10 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1651 vddi heart_block5_enable mbk_sig1097 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1652 mbk_sig1097 heart_block5_b10 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1653 mbk_sig1094 mbk_sig1090 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1654 vddi heart_block5_m_10_3_dff_m mbk_sig1090 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1655 mbk_sig1095 heart_block5_ck10 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1656 heart_block5_m_10_3_dff_s mbk_sig1096 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1657 vddi heart_block5_m_10_3_dff_s mbk_sig1096 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1658 heart_block5_s310 heart_block5_m_10_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1659 heart_block5_m_10_3_dff_m mbk_sig1090 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1660 mbk_sig1092 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1661 heart_block5_a02s heart_block5_s02 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1662 vddi heart_block5_a2 heart_block5_a02s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1663 heart_block5_a010s heart_block5_s010 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1664 vddi heart_block5_a10 heart_block5_a010s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1665 heart_block3_gb0 heart_block3_x10 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1666 vddi heart_block3_x00 heart_block3_gb0 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1667 heart_block3_na23 heart_block3_cout2 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1668 vddi heart_block3_not3 heart_block3_na23 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1669 heart_block3_couta heart_block3_na23 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1670 vddi heart_block3_gb3 heart_block3_couta vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1671 mbk_sig1065 heart_block3_pb0 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1672 heart_block3_no30 heart_block3_n3 mbk_sig1065 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1673 mbk_sig1063 heart_block1_sra1 mbk_sig1064 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1674 mbk_sig1050 heart_block1_srq1 mbk_sig1063 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1675 vddi mbk_sig1050 heart_s_1 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1676 mbk_sig1064 heart_block1_srb1 vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M1677 mbk_sig1061 heart_s_1 mbk_sig1049 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1678 vddi heart_block3_n1 mbk_sig1061 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1679 vddi heart_block3_n1 mbk_sig1062 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1680 mbk_sig1062 heart_s_1 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1681 heart_block3_x11 mbk_sig1049 mbk_sig1062 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1682 mbk_sig1059 heart_block3_cout2 mbk_sig1046 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1683 vddi heart_block3_couta mbk_sig1059 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1684 vddi heart_block3_couta mbk_sig1060 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1685 mbk_sig1060 heart_block3_cout2 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1686 ovrc mbk_sig1046 mbk_sig1060 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1687 vddi mbk_sig1042 heart_block1_srq1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1688 vddi heart_q_1 mbk_sig1042 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1689 mbk_sig1042 heart_block1_selqs vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1690 mbk_sig1058 heart_block3_pb3 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1691 heart_block3_no2_csh heart_block3_gb2 mbk_sig1058 vddi TP L=0.18U 
+ W=4.14U AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1692 vddi heart_block3_gb0 heart_block3_ngb0 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1693 vddi heart_block3_p npc vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1694 vddi mbk_sig1037 coutc vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1695 vddi heart_block3_couta mbk_sig1037 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1696 mbk_sig1037 heart_block3_flag vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1697 vddi heart_block3_nprop heart_block3_propf vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1698 vddi heart_block5_decaldra mbk_sig1035 vddi TP L=0.18U W=2.7U AS=0.972P 
+ AD=0.972P PS=6.12U PD=6.12U 
M1699 vddi mbk_sig1035 decaldrc vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1700 decaldrc mbk_sig1035 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1701 vddi mbk_sig1034 heart_block3_p vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1702 vddi heart_block3_propf mbk_sig1034 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1703 mbk_sig1034 heart_block3_flag vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1704 vddi ii_7 heart_block5_ni7 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1705 vddi mbk_sig1030 heart_block2_syalu3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1706 vddi heart_block2_a28ms_i0 mbk_sig1030 vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1707 mbk_sig1030 heart_block2_selaluy vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1708 vddi mbk_sig1028 heart_block5_decaldra vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1709 vddi ii_8 mbk_sig1028 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1710 mbk_sig1028 heart_block5_ni7 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1711 mbk_sig1057 heart_block2_syra3 vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M1712 mbk_sig1023 heart_block2_syalu3 mbk_sig1057 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1713 vddi mbk_sig1023 yc_3 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1714 vddi mbk_sig1022 s0c vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1715 vddi heart_block5_decaldra mbk_sig1022 vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1716 mbk_sig1022 heart_block2_a25ms_i0 vddi vddi TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M1717 vddi mbk_sig1020 heart_block1_srq0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1718 vddi heart_q_0 mbk_sig1020 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1719 mbk_sig1020 heart_block1_selqs vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1720 vddi mbk_sig1016 heart_block4_decalga vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1721 vddi ii_8 mbk_sig1016 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1722 mbk_sig1016 ii_7 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1723 vddi mbk_sig1013 heart_block1_srb3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1724 vddi heart_rb_3 mbk_sig1013 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1725 mbk_sig1013 heart_block1_selbs vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1726 vddi mbk_sig1012 heart_block5_ck16 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1727 vddi heart_block5_enable mbk_sig1012 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1728 mbk_sig1012 heart_block5_b16 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1729 vddi mbk_sig1011 heart_block5_ck13 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1730 vddi heart_block5_enable mbk_sig1011 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1731 mbk_sig1011 heart_block5_b13 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1732 heart_block5_b113s heart_block5_s113 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1733 vddi heart_block5_b13 heart_block5_b113s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1734 heart_block5_b116s heart_block5_s116 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1735 vddi heart_block5_b16 heart_block5_b116s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1736 mbk_sig1003 mbk_sig1002 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1737 vddi heart_block5_m_6_0_dff_m mbk_sig1002 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1738 mbk_sig1004 heart_block5_ck6 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1739 heart_block5_m_6_0_dff_s mbk_sig1008 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1740 vddi heart_block5_m_6_0_dff_s mbk_sig1008 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1741 heart_block5_s06 heart_block5_m_6_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1742 heart_block5_m_6_0_dff_m mbk_sig1002 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1743 mbk_sig1000 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1744 heart_block5_b316s heart_block5_s316 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1745 vddi heart_block5_b16 heart_block5_b316s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1746 vddi mbk_sig994 heart_block5_ob413s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1747 vddi heart_block5_b314s mbk_sig994 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1748 mbk_sig994 heart_block5_b315s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1749 vddi heart_block5_b316s mbk_sig994 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1750 mbk_sig994 heart_block5_b313s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1751 mbk_sig991 mbk_sig990 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1752 vddi heart_block5_m_16_3_dff_m mbk_sig990 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1753 mbk_sig989 heart_block5_ck16 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1754 heart_block5_m_16_3_dff_s mbk_sig993 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1755 vddi heart_block5_m_16_3_dff_s mbk_sig993 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1756 heart_block5_s316 heart_block5_m_16_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1757 heart_block5_m_16_3_dff_m mbk_sig990 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1758 mbk_sig987 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1759 heart_rb_2 heart_block5_ob442s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1760 vddi heart_block5_ob432s heart_rb_2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1761 heart_rb_2 heart_block5_ob422s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1762 vddi heart_block5_ob412s heart_rb_2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1763 heart_block5_b315s heart_block5_s315 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1764 vddi heart_block5_b15 heart_block5_b315s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1765 vddi mbk_sig974 heart_block5_ob433s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1766 vddi heart_block5_b36s mbk_sig974 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1767 mbk_sig974 heart_block5_b37s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1768 vddi heart_block5_b38s mbk_sig974 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1769 mbk_sig974 heart_block5_b35s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1770 mbk_sig969 mbk_sig971 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1771 vddi heart_block5_m_7_3_dff_m mbk_sig971 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1772 mbk_sig970 heart_block5_ck7 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1773 heart_block5_m_7_3_dff_s mbk_sig973 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1774 vddi heart_block5_m_7_3_dff_s mbk_sig973 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1775 heart_block5_s37 heart_block5_m_7_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1776 heart_block5_m_7_3_dff_m mbk_sig971 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1777 mbk_sig967 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1778 heart_rb_3 heart_block5_ob443s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1779 vddi heart_block5_ob433s heart_rb_3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1780 heart_rb_3 heart_block5_ob423s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1781 vddi heart_block5_ob413s heart_rb_3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1782 mbk_sig958 mbk_sig955 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1783 vddi heart_block5_m_11_2_dff_m mbk_sig955 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1784 mbk_sig960 heart_block5_ck11 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1785 heart_block5_m_11_2_dff_s mbk_sig961 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1786 vddi heart_block5_m_11_2_dff_s mbk_sig961 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1787 heart_block5_s211 heart_block5_m_11_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1788 heart_block5_m_11_2_dff_m mbk_sig955 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1789 mbk_sig957 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1790 heart_block5_b211s heart_block5_s211 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1791 vddi heart_block5_b11 heart_block5_b211s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1792 vddi mbk_sig952 heart_block5_a3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1793 vddi heart_a_1 mbk_sig952 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1794 mbk_sig952 heart_block5_na2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1795 vddi heart_block5_na3 mbk_sig952 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1796 mbk_sig952 heart_block5_na0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1797 vddi mbk_sig948 heart_block5_a5 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1798 vddi heart_block5_na1 mbk_sig948 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1799 mbk_sig948 heart_a_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1800 vddi heart_block5_na3 mbk_sig948 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1801 mbk_sig948 heart_block5_na0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1802 heart_block5_a37s heart_block5_s37 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1803 vddi heart_block5_a7 heart_block5_a37s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1804 heart_block5_b29s heart_block5_s29 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1805 vddi heart_block5_b9 heart_block5_b29s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1806 vddi mbk_sig937 heart_block5_ob422s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1807 vddi heart_block5_b210s mbk_sig937 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1808 mbk_sig937 heart_block5_b211s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1809 vddi heart_block5_b212s mbk_sig937 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1810 mbk_sig937 heart_block5_b29s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1811 vddi mbk_sig933 heart_block5_a7 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1812 vddi heart_a_1 mbk_sig933 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1813 mbk_sig933 heart_a_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1814 vddi heart_block5_na3 mbk_sig933 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1815 mbk_sig933 heart_block5_na0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1816 heart_block5_b210s heart_block5_s210 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1817 vddi heart_block5_b10 heart_block5_b210s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1818 heart_block5_b311s heart_block5_s311 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1819 vddi heart_block5_b11 heart_block5_b311s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1820 vddi mbk_sig927 heart_block5_a4 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1821 vddi heart_a_1 mbk_sig927 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1822 mbk_sig927 heart_block5_na2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1823 vddi heart_block5_na3 mbk_sig927 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1824 mbk_sig927 heart_a_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1825 heart_block5_a311s heart_block5_s311 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1826 vddi heart_block5_a11 heart_block5_a311s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1827 vddi mbk_sig918 heart_block5_ob423s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1828 vddi heart_block5_b310s mbk_sig918 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1829 mbk_sig918 heart_block5_b311s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1830 vddi heart_block5_b312s mbk_sig918 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1831 mbk_sig918 heart_block5_b39s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1832 mbk_sig913 mbk_sig915 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1833 vddi heart_block5_m_10_0_dff_m mbk_sig915 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1834 mbk_sig914 heart_block5_ck10 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1835 heart_block5_m_10_0_dff_s mbk_sig917 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1836 vddi heart_block5_m_10_0_dff_s mbk_sig917 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1837 heart_block5_s010 heart_block5_m_10_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1838 heart_block5_m_10_0_dff_m mbk_sig915 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1839 mbk_sig911 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1840 mbk_sig907 mbk_sig906 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1841 vddi heart_block5_m_10_1_dff_m mbk_sig906 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1842 mbk_sig908 heart_block5_ck10 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1843 heart_block5_m_10_1_dff_s mbk_sig910 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1844 vddi heart_block5_m_10_1_dff_s mbk_sig910 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1845 heart_block5_s110 heart_block5_m_10_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1846 heart_block5_m_10_1_dff_m mbk_sig906 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1847 mbk_sig905 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1848 mbk_sig867 heart_r_0 mbk_sig866 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1849 vddi heart_block3_n0 mbk_sig867 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1850 vddi heart_block3_n0 mbk_sig868 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1851 mbk_sig868 heart_r_0 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1852 heart_block3_x00 mbk_sig866 mbk_sig868 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1853 mbk_sig864 heart_block3_x10 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1854 heart_block3_pb0 heart_block3_x00 mbk_sig864 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1855 vddi heart_block3_pb3 heart_block3_not3 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1856 vddi mbk_sig861 heart_block3_ngen vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1857 vddi heart_block3_na_csh mbk_sig861 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1858 mbk_sig861 heart_block3_no32_csh vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1859 heart_block3_na_csh heart_block3_no30_csh vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1860 vddi heart_block3_ngb0 heart_block3_na_csh vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1861 mbk_sig857 heart_block3_x12 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1862 heart_block3_pb2 heart_block3_x02 mbk_sig857 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1863 mbk_sig854 heart_r_3 mbk_sig853 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1864 vddi heart_block3_n0 mbk_sig854 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1865 vddi heart_block3_n0 mbk_sig855 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1866 mbk_sig855 heart_r_3 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1867 heart_block3_x03 mbk_sig853 mbk_sig855 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1868 mbk_sig851 heart_block3_x13 vddi vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1869 heart_block3_pb3 heart_block3_x03 mbk_sig851 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1870 heart_block3_gb3 heart_block3_x13 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1871 vddi heart_block3_x03 heart_block3_gb3 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1872 vddi heart_block3_ngen heart_block3_genf vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1873 vddi mbk_sig844 heart_block3_g vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1874 vddi heart_block3_genf mbk_sig844 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1875 mbk_sig844 heart_block3_flag vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1876 heart_block3_nprop heart_block3_no30_csh vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1877 vddi heart_block3_npb0 heart_block3_nprop vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1878 mbk_sig838 heart_s_3 mbk_sig837 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1879 vddi heart_block3_n1 mbk_sig838 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1880 vddi heart_block3_n1 mbk_sig839 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M1881 mbk_sig839 heart_s_3 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M1882 heart_block3_x13 mbk_sig837 mbk_sig839 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1883 mbk_sig835 heart_block1_sra3 mbk_sig836 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1884 mbk_sig832 heart_block1_srq3 mbk_sig835 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M1885 vddi mbk_sig832 heart_s_3 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1886 mbk_sig836 heart_block1_srb3 vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M1887 vddi mbk_sig830 heart_block1_srq3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1888 vddi heart_q_3 mbk_sig830 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1889 mbk_sig830 heart_block1_selqs vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1890 mbk_sig828 mbk_sig824 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1891 vddi heart_block5_m_13_0_dff_m mbk_sig824 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1892 mbk_sig826 heart_block5_ck13 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1893 heart_block5_m_13_0_dff_s mbk_sig829 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1894 vddi heart_block5_m_13_0_dff_s mbk_sig829 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1895 heart_block5_s013 heart_block5_m_13_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1896 heart_block5_m_13_0_dff_m mbk_sig824 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1897 mbk_sig822 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1898 mbk_sig820 mbk_sig815 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1899 vddi heart_block5_m_13_2_dff_m mbk_sig815 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1900 mbk_sig821 heart_block5_ck13 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1901 heart_block5_m_13_2_dff_s mbk_sig823 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1902 vddi heart_block5_m_13_2_dff_s mbk_sig823 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1903 heart_block5_s213 heart_block5_m_13_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1904 heart_block5_m_13_2_dff_m mbk_sig815 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1905 mbk_sig818 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1906 heart_block5_a213s heart_block5_s213 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1907 vddi heart_block5_a13 heart_block5_a213s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1908 mbk_sig810 mbk_sig812 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1909 vddi heart_block5_m_16_1_dff_m mbk_sig812 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1910 mbk_sig811 heart_block5_ck16 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1911 heart_block5_m_16_1_dff_s mbk_sig814 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1912 vddi heart_block5_m_16_1_dff_s mbk_sig814 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1913 heart_block5_s116 heart_block5_m_16_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1914 heart_block5_m_16_1_dff_m mbk_sig812 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1915 mbk_sig808 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1916 heart_block5_b214s heart_block5_s214 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1917 vddi heart_block5_b14 heart_block5_b214s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1918 heart_block5_a113s heart_block5_s113 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1919 vddi heart_block5_a13 heart_block5_a113s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1920 heart_block5_b213s heart_block5_s213 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1921 vddi heart_block5_b13 heart_block5_b213s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1922 mbk_sig799 mbk_sig801 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1923 vddi heart_block5_m_6_2_dff_m mbk_sig801 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1924 mbk_sig800 heart_block5_ck6 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1925 heart_block5_m_6_2_dff_s mbk_sig804 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1926 vddi heart_block5_m_6_2_dff_s mbk_sig804 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1927 heart_block5_s26 heart_block5_m_6_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1928 heart_block5_m_6_2_dff_m mbk_sig801 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1929 mbk_sig796 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1930 heart_block5_b216s heart_block5_s216 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1931 vddi heart_block5_b16 heart_block5_b216s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1932 vddi mbk_sig793 heart_block5_ob412s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1933 vddi heart_block5_b214s mbk_sig793 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1934 mbk_sig793 heart_block5_b215s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1935 vddi heart_block5_b216s mbk_sig793 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1936 mbk_sig793 heart_block5_b213s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1937 heart_block5_a216s heart_block5_s216 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1938 vddi heart_block5_a16 heart_block5_a216s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1939 vddi mbk_sig787 heart_block5_oa412s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1940 vddi heart_block5_a214s mbk_sig787 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1941 mbk_sig787 heart_block5_a215s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1942 vddi heart_block5_a216s mbk_sig787 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1943 mbk_sig787 heart_block5_a213s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1944 heart_rb_0 heart_block5_ob440s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1945 vddi heart_block5_ob430s heart_rb_0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1946 heart_rb_0 heart_block5_ob420s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1947 vddi heart_block5_ob410s heart_rb_0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1948 heart_block5_b115s heart_block5_s115 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1949 vddi heart_block5_b15 heart_block5_b115s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1950 vddi mbk_sig779 heart_block5_ob411s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1951 vddi heart_block5_b114s mbk_sig779 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1952 mbk_sig779 heart_block5_b115s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1953 vddi heart_block5_b116s mbk_sig779 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1954 mbk_sig779 heart_block5_b113s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1955 heart_ra_0 heart_block5_oa440s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1956 vddi heart_block5_oa430s heart_ra_0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1957 heart_ra_0 heart_block5_oa420s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1958 vddi heart_block5_oa410s heart_ra_0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1959 heart_block5_b37s heart_block5_s37 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1960 vddi heart_block5_b7 heart_block5_b37s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M1961 vddi mbk_sig773 heart_block5_ck15 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1962 vddi heart_block5_enable mbk_sig773 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1963 mbk_sig773 heart_block5_b15 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1964 vddi mbk_sig768 heart_block5_a8 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1965 vddi heart_a_1 mbk_sig768 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1966 mbk_sig768 heart_a_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1967 vddi heart_block5_na3 mbk_sig768 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1968 mbk_sig768 heart_a_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M1969 mbk_sig762 mbk_sig764 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1970 vddi heart_block5_m_15_1_dff_m mbk_sig764 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1971 mbk_sig763 heart_block5_ck15 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1972 heart_block5_m_15_1_dff_s mbk_sig767 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1973 vddi heart_block5_m_15_1_dff_s mbk_sig767 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1974 heart_block5_s115 heart_block5_m_15_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1975 heart_block5_m_15_1_dff_m mbk_sig764 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1976 mbk_sig759 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1977 vddi mbk_sig758 heart_block5_ck11 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1978 vddi heart_block5_enable mbk_sig758 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1979 mbk_sig758 heart_block5_b11 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1980 mbk_sig753 mbk_sig755 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1981 vddi heart_block5_m_9_3_dff_m mbk_sig755 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1982 mbk_sig754 heart_block5_ck9 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1983 heart_block5_m_9_3_dff_s mbk_sig757 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1984 vddi heart_block5_m_9_3_dff_s mbk_sig757 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1985 heart_block5_s39 heart_block5_m_9_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1986 heart_block5_m_9_3_dff_m mbk_sig755 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1987 mbk_sig750 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1988 vddi mbk_sig749 heart_block5_a1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M1989 vddi heart_block5_na1 mbk_sig749 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1990 mbk_sig749 heart_block5_na2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1991 vddi heart_block5_na3 mbk_sig749 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1992 mbk_sig749 heart_block5_na0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M1993 mbk_sig743 mbk_sig738 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M1994 vddi heart_block5_m_10_2_dff_m mbk_sig738 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1995 mbk_sig745 heart_block5_ck10 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M1996 heart_block5_m_10_2_dff_s mbk_sig744 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M1997 vddi heart_block5_m_10_2_dff_s mbk_sig744 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M1998 heart_block5_s210 heart_block5_m_10_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M1999 heart_block5_m_10_2_dff_m mbk_sig738 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2000 mbk_sig740 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2001 vddi mbk_sig736 heart_block5_a13 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2002 vddi heart_block5_na1 mbk_sig736 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2003 mbk_sig736 heart_a_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2004 vddi heart_a_3 mbk_sig736 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2005 mbk_sig736 heart_block5_na0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2006 heart_block5_b39s heart_block5_s39 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2007 vddi heart_block5_b9 heart_block5_b39s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2008 vddi heart_a_1 heart_block5_na1 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2009 heart_block5_a210s heart_block5_s210 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2010 vddi heart_block5_a10 heart_block5_a210s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2011 vddi mbk_sig729 heart_block5_a2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2012 vddi heart_block5_na1 mbk_sig729 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2013 mbk_sig729 heart_block5_na2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2014 vddi heart_block5_na3 mbk_sig729 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2015 mbk_sig729 heart_a_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2016 heart_block5_b312s heart_block5_s312 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2017 vddi heart_block5_b12 heart_block5_b312s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2018 vddi mbk_sig721 heart_block5_a10 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2019 vddi heart_block5_na1 mbk_sig721 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2020 mbk_sig721 heart_block5_na2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2021 vddi heart_a_3 mbk_sig721 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2022 mbk_sig721 heart_a_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2023 heart_block5_b010s heart_block5_s010 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2024 vddi heart_block5_b10 heart_block5_b010s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2025 vddi heart_a_0 heart_block5_na0 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2026 mbk_sig678 heart_s_2 mbk_sig667 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2027 vddi heart_block3_n1 mbk_sig678 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2028 vddi heart_block3_n1 mbk_sig679 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2029 mbk_sig679 heart_s_2 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M2030 heart_block3_x12 mbk_sig667 mbk_sig679 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2031 vddi heart_block3_nn1 heart_block3_n1 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2032 mbk_sig676 heart_block1_sra0 mbk_sig677 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M2033 mbk_sig663 heart_block1_srq0 mbk_sig676 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M2034 vddi mbk_sig663 heart_s_0 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2035 mbk_sig677 heart_block1_srb0 vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M2036 mbk_sig675 heart_s_0 mbk_sig662 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2037 vddi heart_block3_n1 mbk_sig675 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2038 vddi heart_block3_n1 mbk_sig674 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2039 mbk_sig674 heart_s_0 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M2040 heart_block3_x10 mbk_sig662 mbk_sig674 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2041 vddi heart_block3_pb0 heart_block3_npb0 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2042 vddi mbk_sig656 heart_block1_sra0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2043 vddi heart_ra_0 mbk_sig656 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2044 mbk_sig656 heart_block1_selas vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2045 vddi mbk_sig654 heart_block4_ckin vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2046 vddi cko mbk_sig654 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2047 mbk_sig654 heart_block4_w vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2048 heart_block3_gb2 heart_block3_x12 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2049 vddi heart_block3_x02 heart_block3_gb2 vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2050 mbk_sig673 heart_block4_test_mode vddi vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M2051 mbk_sig648 heart_block4_a231s mbk_sig673 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M2052 vddi mbk_sig648 heart_block4_w vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2053 vddi mbk_sig646 heart_fonc_mode vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2054 vddi fonci mbk_sig646 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2055 mbk_sig646 heart_block4_n15s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2056 vddi ii_6 heart_block4_ni6 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2057 vddi mbk_sig642 heart_block4_a231s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2058 vddi heart_fonc_mode mbk_sig642 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2059 mbk_sig642 heart_block4_waccu vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2060 vddi mbk_sig641 heart_block4_waccu vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2061 vddi heart_block4_o21s mbk_sig641 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2062 mbk_sig641 heart_block4_ni6 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2063 vddi fonci heart_block4_n14s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2064 vddi mbk_sig639 heart_block2_syra3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2065 vddi heart_ra_3 mbk_sig639 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2066 mbk_sig639 heart_block2_selray vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2067 vddi mbk_sig634 heart_block2_syalu2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2068 vddi heart_block2_a27ms_i0 mbk_sig634 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2069 mbk_sig634 heart_block2_selaluy vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2070 heart_block5_a313s heart_block5_s313 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2071 vddi heart_block5_a13 heart_block5_a313s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2072 vddi mbk_sig630 heart_block2_syalu0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2073 vddi heart_block2_a25ms_i0 mbk_sig630 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2074 mbk_sig630 heart_block2_selaluy vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2075 vddi mbk_sig628 heart_block2_syra0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2076 vddi heart_ra_0 mbk_sig628 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2077 mbk_sig628 heart_block2_selray vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2078 mbk_sig672 heart_block2_syra0 vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M2079 mbk_sig624 heart_block2_syalu0 mbk_sig672 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M2080 vddi mbk_sig624 yc_0 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2081 vddi mbk_sig623 heart_block1_srb2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2082 vddi heart_rb_2 mbk_sig623 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2083 mbk_sig623 heart_block1_selbs vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2084 vddi mbk_sig621 heart_block1_srb0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2085 vddi heart_rb_0 mbk_sig621 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2086 mbk_sig621 heart_block1_selbs vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2087 mbk_sig617 mbk_sig612 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2088 vddi heart_block5_m_13_1_dff_m mbk_sig612 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2089 mbk_sig614 heart_block5_ck13 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2090 heart_block5_m_13_1_dff_s mbk_sig619 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2091 vddi heart_block5_m_13_1_dff_s mbk_sig619 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2092 heart_block5_s113 heart_block5_m_13_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2093 heart_block5_m_13_1_dff_m mbk_sig612 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2094 mbk_sig609 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2095 vddi mbk_sig610 heart_block1_srb1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2096 vddi heart_rb_1 mbk_sig610 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2097 mbk_sig610 heart_block1_selbs vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2098 heart_block5_a013s heart_block5_s013 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2099 vddi heart_block5_a13 heart_block5_a013s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2100 vddi mbk_sig605 heart_block5_ob410s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2101 vddi heart_block5_b014s mbk_sig605 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2102 mbk_sig605 heart_block5_b015s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2103 vddi heart_block5_b016s mbk_sig605 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2104 mbk_sig605 heart_block5_b013s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2105 mbk_sig597 mbk_sig593 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2106 vddi heart_block5_m_16_2_dff_m mbk_sig593 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2107 mbk_sig595 heart_block5_ck16 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2108 heart_block5_m_16_2_dff_s mbk_sig599 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2109 vddi heart_block5_m_16_2_dff_s mbk_sig599 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2110 heart_block5_s216 heart_block5_m_16_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2111 heart_block5_m_16_2_dff_m mbk_sig593 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2112 mbk_sig596 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2113 heart_block5_a214s heart_block5_s214 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2114 vddi heart_block5_a14 heart_block5_a214s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2115 vddi mbk_sig589 heart_block5_oa413s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2116 vddi heart_block5_a314s mbk_sig589 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2117 mbk_sig589 heart_block5_a315s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2118 vddi heart_block5_a316s mbk_sig589 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2119 mbk_sig589 heart_block5_a313s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2120 heart_block5_a316s heart_block5_s316 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2121 vddi heart_block5_a16 heart_block5_a316s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2122 heart_block5_b013s heart_block5_s013 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2123 vddi heart_block5_b13 heart_block5_b013s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2124 heart_block5_a315s heart_block5_s315 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2125 vddi heart_block5_a15 heart_block5_a315s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2126 heart_block5_a115s heart_block5_s115 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2127 vddi heart_block5_a15 heart_block5_a115s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2128 heart_block5_b215s heart_block5_s215 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2129 vddi heart_block5_b15 heart_block5_b215s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2130 heart_rb_1 heart_block5_ob441s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2131 vddi heart_block5_ob431s heart_rb_1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2132 heart_rb_1 heart_block5_ob421s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2133 vddi heart_block5_ob411s heart_rb_1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2134 vddi mbk_sig569 heart_block5_ck9 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2135 vddi heart_block5_enable mbk_sig569 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2136 mbk_sig569 heart_block5_b9 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2137 vddi mbk_sig566 heart_block5_a16 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2138 vddi heart_a_1 mbk_sig566 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2139 mbk_sig566 heart_a_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2140 vddi heart_a_3 mbk_sig566 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2141 mbk_sig566 heart_a_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2142 heart_ra_1 heart_block5_oa441s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2143 vddi heart_block5_oa431s heart_ra_1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2144 heart_ra_1 heart_block5_oa421s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2145 vddi heart_block5_oa411s heart_ra_1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2146 mbk_sig556 mbk_sig553 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2147 vddi heart_block5_m_15_2_dff_m mbk_sig553 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2148 mbk_sig558 heart_block5_ck15 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2149 heart_block5_m_15_2_dff_s mbk_sig559 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2150 vddi heart_block5_m_15_2_dff_s mbk_sig559 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2151 heart_block5_s215 heart_block5_m_15_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2152 heart_block5_m_15_2_dff_m mbk_sig553 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2153 mbk_sig555 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2154 mbk_sig549 mbk_sig546 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2155 vddi heart_block5_m_15_3_dff_m mbk_sig546 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2156 mbk_sig548 heart_block5_ck15 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2157 heart_block5_m_15_3_dff_s mbk_sig552 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2158 vddi heart_block5_m_15_3_dff_s mbk_sig552 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2159 heart_block5_s315 heart_block5_m_15_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2160 heart_block5_m_15_3_dff_m mbk_sig546 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2161 mbk_sig543 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2162 mbk_sig540 mbk_sig542 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2163 vddi heart_block5_m_9_2_dff_m mbk_sig542 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2164 mbk_sig541 heart_block5_ck9 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2165 heart_block5_m_9_2_dff_s mbk_sig545 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2166 vddi heart_block5_m_9_2_dff_s mbk_sig545 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2167 heart_block5_s29 heart_block5_m_9_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2168 heart_block5_m_9_2_dff_m mbk_sig542 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2169 mbk_sig539 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2170 vddi mbk_sig536 heart_block5_a6 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2171 vddi heart_block5_na1 mbk_sig536 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2172 mbk_sig536 heart_a_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2173 vddi heart_block5_na3 mbk_sig536 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2174 mbk_sig536 heart_a_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2175 vddi heart_a_3 heart_block5_na3 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2176 vddi mbk_sig528 heart_block5_a14 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2177 vddi heart_block5_na1 mbk_sig528 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2178 mbk_sig528 heart_a_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2179 vddi heart_a_3 mbk_sig528 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2180 mbk_sig528 heart_a_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2181 heart_ra_3 heart_block5_oa443s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2182 vddi heart_block5_oa433s heart_ra_3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2183 heart_ra_3 heart_block5_oa423s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2184 vddi heart_block5_oa413s heart_ra_3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2185 heart_block5_a312s heart_block5_s312 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2186 vddi heart_block5_a12 heart_block5_a312s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2187 vddi mbk_sig517 heart_block5_oa423s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2188 vddi heart_block5_a310s mbk_sig517 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2189 mbk_sig517 heart_block5_a311s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2190 vddi heart_block5_a312s mbk_sig517 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2191 mbk_sig517 heart_block5_a39s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2192 heart_block5_a39s heart_block5_s39 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2193 vddi heart_block5_a9 heart_block5_a39s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2194 vddi mbk_sig514 heart_block5_a11 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2195 vddi heart_a_1 mbk_sig514 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2196 mbk_sig514 heart_block5_na2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2197 vddi heart_a_3 mbk_sig514 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2198 mbk_sig514 heart_block5_na0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2199 heart_block5_b212s heart_block5_s212 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2200 vddi heart_block5_b12 heart_block5_b212s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2201 mbk_sig504 mbk_sig502 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2202 vddi heart_block5_m_2_3_dff_m mbk_sig502 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2203 mbk_sig505 heart_block5_ck2 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2204 heart_block5_m_2_3_dff_s mbk_sig507 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2205 vddi heart_block5_m_2_3_dff_s mbk_sig507 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2206 heart_block5_s32 heart_block5_m_2_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2207 heart_block5_m_2_3_dff_m mbk_sig502 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2208 mbk_sig501 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2209 mbk_sig476 heart_block1_ssa0 vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M2210 mbk_sig465 heart_block1_ssd0 mbk_sig476 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M2211 vddi mbk_sig465 heart_r_0 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2212 vddi heart_block2_selray heart_block2_selaluy vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2213 mbk_sig475 heart_block2_syra1 vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M2214 mbk_sig463 heart_block2_syalu1 mbk_sig475 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M2215 vddi mbk_sig463 yc_1 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2216 vddi mbk_sig461 heart_block2_syra1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2217 vddi heart_ra_1 mbk_sig461 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2218 mbk_sig461 heart_block2_selray vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2219 vddi mbk_sig458 heart_block2_syalu1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2220 vddi heart_block2_a26ms_i0 mbk_sig458 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2221 mbk_sig458 heart_block2_selaluy vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2222 vddi mbk_sig455 heart_block1_ssa0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2223 vddi heart_ra_0 mbk_sig455 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2224 mbk_sig455 heart_block1_selar vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2225 vddi mbk_sig453 heart_block5_enable vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2226 vddi cko mbk_sig453 vddi TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
M2227 mbk_sig453 heart_block5_wram vddi vddi TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M2228 vddi mbk_sig450 heart_block1_sra1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2229 vddi heart_ra_1 mbk_sig450 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2230 mbk_sig450 heart_block1_selas vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2231 vddi mbk_sig446 heart_block5_wram vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2232 vddi heart_fonc_mode mbk_sig446 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2233 mbk_sig446 heart_block5_o21s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2234 mbk_sig473 heart_r_2 mbk_sig443 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2235 vddi heart_block3_n0 mbk_sig473 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2236 vddi heart_block3_n0 mbk_sig474 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2237 mbk_sig474 heart_r_2 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M2238 heart_block3_x02 mbk_sig443 mbk_sig474 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2239 vddi mbk_sig440 heart_block1_sra3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2240 vddi heart_ra_3 mbk_sig440 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2241 mbk_sig440 heart_block1_selas vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2242 mbk_sig472 ii_8 vddi vddi TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
M2243 mbk_sig437 ii_7 mbk_sig472 vddi TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
M2244 vddi mbk_sig437 heart_block5_o21s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2245 vddi mbk_sig436 heart_block1_srq2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2246 vddi heart_q_2 mbk_sig436 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2247 mbk_sig436 heart_block1_selqs vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2248 vddi mbk_sig433 heart_block1_ssa3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2249 vddi heart_ra_3 mbk_sig433 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2250 mbk_sig433 heart_block1_selar vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2251 mbk_sig471 heart_block1_sra2 mbk_sig470 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M2252 mbk_sig430 heart_block1_srq2 mbk_sig471 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M2253 vddi mbk_sig430 heart_s_2 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2254 mbk_sig470 heart_block1_srb2 vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M2255 vddi mbk_sig428 heart_block1_sra2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2256 vddi heart_ra_2 mbk_sig428 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2257 mbk_sig428 heart_block1_selas vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2258 mbk_sig422 mbk_sig424 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2259 vddi heart_block5_m_13_3_dff_m mbk_sig424 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2260 mbk_sig423 heart_block5_ck13 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2261 heart_block5_m_13_3_dff_s mbk_sig426 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2262 vddi heart_block5_m_13_3_dff_s mbk_sig426 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2263 heart_block5_s313 heart_block5_m_13_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2264 heart_block5_m_13_3_dff_m mbk_sig424 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2265 mbk_sig419 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2266 vddi mbk_sig416 heart_block4_test_mode vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2267 vddi testi mbk_sig416 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2268 mbk_sig416 heart_block4_n14s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2269 vddi testi heart_block4_n15s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2270 mbk_sig410 mbk_sig405 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2271 vddi heart_block5_m_16_0_dff_m mbk_sig405 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2272 mbk_sig412 heart_block5_ck16 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2273 heart_block5_m_16_0_dff_s mbk_sig411 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2274 vddi heart_block5_m_16_0_dff_s mbk_sig411 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2275 heart_block5_s016 heart_block5_m_16_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2276 heart_block5_m_16_0_dff_m mbk_sig405 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2277 mbk_sig407 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2278 heart_block5_b016s heart_block5_s016 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2279 vddi heart_block5_b16 heart_block5_b016s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2280 heart_block5_a116s heart_block5_s116 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2281 vddi heart_block5_a16 heart_block5_a116s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2282 heart_block5_a016s heart_block5_s016 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2283 vddi heart_block5_a16 heart_block5_a016s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2284 vddi mbk_sig396 heart_block5_oa411s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2285 vddi heart_block5_a114s mbk_sig396 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2286 mbk_sig396 heart_block5_a115s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2287 vddi heart_block5_a116s mbk_sig396 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2288 mbk_sig396 heart_block5_a113s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2289 mbk_sig387 mbk_sig383 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2290 vddi heart_block5_m_14_2_dff_m mbk_sig383 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2291 mbk_sig385 heart_block5_ck14 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2292 heart_block5_m_14_2_dff_s mbk_sig388 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2293 vddi heart_block5_m_14_2_dff_s mbk_sig388 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2294 heart_block5_s214 heart_block5_m_14_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2295 heart_block5_m_14_2_dff_m mbk_sig383 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2296 mbk_sig382 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2297 vddi mbk_sig381 heart_block5_ck14 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2298 vddi heart_block5_enable mbk_sig381 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2299 mbk_sig381 heart_block5_b14 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2300 heart_block5_a314s heart_block5_s314 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2301 vddi heart_block5_a14 heart_block5_a314s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2302 mbk_sig373 mbk_sig375 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2303 vddi heart_block5_m_9_0_dff_m mbk_sig375 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2304 mbk_sig374 heart_block5_ck9 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2305 heart_block5_m_9_0_dff_s mbk_sig378 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2306 vddi heart_block5_m_9_0_dff_s mbk_sig378 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2307 heart_block5_s09 heart_block5_m_9_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2308 heart_block5_m_9_0_dff_m mbk_sig375 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2309 mbk_sig370 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2310 vddi mbk_sig369 heart_block5_oa410s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2311 vddi heart_block5_a014s mbk_sig369 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2312 mbk_sig369 heart_block5_a015s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2313 vddi heart_block5_a016s mbk_sig369 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2314 mbk_sig369 heart_block5_a013s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2315 heart_block5_a114s heart_block5_s114 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2316 vddi heart_block5_a14 heart_block5_a114s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2317 vddi heart_a_2 heart_block5_na2 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2318 mbk_sig361 mbk_sig356 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2319 vddi heart_block5_m_9_1_dff_m mbk_sig356 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2320 mbk_sig358 heart_block5_ck9 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2321 heart_block5_m_9_1_dff_s mbk_sig362 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2322 vddi heart_block5_m_9_1_dff_s mbk_sig362 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2323 heart_block5_s19 heart_block5_m_9_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2324 heart_block5_m_9_1_dff_m mbk_sig356 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2325 mbk_sig355 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2326 heart_block5_b09s heart_block5_s09 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2327 vddi heart_block5_b9 heart_block5_b09s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2328 heart_block5_a215s heart_block5_s215 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2329 vddi heart_block5_a15 heart_block5_a215s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2330 heart_block5_b19s heart_block5_s19 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2331 vddi heart_block5_b9 heart_block5_b19s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2332 mbk_sig347 mbk_sig343 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2333 vddi heart_block5_m_11_1_dff_m mbk_sig343 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2334 mbk_sig345 heart_block5_ck11 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2335 heart_block5_m_11_1_dff_s mbk_sig348 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2336 vddi heart_block5_m_11_1_dff_s mbk_sig348 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2337 heart_block5_s111 heart_block5_m_11_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2338 heart_block5_m_11_1_dff_m mbk_sig343 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2339 mbk_sig342 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2340 vddi mbk_sig338 heart_block5_ob421s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2341 vddi heart_block5_b110s mbk_sig338 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2342 mbk_sig338 heart_block5_b111s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2343 vddi heart_block5_b112s mbk_sig338 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2344 mbk_sig338 heart_block5_b19s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2345 vddi mbk_sig332 heart_block5_a15 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2346 vddi heart_a_1 mbk_sig332 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2347 mbk_sig332 heart_a_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2348 vddi heart_a_3 mbk_sig332 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2349 mbk_sig332 heart_block5_na0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2350 heart_block5_a211s heart_block5_s211 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2351 vddi heart_block5_a11 heart_block5_a211s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2352 vddi mbk_sig326 heart_block5_a9 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2353 vddi heart_block5_na1 mbk_sig326 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2354 mbk_sig326 heart_block5_na2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2355 vddi heart_a_3 mbk_sig326 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2356 mbk_sig326 heart_block5_na0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2357 heart_block5_a011s heart_block5_s011 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2358 vddi heart_block5_a11 heart_block5_a011s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2359 vddi mbk_sig321 heart_block5_oa420s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2360 vddi heart_block5_a010s mbk_sig321 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2361 mbk_sig321 heart_block5_a011s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2362 vddi heart_block5_a012s mbk_sig321 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2363 mbk_sig321 heart_block5_a09s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2364 heart_block5_a19s heart_block5_s19 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2365 vddi heart_block5_a9 heart_block5_a19s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2366 heart_block5_a09s heart_block5_s09 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2367 vddi heart_block5_a9 heart_block5_a09s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2368 vddi mbk_sig309 heart_block5_a12 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2369 vddi heart_a_1 mbk_sig309 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2370 mbk_sig309 heart_block5_na2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2371 vddi heart_a_3 mbk_sig309 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2372 mbk_sig309 heart_a_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2373 vddi mbk_sig303 heart_block5_oa421s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2374 vddi heart_block5_a110s mbk_sig303 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2375 mbk_sig303 heart_block5_a111s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2376 vddi heart_block5_a112s mbk_sig303 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2377 mbk_sig303 heart_block5_a19s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2378 mbk_sig297 mbk_sig299 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2379 vddi heart_block5_m_12_2_dff_m mbk_sig299 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2380 mbk_sig298 heart_block5_ck12 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2381 heart_block5_m_12_2_dff_s mbk_sig302 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2382 vddi heart_block5_m_12_2_dff_s mbk_sig302 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2383 heart_block5_s212 heart_block5_m_12_2_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2384 heart_block5_m_12_2_dff_m mbk_sig299 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2385 mbk_sig293 heart_block5_shram2 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2386 heart_block5_a310s heart_block5_s310 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2387 vddi heart_block5_a10 heart_block5_a310s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2388 heart_block5_b110s heart_block5_s110 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2389 vddi heart_block5_b10 heart_block5_b110s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2390 heart_block5_a012s heart_block5_s012 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2391 vddi heart_block5_a12 heart_block5_a012s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2392 heart_block5_a110s heart_block5_s110 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2393 vddi heart_block5_a10 heart_block5_a110s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2394 vddi mbk_sig264 heart_block1_ssd0 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2395 vddi heart_d_0 mbk_sig264 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2396 mbk_sig264 heart_block1_seldr vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2397 vddi ii_2 heart_block1_ni2 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2398 vddi mbk_sig262 heart_block1_selas vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2399 vddi heart_block1_ni1 mbk_sig262 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2400 mbk_sig262 ii_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2401 vddi mbk_sig259 heart_block1_selar vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2402 vddi heart_block1_ni2 mbk_sig259 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2403 mbk_sig259 heart_block1_ni1 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2404 vddi ii_1 heart_block1_ni1 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2405 mbk_sig258 heart_block1_ssa3 vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M2406 mbk_sig257 heart_block1_ssd3 mbk_sig258 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M2407 vddi mbk_sig257 heart_r_3 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2408 vddi mbk_sig256 heart_block1_seldr vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2409 vddi heart_block1_o22s mbk_sig256 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2410 mbk_sig256 ii_2 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2411 vddi mbk_sig254 heart_block1_ssd2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2412 vddi heart_d_2 mbk_sig254 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2413 mbk_sig254 heart_block1_seldr vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2414 mbk_sig252 heart_block1_ssa2 vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M2415 mbk_sig251 heart_block1_ssd2 mbk_sig252 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M2416 vddi mbk_sig251 heart_r_2 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2417 mbk_sig248 heart_r_1 mbk_sig247 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2418 vddi heart_block3_n0 mbk_sig248 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2419 vddi heart_block3_n0 mbk_sig250 vddi TP L=0.18U W=4.14U AS=1.4904P 
+ AD=1.4904P PS=9U PD=9U 
M2420 mbk_sig250 heart_r_1 vddi vddi TP L=0.18U W=4.14U AS=1.4904P AD=1.4904P 
+ PS=9U PD=9U 
M2421 heart_block3_x01 mbk_sig247 mbk_sig250 vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2422 mbk_sig246 ii_1 vddi vddi TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
M2423 mbk_sig244 ii_0 mbk_sig246 vddi TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
M2424 vddi mbk_sig244 heart_block1_o22s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2425 vddi mbk_sig243 heart_block2_syra2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2426 vddi heart_ra_2 mbk_sig243 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2427 mbk_sig243 heart_block2_selray vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2428 mbk_sig242 heart_block2_syra2 vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M2429 mbk_sig241 heart_block2_syalu2 mbk_sig242 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M2430 vddi mbk_sig241 yc_2 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2431 mbk_sig240 ii_1 vddi vddi TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
M2432 mbk_sig239 heart_block1_ni2 mbk_sig240 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M2433 vddi mbk_sig239 heart_block1_o21s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2434 vddi mbk_sig238 heart_block1_ssa2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2435 vddi heart_ra_2 mbk_sig238 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2436 mbk_sig238 heart_block1_selar vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2437 vddi mbk_sig236 heart_block1_ssd3 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2438 vddi heart_d_3 mbk_sig236 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2439 mbk_sig236 heart_block1_seldr vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2440 vddi ii_6 heart_block2_ni6 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2441 mbk_sig234 ii_7 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2442 vddi heart_block2_ni6 mbk_sig234 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2443 mbk_sig234 heart_block2_ni8 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2444 vddi mbk_sig234 heart_block2_selray vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2445 vddi ii_8 heart_block2_ni8 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2446 vddi mbk_sig230 heart_block1_ssa1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2447 vddi heart_ra_1 mbk_sig230 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2448 mbk_sig230 heart_block1_selar vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2449 mbk_sig229 heart_block1_ssa1 vddi vddi TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
M2450 mbk_sig228 heart_block1_ssd1 mbk_sig229 vddi TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
M2451 vddi mbk_sig228 heart_r_1 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2452 vddi mbk_sig227 heart_block1_ssd1 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2453 vddi heart_d_1 mbk_sig227 vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2454 mbk_sig227 heart_block1_seldr vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2455 vddi mbk_sig224 heart_block1_selqs vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2456 vddi heart_block1_o21s mbk_sig224 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2457 mbk_sig224 heart_block1_ni0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2458 vddi ii_0 heart_block1_ni0 vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2459 vddi mbk_sig223 heart_block1_selbs vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2460 vddi heart_block1_ni2 mbk_sig223 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2461 mbk_sig223 ii_0 vddi vddi TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M2462 heart_block5_a014s heart_block5_s014 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2463 vddi heart_block5_a14 heart_block5_a014s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2464 heart_block5_b014s heart_block5_s014 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2465 vddi heart_block5_b14 heart_block5_b014s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2466 mbk_sig218 mbk_sig147 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2467 vddi heart_block5_m_14_0_dff_m mbk_sig147 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2468 mbk_sig219 heart_block5_ck14 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2469 heart_block5_m_14_0_dff_s mbk_sig149 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2470 vddi heart_block5_m_14_0_dff_s mbk_sig149 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2471 heart_block5_s014 heart_block5_m_14_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2472 heart_block5_m_14_0_dff_m mbk_sig147 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2473 mbk_sig217 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2474 mbk_sig216 mbk_sig143 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2475 vddi heart_block5_m_14_1_dff_m mbk_sig143 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2476 mbk_sig215 heart_block5_ck14 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2477 heart_block5_m_14_1_dff_s mbk_sig145 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2478 vddi heart_block5_m_14_1_dff_s mbk_sig145 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2479 heart_block5_s114 heart_block5_m_14_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2480 heart_block5_m_14_1_dff_m mbk_sig143 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2481 mbk_sig214 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2482 heart_block5_b015s heart_block5_s015 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2483 vddi heart_block5_b15 heart_block5_b015s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2484 heart_block5_b314s heart_block5_s314 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2485 vddi heart_block5_b14 heart_block5_b314s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2486 heart_block5_a015s heart_block5_s015 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2487 vddi heart_block5_a15 heart_block5_a015s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2488 heart_ra_2 heart_block5_oa442s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2489 vddi heart_block5_oa432s heart_ra_2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2490 heart_ra_2 heart_block5_oa422s vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2491 vddi heart_block5_oa412s heart_ra_2 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2492 mbk_sig210 mbk_sig125 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2493 vddi heart_block5_m_14_3_dff_m mbk_sig125 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2494 mbk_sig209 heart_block5_ck14 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2495 heart_block5_m_14_3_dff_s mbk_sig128 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2496 vddi heart_block5_m_14_3_dff_s mbk_sig128 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2497 heart_block5_s314 heart_block5_m_14_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2498 heart_block5_m_14_3_dff_m mbk_sig125 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2499 mbk_sig208 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2500 heart_block5_b011s heart_block5_s011 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2501 vddi heart_block5_b11 heart_block5_b011s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2502 heart_block5_b114s heart_block5_s114 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2503 vddi heart_block5_b14 heart_block5_b114s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2504 mbk_sig204 mbk_sig115 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2505 vddi heart_block5_m_15_0_dff_m mbk_sig115 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2506 mbk_sig205 heart_block5_ck15 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2507 heart_block5_m_15_0_dff_s mbk_sig119 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2508 vddi heart_block5_m_15_0_dff_s mbk_sig119 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2509 heart_block5_s015 heart_block5_m_15_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2510 heart_block5_m_15_0_dff_m mbk_sig115 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2511 mbk_sig203 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2512 mbk_sig201 mbk_sig110 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2513 vddi heart_block5_m_11_0_dff_m mbk_sig110 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2514 mbk_sig202 heart_block5_ck11 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2515 heart_block5_m_11_0_dff_s mbk_sig113 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2516 vddi heart_block5_m_11_0_dff_s mbk_sig113 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2517 heart_block5_s011 heart_block5_m_11_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2518 heart_block5_m_11_0_dff_m mbk_sig110 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2519 mbk_sig200 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2520 heart_block5_b111s heart_block5_s111 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2521 vddi heart_block5_b11 heart_block5_b111s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2522 vddi mbk_sig105 heart_block5_ob420s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2523 vddi heart_block5_b010s mbk_sig105 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2524 mbk_sig105 heart_block5_b011s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2525 vddi heart_block5_b012s mbk_sig105 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2526 mbk_sig105 heart_block5_b09s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2527 mbk_sig197 mbk_sig94 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2528 vddi heart_block5_m_12_3_dff_m mbk_sig94 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2529 mbk_sig198 heart_block5_ck12 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2530 heart_block5_m_12_3_dff_s mbk_sig97 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2531 vddi heart_block5_m_12_3_dff_s mbk_sig97 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2532 heart_block5_s312 heart_block5_m_12_3_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2533 heart_block5_m_12_3_dff_m mbk_sig94 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2534 mbk_sig196 heart_block5_shram3 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2535 vddi mbk_sig88 heart_block5_oa422s vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2536 vddi heart_block5_a210s mbk_sig88 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2537 mbk_sig88 heart_block5_a211s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2538 vddi heart_block5_a212s mbk_sig88 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2539 mbk_sig88 heart_block5_a29s vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2540 heart_block5_a29s heart_block5_s29 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2541 vddi heart_block5_a9 heart_block5_a29s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2542 mbk_sig193 mbk_sig79 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2543 vddi heart_block5_m_12_0_dff_m mbk_sig79 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2544 mbk_sig194 heart_block5_ck12 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2545 heart_block5_m_12_0_dff_s mbk_sig82 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2546 vddi heart_block5_m_12_0_dff_s mbk_sig82 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2547 heart_block5_s012 heart_block5_m_12_0_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2548 heart_block5_m_12_0_dff_m mbk_sig79 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2549 mbk_sig192 heart_block5_shram0 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2550 heart_block5_b012s heart_block5_s012 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2551 vddi heart_block5_b12 heart_block5_b012s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2552 heart_block5_a111s heart_block5_s111 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2553 vddi heart_block5_a11 heart_block5_a111s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2554 heart_block5_a112s heart_block5_s112 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2555 vddi heart_block5_a12 heart_block5_a112s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2556 heart_block5_b112s heart_block5_s112 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2557 vddi heart_block5_b12 heart_block5_b112s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2558 mbk_sig186 mbk_sig67 vddi vddi TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M2559 vddi heart_block5_m_12_1_dff_m mbk_sig67 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2560 mbk_sig187 heart_block5_ck12 vddi vddi TP L=0.18U W=3.24U AS=1.1664P 
+ AD=1.1664P PS=7.2U PD=7.2U 
M2561 heart_block5_m_12_1_dff_s mbk_sig69 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2562 vddi heart_block5_m_12_1_dff_s mbk_sig69 vddi TP L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M2563 heart_block5_s112 heart_block5_m_12_1_dff_s vddi vddi TP L=0.18U W=4.14U 
+ AS=1.4904P AD=1.4904P PS=9U PD=9U 
M2564 heart_block5_m_12_1_dff_m mbk_sig67 vddi vddi TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
M2565 mbk_sig184 heart_block5_shram1 vddi vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2566 vddi mbk_sig183 heart_block5_ck12 vddi TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M2567 vddi heart_block5_enable mbk_sig183 vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2568 mbk_sig183 heart_block5_b12 vddi vddi TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M2569 heart_block5_a212s heart_block5_s212 vddi vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2570 vddi heart_block5_a12 heart_block5_a212s vddi TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M2571 vsse mbk_sig55 signe vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2572 signe mbk_sig55 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2573 vsse mbk_sig55 signe vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2574 signe mbk_sig55 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2575 vsse mbk_sig55 signe vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2576 signe mbk_sig55 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2577 vsse mbk_sig55 signe vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2578 signe mbk_sig55 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2579 vsse mbk_sig55 signe vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2580 signe mbk_sig55 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2581 vsse mbk_sig55 signe vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2582 signe mbk_sig55 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2583 vsse mbk_sig55 signe vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2584 signe mbk_sig55 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2585 vsse mbk_sig55 signe vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2586 signe mbk_sig55 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2587 vsse mbk_sig55 signe vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2588 signe mbk_sig55 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2589 vsse mbk_sig55 signe vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2590 signe mbk_sig55 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2591 vsse mbk_sig55 signe vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2592 signe mbk_sig55 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2593 vsse mbk_sig55 signe vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2594 signe mbk_sig55 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2595 vssi mbk_sig178 mbk_sig55 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2596 mbk_sig55 mbk_sig178 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2597 vssi mbk_sig178 mbk_sig55 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2598 mbk_sig55 mbk_sig178 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2599 vssi mbk_sig179 mbk_sig178 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2600 mbk_sig179 signec vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2601 vsse mbk_sig467 ovr vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2602 ovr mbk_sig467 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2603 vsse mbk_sig467 ovr vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2604 ovr mbk_sig467 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2605 vsse mbk_sig467 ovr vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2606 ovr mbk_sig467 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2607 vsse mbk_sig467 ovr vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2608 ovr mbk_sig467 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2609 vsse mbk_sig467 ovr vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2610 ovr mbk_sig467 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2611 vsse mbk_sig467 ovr vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2612 ovr mbk_sig467 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2613 vsse mbk_sig467 ovr vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2614 ovr mbk_sig467 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2615 vsse mbk_sig467 ovr vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2616 ovr mbk_sig467 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2617 vsse mbk_sig467 ovr vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2618 ovr mbk_sig467 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2619 vsse mbk_sig467 ovr vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2620 ovr mbk_sig467 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2621 vsse mbk_sig467 ovr vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2622 ovr mbk_sig467 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2623 vsse mbk_sig467 ovr vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2624 ovr mbk_sig467 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2625 vssi mbk_sig478 mbk_sig467 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2626 mbk_sig467 mbk_sig478 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2627 vssi mbk_sig478 mbk_sig467 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2628 mbk_sig467 mbk_sig478 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2629 vssi mbk_sig479 mbk_sig478 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2630 mbk_sig479 ovrc vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2631 vsse mbk_sig682 cout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2632 cout mbk_sig682 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2633 vsse mbk_sig682 cout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2634 cout mbk_sig682 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2635 vsse mbk_sig682 cout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2636 cout mbk_sig682 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2637 vsse mbk_sig682 cout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2638 cout mbk_sig682 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2639 vsse mbk_sig682 cout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2640 cout mbk_sig682 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2641 vsse mbk_sig682 cout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2642 cout mbk_sig682 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2643 vsse mbk_sig682 cout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2644 cout mbk_sig682 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2645 vsse mbk_sig682 cout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2646 cout mbk_sig682 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2647 vsse mbk_sig682 cout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2648 cout mbk_sig682 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2649 vsse mbk_sig682 cout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2650 cout mbk_sig682 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2651 vsse mbk_sig682 cout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2652 cout mbk_sig682 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2653 vsse mbk_sig682 cout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2654 cout mbk_sig682 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2655 vssi mbk_sig687 mbk_sig682 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2656 mbk_sig682 mbk_sig687 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2657 vssi mbk_sig687 mbk_sig682 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2658 mbk_sig682 mbk_sig687 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2659 vssi mbk_sig686 mbk_sig687 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2660 mbk_sig686 coutc vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2661 vsse mbk_sig871 zero vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2662 zero mbk_sig871 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2663 vsse mbk_sig871 zero vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2664 zero mbk_sig871 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2665 vsse mbk_sig871 zero vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2666 zero mbk_sig871 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2667 vsse mbk_sig871 zero vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2668 zero mbk_sig871 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2669 vsse mbk_sig871 zero vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2670 zero mbk_sig871 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2671 vsse mbk_sig871 zero vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2672 zero mbk_sig871 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2673 vsse mbk_sig871 zero vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2674 zero mbk_sig871 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2675 vsse mbk_sig871 zero vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2676 zero mbk_sig871 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2677 vsse mbk_sig871 zero vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2678 zero mbk_sig871 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2679 vsse mbk_sig871 zero vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2680 zero mbk_sig871 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2681 vsse mbk_sig871 zero vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2682 zero mbk_sig871 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2683 vsse mbk_sig871 zero vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2684 zero mbk_sig871 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2685 vssi mbk_sig878 mbk_sig871 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2686 mbk_sig871 mbk_sig878 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2687 vssi mbk_sig878 mbk_sig871 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2688 mbk_sig871 mbk_sig878 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2689 vssi mbk_sig879 mbk_sig878 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2690 mbk_sig879 zeroc vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2691 fonc vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2692 vsse vsse fonc vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2693 fonc vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2694 vsse vsse fonc vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2695 vssi fonc mbk_sig1066 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2696 mbk_sig1066 fonc vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2697 vssi fonc mbk_sig1066 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2698 vssi mbk_sig1066 fonci vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2699 fonci mbk_sig1066 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2700 test vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2701 vsse vsse test vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2702 test vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2703 vsse vsse test vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2704 vssi test mbk_sig1271 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2705 mbk_sig1271 test vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2706 vssi test mbk_sig1271 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2707 vssi mbk_sig1271 testi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2708 testi mbk_sig1271 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2709 scin vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2710 vsse vsse scin vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2711 scin vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2712 vsse vsse scin vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2713 vssi scin mbk_sig1466 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2714 mbk_sig1466 scin vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2715 vssi scin mbk_sig1466 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2716 vssi mbk_sig1466 scini vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2717 scini mbk_sig1466 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2718 q0 mbk_sig1639 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2719 vsse mbk_sig1639 q0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2720 q0 mbk_sig1639 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2721 vsse mbk_sig1639 q0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2722 vsse mbk_sig1639 q0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2723 q0 mbk_sig1639 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2724 vsse mbk_sig1639 q0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2725 q0 mbk_sig1639 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2726 vsse mbk_sig1639 q0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2727 q0 mbk_sig1639 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2728 vsse mbk_sig1639 q0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2729 q0 mbk_sig1639 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2730 vsse mbk_sig1639 q0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2731 q0 mbk_sig1639 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2732 vsse mbk_sig1639 q0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2733 q0 mbk_sig1639 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2734 vsse mbk_sig1639 q0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2735 q0 mbk_sig1639 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2736 vsse mbk_sig1639 q0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2737 q0 mbk_sig1639 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2738 vsse mbk_sig1639 q0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2739 q0 mbk_sig1639 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2740 vsse mbk_sig1639 q0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2741 q0 mbk_sig1639 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2742 mbk_sig1636 q0 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2743 vssi q0 mbk_sig1636 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2744 vssi mbk_sig1636 q0i vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2745 q0i mbk_sig1636 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2746 vssi q0 mbk_sig1636 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2747 vssi mbk_sig1652 mbk_sig1639 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2748 mbk_sig1639 mbk_sig1652 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2749 mbk_sig1647 f0c vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2750 vssi mbk_sig1652 mbk_sig1639 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2751 mbk_sig1639 mbk_sig1652 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2752 vssi mbk_sig1647 mbk_sig1646 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2753 mbk_sig1639 mbk_sig1646 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2754 vssi mbk_sig1646 mbk_sig1639 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2755 mbk_sig1639 mbk_sig1646 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2756 vssi mbk_sig1646 mbk_sig1639 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2757 mbk_sig1639 mbk_sig1653 mbk_sig1638 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2758 mbk_sig1638 mbk_sig1653 mbk_sig1639 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2759 mbk_sig1639 mbk_sig1653 mbk_sig1638 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2760 mbk_sig1638 mbk_sig1653 mbk_sig1639 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2761 mbk_sig1652 decaldc vssi vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
M2762 vssi mbk_sig1652 mbk_sig1653 vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
M2763 q3 mbk_sig1818 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2764 vsse mbk_sig1818 q3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2765 q3 mbk_sig1818 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2766 vsse mbk_sig1818 q3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2767 vsse mbk_sig1818 q3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2768 q3 mbk_sig1818 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2769 vsse mbk_sig1818 q3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2770 q3 mbk_sig1818 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2771 vsse mbk_sig1818 q3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2772 q3 mbk_sig1818 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2773 vsse mbk_sig1818 q3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2774 q3 mbk_sig1818 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2775 vsse mbk_sig1818 q3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2776 q3 mbk_sig1818 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2777 vsse mbk_sig1818 q3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2778 q3 mbk_sig1818 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2779 vsse mbk_sig1818 q3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2780 q3 mbk_sig1818 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2781 vsse mbk_sig1818 q3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2782 q3 mbk_sig1818 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2783 vsse mbk_sig1818 q3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2784 q3 mbk_sig1818 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2785 vsse mbk_sig1818 q3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2786 q3 mbk_sig1818 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2787 mbk_sig1815 q3 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2788 vssi q3 mbk_sig1815 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2789 vssi mbk_sig1815 q3i vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2790 q3i mbk_sig1815 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2791 vssi q3 mbk_sig1815 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2792 vssi mbk_sig1835 mbk_sig1818 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2793 mbk_sig1818 mbk_sig1835 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2794 mbk_sig1827 f3c vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2795 vssi mbk_sig1835 mbk_sig1818 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2796 mbk_sig1818 mbk_sig1835 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2797 vssi mbk_sig1827 mbk_sig1826 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2798 mbk_sig1818 mbk_sig1826 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2799 vssi mbk_sig1826 mbk_sig1818 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2800 mbk_sig1818 mbk_sig1826 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2801 vssi mbk_sig1826 mbk_sig1818 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2802 mbk_sig1818 mbk_sig1836 mbk_sig1817 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2803 mbk_sig1817 mbk_sig1836 mbk_sig1818 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2804 mbk_sig1818 mbk_sig1836 mbk_sig1817 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2805 mbk_sig1817 mbk_sig1836 mbk_sig1818 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2806 mbk_sig1835 decalgc vssi vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
M2807 vssi mbk_sig1835 mbk_sig1836 vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
M2808 cin vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2809 vsse vsse cin vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2810 cin vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2811 vsse vsse cin vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2812 vssi cin mbk_sig44 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2813 mbk_sig44 cin vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2814 vssi cin mbk_sig44 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2815 vssi mbk_sig44 cini vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2816 cini mbk_sig44 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M2817 vsse mbk_sig57 np vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2818 np mbk_sig57 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2819 vsse mbk_sig57 np vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2820 np mbk_sig57 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2821 vsse mbk_sig57 np vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2822 np mbk_sig57 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2823 vsse mbk_sig57 np vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2824 np mbk_sig57 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2825 vsse mbk_sig57 np vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2826 np mbk_sig57 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2827 vsse mbk_sig57 np vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2828 np mbk_sig57 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2829 vsse mbk_sig57 np vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2830 np mbk_sig57 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2831 vsse mbk_sig57 np vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2832 np mbk_sig57 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2833 vsse mbk_sig57 np vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2834 np mbk_sig57 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2835 vsse mbk_sig57 np vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2836 np mbk_sig57 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2837 vsse mbk_sig57 np vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2838 np mbk_sig57 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2839 vsse mbk_sig57 np vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2840 np mbk_sig57 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2841 vssi mbk_sig265 mbk_sig57 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2842 mbk_sig57 mbk_sig265 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2843 vssi mbk_sig265 mbk_sig57 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2844 mbk_sig57 mbk_sig265 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2845 vssi mbk_sig180 mbk_sig265 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2846 mbk_sig180 npc vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2847 vsse mbk_sig469 ng vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2848 ng mbk_sig469 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2849 vsse mbk_sig469 ng vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2850 ng mbk_sig469 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2851 vsse mbk_sig469 ng vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2852 ng mbk_sig469 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2853 vsse mbk_sig469 ng vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2854 ng mbk_sig469 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2855 vsse mbk_sig469 ng vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2856 ng mbk_sig469 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2857 vsse mbk_sig469 ng vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2858 ng mbk_sig469 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2859 vsse mbk_sig469 ng vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2860 ng mbk_sig469 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2861 vsse mbk_sig469 ng vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2862 ng mbk_sig469 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2863 vsse mbk_sig469 ng vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2864 ng mbk_sig469 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2865 vsse mbk_sig469 ng vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2866 ng mbk_sig469 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2867 vsse mbk_sig469 ng vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2868 ng mbk_sig469 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2869 vsse mbk_sig469 ng vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2870 ng mbk_sig469 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2871 vssi mbk_sig480 mbk_sig469 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2872 mbk_sig469 mbk_sig480 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2873 vssi mbk_sig480 mbk_sig469 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2874 mbk_sig469 mbk_sig480 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2875 vssi mbk_sig481 mbk_sig480 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2876 mbk_sig481 ngc vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2877 r0 mbk_sig669 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2878 vsse mbk_sig669 r0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2879 r0 mbk_sig669 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2880 vsse mbk_sig669 r0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2881 vsse mbk_sig669 r0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2882 r0 mbk_sig669 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2883 vsse mbk_sig669 r0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2884 r0 mbk_sig669 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2885 vsse mbk_sig669 r0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2886 r0 mbk_sig669 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2887 vsse mbk_sig669 r0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2888 r0 mbk_sig669 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2889 vsse mbk_sig669 r0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2890 r0 mbk_sig669 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2891 vsse mbk_sig669 r0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2892 r0 mbk_sig669 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2893 vsse mbk_sig669 r0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2894 r0 mbk_sig669 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2895 vsse mbk_sig669 r0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2896 r0 mbk_sig669 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2897 vsse mbk_sig669 r0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2898 r0 mbk_sig669 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2899 vsse mbk_sig669 r0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2900 r0 mbk_sig669 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2901 mbk_sig671 r0 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2902 vssi r0 mbk_sig671 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2903 vssi mbk_sig671 r0i vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2904 r0i mbk_sig671 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2905 vssi r0 mbk_sig671 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2906 vssi mbk_sig690 mbk_sig669 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2907 mbk_sig669 mbk_sig690 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2908 mbk_sig683 s0c vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2909 vssi mbk_sig690 mbk_sig669 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2910 mbk_sig669 mbk_sig690 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2911 vssi mbk_sig683 mbk_sig688 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2912 mbk_sig669 mbk_sig688 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2913 vssi mbk_sig688 mbk_sig669 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2914 mbk_sig669 mbk_sig688 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2915 vssi mbk_sig688 mbk_sig669 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2916 mbk_sig669 mbk_sig689 mbk_sig670 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2917 mbk_sig670 mbk_sig689 mbk_sig669 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2918 mbk_sig669 mbk_sig689 mbk_sig670 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2919 mbk_sig670 mbk_sig689 mbk_sig669 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2920 mbk_sig690 decaldrc vssi vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
M2921 vssi mbk_sig690 mbk_sig689 vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
M2922 r3 mbk_sig873 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2923 vsse mbk_sig873 r3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2924 r3 mbk_sig873 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2925 vsse mbk_sig873 r3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2926 vsse mbk_sig873 r3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2927 r3 mbk_sig873 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2928 vsse mbk_sig873 r3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2929 r3 mbk_sig873 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2930 vsse mbk_sig873 r3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2931 r3 mbk_sig873 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2932 vsse mbk_sig873 r3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2933 r3 mbk_sig873 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2934 vsse mbk_sig873 r3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2935 r3 mbk_sig873 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2936 vsse mbk_sig873 r3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2937 r3 mbk_sig873 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2938 vsse mbk_sig873 r3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2939 r3 mbk_sig873 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2940 vsse mbk_sig873 r3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2941 r3 mbk_sig873 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2942 vsse mbk_sig873 r3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2943 r3 mbk_sig873 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2944 vsse mbk_sig873 r3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2945 r3 mbk_sig873 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M2946 mbk_sig876 r3 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2947 vssi r3 mbk_sig876 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2948 vssi mbk_sig876 r3i vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2949 r3i mbk_sig876 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2950 vssi r3 mbk_sig876 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2951 vssi mbk_sig885 mbk_sig873 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2952 mbk_sig873 mbk_sig885 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2953 mbk_sig881 s3c vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P PS=11.52U 
+ PD=11.52U 
M2954 vssi mbk_sig885 mbk_sig873 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2955 mbk_sig873 mbk_sig885 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2956 vssi mbk_sig881 mbk_sig880 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2957 mbk_sig873 mbk_sig880 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2958 vssi mbk_sig880 mbk_sig873 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2959 mbk_sig873 mbk_sig880 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2960 vssi mbk_sig880 mbk_sig873 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2961 mbk_sig873 mbk_sig884 mbk_sig874 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2962 mbk_sig874 mbk_sig884 mbk_sig873 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2963 mbk_sig873 mbk_sig884 mbk_sig874 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2964 mbk_sig874 mbk_sig884 mbk_sig873 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2965 mbk_sig885 decalgrc vssi vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
M2966 vssi mbk_sig885 mbk_sig884 vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
M2967 y_0 mbk_sig1075 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2968 vsse mbk_sig1075 y_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2969 y_0 mbk_sig1075 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2970 vsse mbk_sig1075 y_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2971 vsse mbk_sig1075 y_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2972 y_0 mbk_sig1075 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2973 vsse mbk_sig1075 y_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2974 y_0 mbk_sig1075 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2975 vsse mbk_sig1075 y_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2976 y_0 mbk_sig1075 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2977 vsse mbk_sig1075 y_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2978 y_0 mbk_sig1075 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2979 vsse mbk_sig1075 y_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2980 y_0 mbk_sig1075 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2981 vsse mbk_sig1075 y_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2982 y_0 mbk_sig1075 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2983 vsse mbk_sig1075 y_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2984 y_0 mbk_sig1075 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2985 vsse mbk_sig1075 y_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2986 y_0 mbk_sig1075 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2987 vsse mbk_sig1075 y_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2988 y_0 mbk_sig1075 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2989 vsse mbk_sig1075 y_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2990 y_0 mbk_sig1075 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M2991 vssi mbk_sig1224 mbk_sig1223 vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
M2992 mbk_sig1224 oec vssi vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
M2993 mbk_sig1075 mbk_sig1223 mbk_sig1076 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2994 mbk_sig1076 mbk_sig1223 mbk_sig1075 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2995 mbk_sig1075 mbk_sig1223 mbk_sig1076 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2996 mbk_sig1076 mbk_sig1223 mbk_sig1075 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M2997 mbk_sig1075 mbk_sig1084 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2998 vssi mbk_sig1084 mbk_sig1075 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M2999 vssi mbk_sig1085 mbk_sig1084 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3000 mbk_sig1075 mbk_sig1084 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3001 vssi mbk_sig1084 mbk_sig1075 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3002 vssi mbk_sig1224 mbk_sig1075 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3003 mbk_sig1075 mbk_sig1224 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3004 vssi mbk_sig1224 mbk_sig1075 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3005 mbk_sig1075 mbk_sig1224 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3006 mbk_sig1085 yc_0 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3007 y_1 mbk_sig1247 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3008 vsse mbk_sig1247 y_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3009 y_1 mbk_sig1247 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3010 vsse mbk_sig1247 y_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3011 vsse mbk_sig1247 y_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3012 y_1 mbk_sig1247 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3013 vsse mbk_sig1247 y_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3014 y_1 mbk_sig1247 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3015 vsse mbk_sig1247 y_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3016 y_1 mbk_sig1247 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3017 vsse mbk_sig1247 y_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3018 y_1 mbk_sig1247 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3019 vsse mbk_sig1247 y_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3020 y_1 mbk_sig1247 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3021 vsse mbk_sig1247 y_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3022 y_1 mbk_sig1247 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3023 vsse mbk_sig1247 y_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3024 y_1 mbk_sig1247 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3025 vsse mbk_sig1247 y_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3026 y_1 mbk_sig1247 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3027 vsse mbk_sig1247 y_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3028 y_1 mbk_sig1247 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3029 vsse mbk_sig1247 y_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3030 y_1 mbk_sig1247 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3031 vssi mbk_sig1261 mbk_sig1260 vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
M3032 mbk_sig1261 oec vssi vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
M3033 mbk_sig1247 mbk_sig1260 mbk_sig1248 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M3034 mbk_sig1248 mbk_sig1260 mbk_sig1247 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M3035 mbk_sig1247 mbk_sig1260 mbk_sig1248 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M3036 mbk_sig1248 mbk_sig1260 mbk_sig1247 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M3037 mbk_sig1247 mbk_sig1251 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3038 vssi mbk_sig1251 mbk_sig1247 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3039 vssi mbk_sig1250 mbk_sig1251 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3040 mbk_sig1247 mbk_sig1251 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3041 vssi mbk_sig1251 mbk_sig1247 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3042 vssi mbk_sig1261 mbk_sig1247 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3043 mbk_sig1247 mbk_sig1261 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3044 vssi mbk_sig1261 mbk_sig1247 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3045 mbk_sig1247 mbk_sig1261 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3046 mbk_sig1250 yc_1 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3047 y_2 mbk_sig1448 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3048 vsse mbk_sig1448 y_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3049 y_2 mbk_sig1448 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3050 vsse mbk_sig1448 y_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3051 vsse mbk_sig1448 y_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3052 y_2 mbk_sig1448 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3053 vsse mbk_sig1448 y_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3054 y_2 mbk_sig1448 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3055 vsse mbk_sig1448 y_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3056 y_2 mbk_sig1448 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3057 vsse mbk_sig1448 y_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3058 y_2 mbk_sig1448 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3059 vsse mbk_sig1448 y_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3060 y_2 mbk_sig1448 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3061 vsse mbk_sig1448 y_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3062 y_2 mbk_sig1448 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3063 vsse mbk_sig1448 y_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3064 y_2 mbk_sig1448 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3065 vsse mbk_sig1448 y_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3066 y_2 mbk_sig1448 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3067 vsse mbk_sig1448 y_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3068 y_2 mbk_sig1448 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3069 vsse mbk_sig1448 y_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3070 y_2 mbk_sig1448 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3071 vssi mbk_sig1459 mbk_sig1458 vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
M3072 mbk_sig1459 oec vssi vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
M3073 mbk_sig1448 mbk_sig1458 mbk_sig1449 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M3074 mbk_sig1449 mbk_sig1458 mbk_sig1448 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M3075 mbk_sig1448 mbk_sig1458 mbk_sig1449 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M3076 mbk_sig1449 mbk_sig1458 mbk_sig1448 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M3077 mbk_sig1448 mbk_sig1454 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3078 vssi mbk_sig1454 mbk_sig1448 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3079 vssi mbk_sig1450 mbk_sig1454 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3080 mbk_sig1448 mbk_sig1454 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3081 vssi mbk_sig1454 mbk_sig1448 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3082 vssi mbk_sig1459 mbk_sig1448 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3083 mbk_sig1448 mbk_sig1459 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3084 vssi mbk_sig1459 mbk_sig1448 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3085 mbk_sig1448 mbk_sig1459 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3086 mbk_sig1450 yc_2 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3087 y_3 mbk_sig1632 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3088 vsse mbk_sig1632 y_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3089 y_3 mbk_sig1632 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3090 vsse mbk_sig1632 y_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3091 vsse mbk_sig1632 y_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3092 y_3 mbk_sig1632 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3093 vsse mbk_sig1632 y_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3094 y_3 mbk_sig1632 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3095 vsse mbk_sig1632 y_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3096 y_3 mbk_sig1632 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3097 vsse mbk_sig1632 y_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3098 y_3 mbk_sig1632 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3099 vsse mbk_sig1632 y_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3100 y_3 mbk_sig1632 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3101 vsse mbk_sig1632 y_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3102 y_3 mbk_sig1632 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3103 vsse mbk_sig1632 y_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3104 y_3 mbk_sig1632 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3105 vsse mbk_sig1632 y_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3106 y_3 mbk_sig1632 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3107 vsse mbk_sig1632 y_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3108 y_3 mbk_sig1632 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3109 vsse mbk_sig1632 y_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3110 y_3 mbk_sig1632 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3111 vssi mbk_sig1641 mbk_sig1640 vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
M3112 mbk_sig1641 oec vssi vsse TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
M3113 mbk_sig1632 mbk_sig1640 mbk_sig1633 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M3114 mbk_sig1633 mbk_sig1640 mbk_sig1632 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M3115 mbk_sig1632 mbk_sig1640 mbk_sig1633 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M3116 mbk_sig1633 mbk_sig1640 mbk_sig1632 vsse TN L=0.18U W=5.22U AS=1.8792P 
+ AD=1.8792P PS=11.16U PD=11.16U 
M3117 mbk_sig1632 mbk_sig1634 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3118 vssi mbk_sig1634 mbk_sig1632 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3119 vssi mbk_sig1635 mbk_sig1634 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3120 mbk_sig1632 mbk_sig1634 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3121 vssi mbk_sig1634 mbk_sig1632 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3122 vssi mbk_sig1641 mbk_sig1632 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3123 mbk_sig1632 mbk_sig1641 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3124 vssi mbk_sig1641 mbk_sig1632 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3125 mbk_sig1632 mbk_sig1641 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3126 mbk_sig1635 yc_3 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3127 noe vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3128 vsse vsse noe vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3129 noe vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3130 vsse vsse noe vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3131 vssi noe mbk_sig1975 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3132 mbk_sig1975 noe vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3133 vssi noe mbk_sig1975 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3134 vssi mbk_sig1975 noei vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3135 noei mbk_sig1975 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3136 vsse mbk_sig13 scout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3137 scout mbk_sig13 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3138 vsse mbk_sig13 scout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3139 scout mbk_sig13 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3140 vsse mbk_sig13 scout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3141 scout mbk_sig13 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3142 vsse mbk_sig13 scout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3143 scout mbk_sig13 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3144 vsse mbk_sig13 scout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3145 scout mbk_sig13 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3146 vsse mbk_sig13 scout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3147 scout mbk_sig13 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3148 vsse mbk_sig13 scout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3149 scout mbk_sig13 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3150 vsse mbk_sig13 scout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3151 scout mbk_sig13 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3152 vsse mbk_sig13 scout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3153 scout mbk_sig13 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3154 vsse mbk_sig13 scout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3155 scout mbk_sig13 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3156 vsse mbk_sig13 scout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3157 scout mbk_sig13 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3158 vsse mbk_sig13 scout vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3159 scout mbk_sig13 vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P 
+ PS=13.32U PD=13.32U 
M3160 vssi mbk_sig16 mbk_sig13 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3161 mbk_sig13 mbk_sig16 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3162 vssi mbk_sig16 mbk_sig13 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3163 mbk_sig13 mbk_sig16 vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3164 vssi mbk_sig17 mbk_sig16 vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3165 mbk_sig17 scoutc vssi vsse TN L=0.18U W=5.4U AS=1.944P AD=1.944P 
+ PS=11.52U PD=11.52U 
M3166 i_8 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3167 vsse vsse i_8 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3168 i_8 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3169 vsse vsse i_8 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3170 vssi i_8 mbk_sig20 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3171 mbk_sig20 i_8 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3172 vssi i_8 mbk_sig20 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3173 vssi mbk_sig20 ii_8 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3174 ii_8 mbk_sig20 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3175 i_7 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3176 vsse vsse i_7 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3177 i_7 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3178 vsse vsse i_7 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3179 vssi i_7 mbk_sig22 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3180 mbk_sig22 i_7 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3181 vssi i_7 mbk_sig22 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3182 vssi mbk_sig22 ii_7 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3183 ii_7 mbk_sig22 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3184 i_6 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3185 vsse vsse i_6 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3186 i_6 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3187 vsse vsse i_6 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3188 vssi i_6 mbk_sig24 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3189 mbk_sig24 i_6 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3190 vssi i_6 mbk_sig24 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3191 vssi mbk_sig24 ii_6 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3192 ii_6 mbk_sig24 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3193 cko mbk_sig40 vssi vsse TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
M3194 vssi mbk_sig40 cko vsse TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
M3195 cko mbk_sig40 vssi vsse TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
M3196 mbk_sig40 ck_log_log_ck vssi vsse TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
M3197 cko mbk_sig40 vssi vsse TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
M3198 vssi mbk_sig40 cko vsse TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
M3199 i_5 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3200 vsse vsse i_5 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3201 i_5 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3202 vsse vsse i_5 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3203 vssi i_5 mbk_sig26 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3204 mbk_sig26 i_5 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3205 vssi i_5 mbk_sig26 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3206 vssi mbk_sig26 ii_5 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3207 ii_5 mbk_sig26 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3208 i_4 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3209 vsse vsse i_4 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3210 i_4 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3211 vsse vsse i_4 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3212 vssi i_4 mbk_sig28 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3213 mbk_sig28 i_4 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3214 vssi i_4 mbk_sig28 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3215 vssi mbk_sig28 ii_4 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3216 ii_4 mbk_sig28 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3217 i_3 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3218 vsse vsse i_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3219 i_3 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3220 vsse vsse i_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3221 vssi i_3 mbk_sig30 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3222 mbk_sig30 i_3 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3223 vssi i_3 mbk_sig30 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3224 vssi mbk_sig30 ii_3 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3225 ii_3 mbk_sig30 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3226 i_2 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3227 vsse vsse i_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3228 i_2 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3229 vsse vsse i_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3230 vssi i_2 mbk_sig32 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3231 mbk_sig32 i_2 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3232 vssi i_2 mbk_sig32 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3233 vssi mbk_sig32 ii_2 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3234 ii_2 mbk_sig32 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3235 i_1 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3236 vsse vsse i_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3237 i_1 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3238 vsse vsse i_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3239 vssi i_1 mbk_sig34 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3240 mbk_sig34 i_1 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3241 vssi i_1 mbk_sig34 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3242 vssi mbk_sig34 ii_1 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3243 ii_1 mbk_sig34 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3244 i_0 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3245 vsse vsse i_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3246 i_0 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3247 vsse vsse i_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3248 vssi i_0 mbk_sig36 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3249 mbk_sig36 i_0 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3250 vssi i_0 mbk_sig36 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3251 vssi mbk_sig36 ii_0 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3252 ii_0 mbk_sig36 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3253 vsse vsse cke vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3254 cke vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3255 vsse vsse cke vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3256 cke vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3257 vssi mbk_sig38 ck_log_log_ck vsse TN L=0.18U W=4.86U AS=1.7496P 
+ AD=1.7496P PS=10.44U PD=10.44U 
M3258 ck_log_log_ck mbk_sig38 vssi vsse TN L=0.18U W=4.86U AS=1.7496P 
+ AD=1.7496P PS=10.44U PD=10.44U 
M3259 vssi mbk_sig38 ck_log_log_ck vsse TN L=0.18U W=4.86U AS=1.7496P 
+ AD=1.7496P PS=10.44U PD=10.44U 
M3260 vssi mbk_sig38 ck_log_log_ck vsse TN L=0.18U W=4.86U AS=1.7496P 
+ AD=1.7496P PS=10.44U PD=10.44U 
M3261 ck_log_log_ck mbk_sig38 vssi vsse TN L=0.18U W=4.86U AS=1.7496P 
+ AD=1.7496P PS=10.44U PD=10.44U 
M3262 ck_log_log_ck mbk_sig38 vssi vsse TN L=0.18U W=4.86U AS=1.7496P 
+ AD=1.7496P PS=10.44U PD=10.44U 
M3263 vssi mbk_sig38 ck_log_log_ck vsse TN L=0.18U W=4.86U AS=1.7496P 
+ AD=1.7496P PS=10.44U PD=10.44U 
M3264 ck_log_log_ck mbk_sig38 vssi vsse TN L=0.18U W=4.86U AS=1.7496P 
+ AD=1.7496P PS=10.44U PD=10.44U 
M3265 vssi cke mbk_sig38 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3266 mbk_sig38 cke vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3267 vssi cke mbk_sig38 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3268 mbk_sig38 cke vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3269 mbk_sig38 cke vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3270 vssi cke mbk_sig38 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3271 vssi cke mbk_sig38 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3272 vssi cke mbk_sig38 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3273 mbk_sig38 cke vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3274 mbk_sig38 cke vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3275 mbk_sig38 cke vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3276 vssi cke mbk_sig38 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3277 a_3 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3278 vsse vsse a_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3279 a_3 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3280 vsse vsse a_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3281 vssi a_3 mbk_sig1976 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3282 mbk_sig1976 a_3 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3283 vssi a_3 mbk_sig1976 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3284 vssi mbk_sig1976 heart_a_3 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3285 heart_a_3 mbk_sig1976 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3286 a_2 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3287 vsse vsse a_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3288 a_2 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3289 vsse vsse a_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3290 vssi a_2 mbk_sig1977 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3291 mbk_sig1977 a_2 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3292 vssi a_2 mbk_sig1977 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3293 vssi mbk_sig1977 heart_a_2 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3294 heart_a_2 mbk_sig1977 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3295 a_1 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3296 vsse vsse a_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3297 a_1 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3298 vsse vsse a_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3299 vssi a_1 mbk_sig1978 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3300 mbk_sig1978 a_1 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3301 vssi a_1 mbk_sig1978 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3302 vssi mbk_sig1978 heart_a_1 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3303 heart_a_1 mbk_sig1978 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3304 a_0 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3305 vsse vsse a_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3306 a_0 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3307 vsse vsse a_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3308 vssi a_0 mbk_sig1979 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3309 mbk_sig1979 a_0 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3310 vssi a_0 mbk_sig1979 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3311 vssi mbk_sig1979 heart_a_0 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3312 heart_a_0 mbk_sig1979 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3313 b_3 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3314 vsse vsse b_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3315 b_3 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3316 vsse vsse b_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3317 vssi b_3 mbk_sig1980 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3318 mbk_sig1980 b_3 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3319 vssi b_3 mbk_sig1980 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3320 vssi mbk_sig1980 heart_b_3 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3321 heart_b_3 mbk_sig1980 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3322 b_2 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3323 vsse vsse b_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3324 b_2 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3325 vsse vsse b_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3326 vssi b_2 mbk_sig1981 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3327 mbk_sig1981 b_2 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3328 vssi b_2 mbk_sig1981 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3329 vssi mbk_sig1981 heart_b_2 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3330 heart_b_2 mbk_sig1981 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3331 b_1 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3332 vsse vsse b_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3333 b_1 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3334 vsse vsse b_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3335 vssi b_1 mbk_sig1982 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3336 mbk_sig1982 b_1 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3337 vssi b_1 mbk_sig1982 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3338 vssi mbk_sig1982 heart_b_1 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3339 heart_b_1 mbk_sig1982 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3340 b_0 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3341 vsse vsse b_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3342 b_0 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3343 vsse vsse b_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3344 vssi b_0 mbk_sig1983 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3345 mbk_sig1983 b_0 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3346 vssi b_0 mbk_sig1983 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3347 vssi mbk_sig1983 heart_b_0 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3348 heart_b_0 mbk_sig1983 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3349 d_3 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3350 vsse vsse d_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3351 d_3 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3352 vsse vsse d_3 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3353 vssi d_3 mbk_sig1984 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3354 mbk_sig1984 d_3 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3355 vssi d_3 mbk_sig1984 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3356 vssi mbk_sig1984 heart_d_3 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3357 heart_d_3 mbk_sig1984 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3358 d_2 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3359 vsse vsse d_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3360 d_2 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3361 vsse vsse d_2 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3362 vssi d_2 mbk_sig1985 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3363 mbk_sig1985 d_2 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3364 vssi d_2 mbk_sig1985 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3365 vssi mbk_sig1985 heart_d_2 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3366 heart_d_2 mbk_sig1985 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3367 d_1 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3368 vsse vsse d_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3369 d_1 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3370 vsse vsse d_1 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3371 vssi d_1 mbk_sig1986 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3372 mbk_sig1986 d_1 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3373 vssi d_1 mbk_sig1986 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3374 vssi mbk_sig1986 heart_d_1 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3375 heart_d_1 mbk_sig1986 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3376 d_0 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3377 vsse vsse d_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3378 d_0 vsse vsse vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3379 vsse vsse d_0 vsse TN L=0.18U W=6.3U AS=2.268P AD=2.268P PS=13.32U 
+ PD=13.32U 
M3380 vssi d_0 mbk_sig1987 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3381 mbk_sig1987 d_0 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3382 vssi d_0 mbk_sig1987 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3383 vssi mbk_sig1987 heart_d_0 vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3384 heart_d_0 mbk_sig1987 vssi vsse TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
M3385 heart_block3_no31 heart_block3_pb1 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3386 vssi heart_block3_n3 heart_block3_no31 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3387 mbk_sig1967 heart_block3_no21 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3388 vssi heart_block3_no31 mbk_sig1967 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3389 mbk_sig1969 heart_block3_no31 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3390 heart_block3_x21 heart_block3_no21 mbk_sig1969 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3391 vssi mbk_sig1967 heart_block3_x21 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3392 heart_block3_no21 heart_block3_gb1 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3393 vssi heart_block3_n2 heart_block3_no21 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3394 mbk_sig1965 heart_block4_a29s vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3395 vssi heart_block4_a213s mbk_sig1965 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3396 vssi mbk_sig1965 heart_block4_insh1 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3397 mbk_sig1961 heart_block3_x21 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3398 vssi heart_block3_no41 mbk_sig1961 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3399 mbk_sig1963 heart_block3_no41 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3400 heart_block3_fb1 heart_block3_x21 mbk_sig1963 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3401 vssi mbk_sig1961 heart_block3_fb1 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3402 mbk_sig1960 heart_block3_fb1 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3403 heart_block3_na0_csb heart_block3_fb0 mbk_sig1960 vsse TN L=0.18U 
+ W=2.16U AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3404 vssi heart_block4_decalga mbk_sig1959 vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3405 vssi mbk_sig1959 decalgc vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3406 decalgc mbk_sig1959 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3407 vssi mbk_sig1958 heart_block4_a221s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3408 mbk_sig1958 heart_block4_insh1 mbk_sig1956 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3409 mbk_sig1956 heart_block4_decalga vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3410 vssi mbk_sig1955 heart_block4_a29s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3411 mbk_sig1955 heart_block2_a26ms_i0 mbk_sig1957 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3412 mbk_sig1957 heart_block4_selalu vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3413 vssi heart_block3_fb1 heart_block2_a26ms_i0 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3414 vssi mbk_sig1953 heart_block4_a28s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3415 mbk_sig1953 heart_block2_a27ms_i0 mbk_sig1954 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3416 mbk_sig1954 heart_block4_selalu vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3417 vssi mbk_sig1952 heart_block4_a212s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3418 mbk_sig1952 heart_q_2 mbk_sig1951 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3419 mbk_sig1951 ii_8 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M3420 vssi mbk_sig1949 heart_block4_a219s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3421 mbk_sig1949 heart_block4_insh3 mbk_sig1950 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3422 mbk_sig1950 heart_block4_decalda vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3423 vssi mbk_sig1946 heart_block4_shacc2 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3424 mbk_sig1946 heart_block4_a221s vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3425 vssi heart_block4_a220s mbk_sig1946 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3426 mbk_sig1946 heart_block4_a219s vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3427 vssi mbk_sig1945 heart_block4_a220s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3428 mbk_sig1945 heart_block4_insh2 mbk_sig1943 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3429 mbk_sig1943 heart_block4_decaln vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3430 mbk_sig1942 heart_block4_a28s vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3431 vssi heart_block4_a212s mbk_sig1942 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3432 vssi mbk_sig1942 heart_block4_insh2 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3433 vssi mbk_sig1940 heart_block4_a223s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3434 mbk_sig1940 heart_block4_insh1 mbk_sig1941 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3435 mbk_sig1941 heart_block4_decaln vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3436 vssi mbk_sig1939 heart_block4_a227s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3437 mbk_sig1939 q0i mbk_sig1938 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3438 mbk_sig1938 heart_block4_decalga vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3439 vssi ii_8 heart_block4_decaln vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3440 vssi mbk_sig1936 heart_block4_a217s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3441 mbk_sig1936 heart_block4_insh3 mbk_sig1937 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3442 mbk_sig1937 heart_block4_decaln vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3443 vssi mbk_sig1935 f3c vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M3444 mbk_sig1935 heart_block4_decalga mbk_sig1934 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3445 mbk_sig1934 heart_block4_insh3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3446 vssi mbk_sig1933 heart_block4_a225s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3447 mbk_sig1933 heart_block4_insh1 mbk_sig1932 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3448 mbk_sig1932 heart_block4_decalda vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3449 vssi mbk_sig1925 heart_block5_m_1_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3450 mbk_sig1929 mbk_sig1925 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3451 heart_block5_m_1_2_dff_s mbk_sig1930 mbk_sig1929 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3452 vssi mbk_sig1931 heart_block5_m_1_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3453 vssi heart_block5_m_1_2_dff_m mbk_sig1925 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3454 heart_block5_m_1_2_dff_m heart_block5_ck1 mbk_sig1927 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3455 mbk_sig1930 heart_block5_ck1 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3456 vssi heart_block5_m_1_2_dff_s mbk_sig1931 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3457 heart_block5_s21 heart_block5_m_1_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3458 mbk_sig1927 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3459 vssi heart_b_1 heart_block5_nb1 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3460 vssi mbk_sig1922 heart_block4_shacc0 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3461 mbk_sig1922 heart_block4_a227s vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3462 vssi heart_block4_a226s mbk_sig1922 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3463 mbk_sig1922 heart_block4_a225s vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3464 vssi mbk_sig1921 heart_block4_a224s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3465 mbk_sig1921 heart_block4_insh0 mbk_sig1920 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3466 mbk_sig1920 heart_block4_decalga vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3467 vssi mbk_sig1919 heart_block5_b16 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3468 mbk_sig1919 heart_b_1 mbk_sig1917 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3469 mbk_sig1917 heart_b_2 mbk_sig1918 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3470 mbk_sig1918 heart_b_3 mbk_sig1916 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3471 mbk_sig1916 heart_b_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3472 vssi mbk_sig1914 heart_block5_b14 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3473 mbk_sig1914 heart_block5_nb1 mbk_sig1912 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3474 mbk_sig1912 heart_b_2 mbk_sig1913 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3475 mbk_sig1913 heart_b_3 mbk_sig1915 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3476 mbk_sig1915 heart_b_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3477 vssi mbk_sig1911 heart_block4_a226s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3478 mbk_sig1911 heart_block4_insh0 mbk_sig1910 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3479 mbk_sig1910 heart_block4_decaln vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3480 vssi mbk_sig1909 heart_block5_b8 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3481 mbk_sig1909 heart_b_1 mbk_sig1908 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3482 mbk_sig1908 heart_b_2 mbk_sig1906 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3483 mbk_sig1906 heart_block5_nb3 mbk_sig1907 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3484 mbk_sig1907 heart_b_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3485 vssi mbk_sig1905 heart_block5_b15 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3486 mbk_sig1905 heart_b_1 mbk_sig1903 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3487 mbk_sig1903 heart_b_2 mbk_sig1904 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3488 mbk_sig1904 heart_b_3 mbk_sig1902 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3489 mbk_sig1902 heart_block5_nb0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3490 vssi mbk_sig1900 heart_block5_b13 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3491 mbk_sig1900 heart_block5_nb1 mbk_sig1898 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3492 mbk_sig1898 heart_b_2 mbk_sig1899 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3493 mbk_sig1899 heart_b_3 mbk_sig1901 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3494 mbk_sig1901 heart_block5_nb0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3495 vssi mbk_sig1894 heart_block5_b5 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3496 mbk_sig1894 heart_block5_nb1 mbk_sig1895 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3497 mbk_sig1895 heart_b_2 mbk_sig1896 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3498 mbk_sig1896 heart_block5_nb3 mbk_sig1897 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3499 mbk_sig1897 heart_block5_nb0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3500 vssi mbk_sig1890 heart_block5_b1 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3501 mbk_sig1890 heart_block5_nb1 mbk_sig1892 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3502 mbk_sig1892 heart_block5_nb2 mbk_sig1891 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3503 mbk_sig1891 heart_block5_nb3 mbk_sig1893 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3504 mbk_sig1893 heart_block5_nb0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3505 mbk_sig1889 heart_block5_s18 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3506 heart_block5_b18s heart_block5_b8 mbk_sig1889 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3507 vssi mbk_sig1883 heart_block5_m_8_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3508 mbk_sig1887 mbk_sig1883 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3509 heart_block5_m_8_1_dff_s mbk_sig1885 mbk_sig1887 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3510 vssi mbk_sig1888 heart_block5_m_8_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3511 vssi heart_block5_m_8_1_dff_m mbk_sig1883 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3512 heart_block5_m_8_1_dff_m heart_block5_ck8 mbk_sig1881 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3513 mbk_sig1885 heart_block5_ck8 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3514 vssi heart_block5_m_8_1_dff_s mbk_sig1888 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3515 heart_block5_s18 heart_block5_m_8_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3516 mbk_sig1881 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3517 mbk_sig1882 heart_block5_s18 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3518 heart_block5_a18s heart_block5_a8 mbk_sig1882 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3519 vssi mbk_sig1880 heart_block5_b10 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3520 mbk_sig1880 heart_block5_nb1 mbk_sig1878 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3521 mbk_sig1878 heart_block5_nb2 mbk_sig1879 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3522 mbk_sig1879 heart_b_3 mbk_sig1877 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3523 mbk_sig1877 heart_b_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3524 vssi mbk_sig1876 heart_block5_ck5 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3525 mbk_sig1876 heart_block5_enable mbk_sig1875 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3526 mbk_sig1875 heart_block5_b5 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3527 vssi mbk_sig1874 heart_block5_ck8 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3528 mbk_sig1874 heart_block5_enable mbk_sig1873 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3529 mbk_sig1873 heart_block5_b8 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3530 vssi mbk_sig1866 heart_block5_m_8_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3531 mbk_sig1870 mbk_sig1866 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3532 heart_block5_m_8_2_dff_s mbk_sig1872 mbk_sig1870 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3533 vssi mbk_sig1871 heart_block5_m_8_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3534 vssi heart_block5_m_8_2_dff_m mbk_sig1866 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3535 heart_block5_m_8_2_dff_m heart_block5_ck8 mbk_sig1868 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3536 mbk_sig1872 heart_block5_ck8 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3537 vssi heart_block5_m_8_2_dff_s mbk_sig1871 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3538 heart_block5_s28 heart_block5_m_8_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3539 mbk_sig1868 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3540 mbk_sig1864 heart_block5_s38 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3541 heart_block5_b38s heart_block5_b8 mbk_sig1864 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3542 vssi mbk_sig1857 heart_block5_m_5_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3543 mbk_sig1862 mbk_sig1857 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3544 heart_block5_m_5_1_dff_s mbk_sig1863 mbk_sig1862 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3545 vssi mbk_sig1865 heart_block5_m_5_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3546 vssi heart_block5_m_5_1_dff_m mbk_sig1857 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3547 heart_block5_m_5_1_dff_m heart_block5_ck5 mbk_sig1860 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3548 mbk_sig1863 heart_block5_ck5 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3549 vssi heart_block5_m_5_1_dff_s mbk_sig1865 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3550 heart_block5_s15 heart_block5_m_5_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3551 mbk_sig1860 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3552 mbk_sig1859 heart_block5_s04 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3553 heart_block5_b04s heart_block5_b4 mbk_sig1859 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3554 vssi mbk_sig1854 heart_block5_m_4_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3555 mbk_sig1852 mbk_sig1854 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3556 heart_block5_m_4_0_dff_s mbk_sig1853 mbk_sig1852 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3557 vssi mbk_sig1856 heart_block5_m_4_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3558 vssi heart_block5_m_4_0_dff_m mbk_sig1854 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3559 heart_block5_m_4_0_dff_m heart_block5_ck4 mbk_sig1851 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3560 mbk_sig1853 heart_block5_ck4 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3561 vssi heart_block5_m_4_0_dff_s mbk_sig1856 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3562 heart_block5_s04 heart_block5_m_4_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3563 mbk_sig1851 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3564 vssi heart_b_0 heart_block5_nb0 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3565 vssi mbk_sig1844 heart_block5_m_8_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3566 mbk_sig1848 mbk_sig1844 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3567 heart_block5_m_8_3_dff_s mbk_sig1846 mbk_sig1848 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3568 vssi mbk_sig1849 heart_block5_m_8_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3569 vssi heart_block5_m_8_3_dff_m mbk_sig1844 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3570 heart_block5_m_8_3_dff_m heart_block5_ck8 mbk_sig1843 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3571 mbk_sig1846 heart_block5_ck8 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3572 vssi heart_block5_m_8_3_dff_s mbk_sig1849 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3573 heart_block5_s38 heart_block5_m_8_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3574 mbk_sig1843 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3575 mbk_sig1842 heart_block5_s33 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3576 heart_block5_a33s heart_block5_a3 mbk_sig1842 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3577 vssi mbk_sig1841 heart_block5_ck2 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3578 mbk_sig1841 heart_block5_enable mbk_sig1839 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3579 mbk_sig1839 heart_block5_b2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3580 vssi mbk_sig1838 heart_block5_ck3 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3581 mbk_sig1838 heart_block5_enable mbk_sig1840 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3582 mbk_sig1840 heart_block5_b3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3583 mbk_sig1837 heart_block5_s33 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3584 heart_block5_b33s heart_block5_b3 mbk_sig1837 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3585 vssi heart_block3_pb1 heart_block3_not1 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3586 mbk_sig1788 heart_block3_cout0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3587 heart_block3_na21 heart_block3_not1 mbk_sig1788 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3588 mbk_sig1787 heart_block3_ni5 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3589 mbk_sig1786 ii_4 mbk_sig1787 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3590 heart_block3_nn3 ii_3 mbk_sig1786 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3591 mbk_sig1784 heart_block3_na20 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3592 heart_block3_cout0 heart_block3_gb0 mbk_sig1784 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3593 heart_block3_no41 heart_block3_cout0 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3594 vssi heart_block3_n4 heart_block3_no41 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3595 heart_block3_n2 heart_block3_ni5 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3596 vssi ii_4 heart_block3_n2 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M3597 mbk_sig1783 ii_3 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3598 heart_block3_flag1 ii_4 mbk_sig1783 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3599 mbk_sig1782 heart_block3_nn3 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3600 heart_block3_n4 heart_block3_ni5 mbk_sig1782 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3601 mbk_sig1781 heart_block3_na21 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3602 heart_block3_cout1 heart_block3_gb1 mbk_sig1781 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3603 vssi mbk_sig1779 heart_block4_a213s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3604 mbk_sig1779 heart_q_1 mbk_sig1809 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3605 mbk_sig1809 ii_8 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M3606 mbk_sig1777 heart_block3_signea vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3607 heart_block3_na1_csb heart_block3_fb2 mbk_sig1777 vsse TN L=0.18U 
+ W=2.16U AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3608 zeroc heart_block3_na1_csb vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3609 vssi heart_block3_na0_csb zeroc vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3610 mbk_sig1805 heart_block3_x22 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3611 vssi heart_block3_no42 mbk_sig1805 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3612 mbk_sig1775 heart_block3_no42 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3613 heart_block3_fb2 heart_block3_x22 mbk_sig1775 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3614 vssi mbk_sig1805 heart_block3_fb2 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3615 vssi mbk_sig1774 heart_block5_a26sh vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3616 mbk_sig1774 heart_block2_a26ms_i0 mbk_sig1804 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3617 mbk_sig1804 heart_block5_decalgra vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3618 heart_block3_no42 heart_block3_cout1 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3619 vssi heart_block3_n4 heart_block3_no42 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3620 vssi mbk_sig1773 heart_block3_flag vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3621 mbk_sig1773 heart_block3_ni5 mbk_sig1802 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3622 mbk_sig1802 heart_block3_flag1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3623 mbk_sig1763 mbk_sig1765 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3624 mbk_sig1764 heart_block4_shacc1 mbk_sig1763 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3625 vssi heart_block4_test_mode mbk_sig1765 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3626 vssi mbk_sig1772 heart_block4_m1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3627 heart_block4_m1_dff_s mbk_sig1768 mbk_sig1770 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3628 mbk_sig1766 heart_q_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3629 mbk_sig1764 heart_block4_test_mode mbk_sig1766 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3630 heart_q_1 heart_block4_m1_dff_s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3631 vssi heart_block4_m1_dff_s mbk_sig1772 vsse TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M3632 mbk_sig1770 mbk_sig1769 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3633 vssi mbk_sig1769 heart_block4_m1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3634 heart_block4_m1_dff_m heart_block4_ckin mbk_sig1764 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3635 vssi heart_block4_m1_dff_m mbk_sig1769 vsse TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M3636 mbk_sig1768 heart_block4_ckin vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3637 vssi mbk_sig1762 heart_block4_shacc1 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3638 mbk_sig1762 heart_block4_a224s vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3639 vssi heart_block4_a223s mbk_sig1762 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3640 mbk_sig1762 heart_block4_a222s vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3641 vssi mbk_sig1757 heart_block4_a222s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3642 mbk_sig1757 heart_block4_insh2 mbk_sig1798 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3643 mbk_sig1798 heart_block4_decalda vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3644 vssi mbk_sig1756 heart_block5_shram2 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3645 mbk_sig1756 heart_block5_a28sh vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3646 vssi heart_block5_a27sh mbk_sig1756 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3647 mbk_sig1756 heart_block5_a26sh vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3648 vssi mbk_sig1754 heart_block4_a27s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3649 mbk_sig1754 heart_block2_a28ms_i0 mbk_sig1794 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3650 mbk_sig1794 heart_block4_selalu vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3651 mbk_sig1752 heart_block4_a27s vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3652 vssi heart_block4_a211s mbk_sig1752 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M3653 vssi mbk_sig1752 heart_block4_insh3 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3654 vssi heart_b_3 heart_block5_nb3 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3655 vssi mbk_sig1751 heart_block4_decalda vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3656 mbk_sig1751 ii_8 mbk_sig1793 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3657 mbk_sig1793 heart_block4_ni7 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3658 vssi mbk_sig1746 heart_block5_m_1_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3659 mbk_sig1748 mbk_sig1746 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3660 heart_block5_m_1_1_dff_s mbk_sig1749 mbk_sig1748 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3661 vssi mbk_sig1750 heart_block5_m_1_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3662 vssi heart_block5_m_1_1_dff_m mbk_sig1746 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3663 heart_block5_m_1_1_dff_m heart_block5_ck1 mbk_sig1745 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3664 mbk_sig1749 heart_block5_ck1 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3665 vssi heart_block5_m_1_1_dff_s mbk_sig1750 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3666 heart_block5_s11 heart_block5_m_1_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3667 mbk_sig1745 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3668 vssi heart_b_2 heart_block5_nb2 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3669 vssi mbk_sig1743 f0c vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M3670 mbk_sig1743 heart_block4_decalda mbk_sig1792 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3671 mbk_sig1792 heart_block4_insh0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3672 vssi mbk_sig1739 heart_block5_b6 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3673 mbk_sig1739 heart_block5_nb1 mbk_sig1740 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3674 mbk_sig1740 heart_b_2 mbk_sig1741 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3675 mbk_sig1741 heart_block5_nb3 mbk_sig1742 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3676 mbk_sig1742 heart_b_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3677 mbk_sig1738 heart_block5_s27 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3678 heart_block5_b27s heart_block5_b7 mbk_sig1738 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3679 vssi mbk_sig1735 heart_block5_b7 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3680 mbk_sig1735 heart_b_1 mbk_sig1736 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3681 mbk_sig1736 heart_b_2 mbk_sig1732 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3682 mbk_sig1732 heart_block5_nb3 mbk_sig1733 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3683 mbk_sig1733 heart_block5_nb0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3684 mbk_sig1734 heart_block5_s11 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3685 heart_block5_b11s heart_block5_b1 mbk_sig1734 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3686 vssi mbk_sig1728 heart_block5_b4 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3687 mbk_sig1728 heart_b_1 mbk_sig1730 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3688 mbk_sig1730 heart_block5_nb2 mbk_sig1729 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3689 mbk_sig1729 heart_block5_nb3 mbk_sig1731 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3690 mbk_sig1731 heart_b_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3691 vssi mbk_sig1724 heart_block5_ob431s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3692 mbk_sig1724 heart_block5_b16s mbk_sig1726 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3693 mbk_sig1726 heart_block5_b17s mbk_sig1727 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3694 mbk_sig1727 heart_block5_b18s mbk_sig1723 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3695 mbk_sig1723 heart_block5_b15s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3696 vssi mbk_sig1721 heart_block5_b2 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3697 mbk_sig1721 heart_block5_nb1 mbk_sig1722 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3698 mbk_sig1722 heart_block5_nb2 mbk_sig1720 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3699 mbk_sig1720 heart_block5_nb3 mbk_sig1719 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3700 mbk_sig1719 heart_b_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3701 vssi mbk_sig1714 heart_block5_m_1_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3702 mbk_sig1716 mbk_sig1714 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3703 heart_block5_m_1_0_dff_s mbk_sig1717 mbk_sig1716 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3704 vssi mbk_sig1718 heart_block5_m_1_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3705 vssi heart_block5_m_1_0_dff_m mbk_sig1714 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3706 heart_block5_m_1_0_dff_m heart_block5_ck1 mbk_sig1713 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3707 mbk_sig1717 heart_block5_ck1 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3708 vssi heart_block5_m_1_0_dff_s mbk_sig1718 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3709 heart_block5_s01 heart_block5_m_1_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3710 mbk_sig1713 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3711 mbk_sig1709 heart_block5_s25 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3712 heart_block5_b25s heart_block5_b5 mbk_sig1709 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3713 mbk_sig1711 heart_block5_s17 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3714 heart_block5_b17s heart_block5_b7 mbk_sig1711 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3715 vssi mbk_sig1704 heart_block5_b12 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3716 mbk_sig1704 heart_b_1 mbk_sig1706 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3717 mbk_sig1706 heart_block5_nb2 mbk_sig1705 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3718 mbk_sig1705 heart_b_3 mbk_sig1707 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3719 mbk_sig1707 heart_b_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3720 mbk_sig1703 heart_block5_s24 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3721 heart_block5_b24s heart_block5_b4 mbk_sig1703 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3722 mbk_sig1702 heart_block5_s17 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3723 heart_block5_a17s heart_block5_a7 mbk_sig1702 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3724 vssi mbk_sig1698 heart_block5_b3 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3725 mbk_sig1698 heart_b_1 mbk_sig1700 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3726 mbk_sig1700 heart_block5_nb2 mbk_sig1701 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3727 mbk_sig1701 heart_block5_nb3 mbk_sig1697 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3728 mbk_sig1697 heart_block5_nb0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3729 vssi mbk_sig1692 heart_block5_m_5_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3730 mbk_sig1694 mbk_sig1692 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3731 heart_block5_m_5_2_dff_s mbk_sig1695 mbk_sig1694 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3732 vssi mbk_sig1696 heart_block5_m_5_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3733 vssi heart_block5_m_5_2_dff_m mbk_sig1692 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3734 heart_block5_m_5_2_dff_m heart_block5_ck5 mbk_sig1691 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3735 mbk_sig1695 heart_block5_ck5 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3736 vssi heart_block5_m_5_2_dff_s mbk_sig1696 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3737 heart_block5_s25 heart_block5_m_5_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3738 mbk_sig1691 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3739 mbk_sig1688 heart_block5_s28 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3740 heart_block5_a28s heart_block5_a8 mbk_sig1688 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3741 mbk_sig1687 heart_block5_s38 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3742 heart_block5_a38s heart_block5_a8 mbk_sig1687 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3743 vssi mbk_sig1683 heart_block5_m_4_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3744 mbk_sig1685 mbk_sig1683 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3745 heart_block5_m_4_2_dff_s mbk_sig1680 mbk_sig1685 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3746 vssi mbk_sig1686 heart_block5_m_4_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3747 vssi heart_block5_m_4_2_dff_m mbk_sig1683 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3748 heart_block5_m_4_2_dff_m heart_block5_ck4 mbk_sig1682 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3749 mbk_sig1680 heart_block5_ck4 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3750 vssi heart_block5_m_4_2_dff_s mbk_sig1686 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3751 heart_block5_s24 heart_block5_m_4_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3752 mbk_sig1682 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3753 vssi mbk_sig1679 heart_block5_ck1 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3754 mbk_sig1679 heart_block5_enable mbk_sig1791 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3755 mbk_sig1791 heart_block5_b1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3756 mbk_sig1676 heart_block5_s04 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3757 heart_block5_a04s heart_block5_a4 mbk_sig1676 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3758 mbk_sig1677 heart_block5_s31 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3759 heart_block5_b31s heart_block5_b1 mbk_sig1677 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3760 vssi mbk_sig1673 heart_block5_m_1_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3761 mbk_sig1671 mbk_sig1673 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3762 heart_block5_m_1_3_dff_s mbk_sig1672 mbk_sig1671 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3763 vssi mbk_sig1675 heart_block5_m_1_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3764 vssi heart_block5_m_1_3_dff_m mbk_sig1673 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3765 heart_block5_m_1_3_dff_m heart_block5_ck1 mbk_sig1666 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3766 mbk_sig1672 heart_block5_ck1 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3767 vssi heart_block5_m_1_3_dff_s mbk_sig1675 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3768 heart_block5_s31 heart_block5_m_1_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3769 mbk_sig1666 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3770 vssi mbk_sig1664 heart_block5_ob443s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3771 mbk_sig1664 heart_block5_b32s mbk_sig1667 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3772 mbk_sig1667 heart_block5_b33s mbk_sig1665 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3773 mbk_sig1665 heart_block5_b34s mbk_sig1661 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3774 mbk_sig1661 heart_block5_b31s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3775 vssi mbk_sig1656 heart_block5_m_3_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3776 mbk_sig1658 mbk_sig1656 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3777 heart_block5_m_3_3_dff_s mbk_sig1659 mbk_sig1658 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3778 vssi mbk_sig1660 heart_block5_m_3_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3779 vssi heart_block5_m_3_3_dff_m mbk_sig1656 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3780 heart_block5_m_3_3_dff_m heart_block5_ck3 mbk_sig1655 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3781 mbk_sig1659 heart_block5_ck3 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3782 vssi heart_block5_m_3_3_dff_s mbk_sig1660 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3783 heart_block5_s33 heart_block5_m_3_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3784 mbk_sig1655 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3785 vssi heart_block3_nn3 heart_block3_n3 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3786 mbk_sig1626 heart_block3_x23 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3787 vssi heart_block3_no43 mbk_sig1626 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3788 mbk_sig1628 heart_block3_no43 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3789 heart_block3_signea heart_block3_x23 mbk_sig1628 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3790 vssi mbk_sig1626 heart_block3_signea vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3791 mbk_sig1623 heart_block3_no23 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3792 vssi heart_block3_no33 mbk_sig1623 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3793 mbk_sig1622 heart_block3_no33 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3794 heart_block3_x23 heart_block3_no23 mbk_sig1622 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3795 vssi mbk_sig1623 heart_block3_x23 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3796 mbk_sig1621 cini vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3797 heart_block3_na20 heart_block3_not0 mbk_sig1621 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3798 heart_block3_no23 heart_block3_gb3 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3799 vssi heart_block3_n2 heart_block3_no23 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3800 heart_block3_no40 cini vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3801 vssi heart_block3_n4 heart_block3_no40 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3802 mbk_sig1614 heart_block3_x20 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3803 vssi heart_block3_no40 mbk_sig1614 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3804 mbk_sig1616 heart_block3_no40 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3805 heart_block3_fb0 heart_block3_x20 mbk_sig1616 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3806 vssi mbk_sig1614 heart_block3_fb0 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3807 vssi heart_block3_signea heart_block2_a28ms_i0 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3808 vssi heart_block3_signea signec vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3809 mbk_sig1601 mbk_sig1602 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3810 mbk_sig1603 heart_block4_shacc2 mbk_sig1601 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3811 vssi heart_block4_test_mode mbk_sig1602 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3812 vssi mbk_sig1612 heart_block4_m2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3813 heart_block4_m2_dff_s mbk_sig1608 mbk_sig1610 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3814 mbk_sig1604 heart_q_1 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3815 mbk_sig1603 heart_block4_test_mode mbk_sig1604 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3816 heart_q_2 heart_block4_m2_dff_s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3817 vssi heart_block4_m2_dff_s mbk_sig1612 vsse TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M3818 mbk_sig1610 mbk_sig1609 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3819 vssi mbk_sig1609 heart_block4_m2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3820 heart_block4_m2_dff_m heart_block4_ckin mbk_sig1603 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3821 vssi heart_block4_m2_dff_m mbk_sig1609 vsse TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M3822 mbk_sig1608 heart_block4_ckin vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3823 vssi mbk_sig1597 heart_block5_a27sh vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3824 mbk_sig1597 heart_block2_a27ms_i0 mbk_sig1600 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3825 mbk_sig1600 heart_block5_decalnr vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3826 vssi heart_block3_fb0 heart_block2_a25ms_i0 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3827 vssi heart_block3_fb2 heart_block2_a27ms_i0 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3828 vssi mbk_sig1590 heart_block5_m_3_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3829 mbk_sig1594 mbk_sig1590 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3830 heart_block5_m_3_2_dff_s mbk_sig1592 mbk_sig1594 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3831 vssi mbk_sig1595 heart_block5_m_3_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3832 vssi heart_block5_m_3_2_dff_m mbk_sig1590 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3833 heart_block5_m_3_2_dff_m heart_block5_ck3 mbk_sig1587 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3834 mbk_sig1592 heart_block5_ck3 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3835 vssi heart_block5_m_3_2_dff_s mbk_sig1595 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3836 heart_block5_s23 heart_block5_m_3_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3837 mbk_sig1587 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3838 vssi mbk_sig1588 heart_block4_a210s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3839 mbk_sig1588 heart_block2_a25ms_i0 mbk_sig1589 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3840 mbk_sig1589 heart_block4_selalu vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3841 vssi mbk_sig1586 s3c vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M3842 mbk_sig1586 heart_block5_decalgra mbk_sig1585 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3843 mbk_sig1585 heart_block2_a28ms_i0 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3844 vssi mbk_sig1584 heart_block5_a28sh vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3845 mbk_sig1584 heart_block2_a28ms_i0 mbk_sig1583 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3846 mbk_sig1583 heart_block5_decaldra vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3847 vssi mbk_sig1580 heart_block4_a216s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3848 mbk_sig1580 q3i mbk_sig1582 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3849 mbk_sig1582 heart_block4_decalda vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3850 vssi mbk_sig1573 heart_block5_m_6_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3851 mbk_sig1577 mbk_sig1573 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3852 heart_block5_m_6_3_dff_s mbk_sig1578 mbk_sig1577 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3853 vssi mbk_sig1579 heart_block5_m_6_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3854 vssi heart_block5_m_6_3_dff_m mbk_sig1573 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3855 heart_block5_m_6_3_dff_m heart_block5_ck6 mbk_sig1575 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3856 mbk_sig1578 heart_block5_ck6 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3857 vssi heart_block5_m_6_3_dff_s mbk_sig1579 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3858 heart_block5_s36 heart_block5_m_6_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3859 mbk_sig1575 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3860 vssi mbk_sig1572 heart_block4_a211s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3861 mbk_sig1572 heart_q_3 mbk_sig1570 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3862 mbk_sig1570 ii_8 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M3863 vssi heart_block4_decalda mbk_sig1567 vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3864 vssi mbk_sig1567 decaldc vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3865 decaldc mbk_sig1567 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3866 mbk_sig1568 heart_block5_s21 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3867 heart_block5_b21s heart_block5_b1 mbk_sig1568 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3868 mbk_sig1564 heart_block5_s23 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3869 heart_block5_b23s heart_block5_b3 mbk_sig1564 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3870 mbk_sig1565 heart_block5_s21 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3871 heart_block5_a21s heart_block5_a1 mbk_sig1565 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3872 mbk_sig1563 heart_block5_s26 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3873 heart_block5_b26s heart_block5_b6 mbk_sig1563 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3874 vssi mbk_sig1558 heart_block5_ob432s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3875 mbk_sig1558 heart_block5_b26s mbk_sig1560 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3876 mbk_sig1560 heart_block5_b27s mbk_sig1561 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3877 mbk_sig1561 heart_block5_b28s mbk_sig1556 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3878 mbk_sig1556 heart_block5_b25s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3879 vssi mbk_sig1554 heart_block5_ck7 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3880 mbk_sig1554 heart_block5_enable mbk_sig1557 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3881 mbk_sig1557 heart_block5_b7 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3882 vssi mbk_sig1549 heart_block5_ob442s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3883 mbk_sig1549 heart_block5_b22s mbk_sig1551 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3884 mbk_sig1551 heart_block5_b23s mbk_sig1552 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3885 mbk_sig1552 heart_block5_b24s mbk_sig1553 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3886 mbk_sig1553 heart_block5_b21s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3887 vssi mbk_sig1546 heart_block5_b11 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3888 mbk_sig1546 heart_b_1 mbk_sig1547 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3889 mbk_sig1547 heart_block5_nb2 mbk_sig1548 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3890 mbk_sig1548 heart_b_3 mbk_sig1545 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3891 mbk_sig1545 heart_block5_nb0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3892 mbk_sig1543 heart_block5_s15 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3893 heart_block5_b15s heart_block5_b5 mbk_sig1543 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3894 vssi mbk_sig1536 heart_block5_m_7_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3895 mbk_sig1540 mbk_sig1536 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3896 heart_block5_m_7_1_dff_s mbk_sig1538 mbk_sig1540 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3897 vssi mbk_sig1542 heart_block5_m_7_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3898 vssi heart_block5_m_7_1_dff_m mbk_sig1536 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3899 heart_block5_m_7_1_dff_m heart_block5_ck7 mbk_sig1534 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3900 mbk_sig1538 heart_block5_ck7 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3901 vssi heart_block5_m_7_1_dff_s mbk_sig1542 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3902 heart_block5_s17 heart_block5_m_7_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3903 mbk_sig1534 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3904 vssi mbk_sig1526 heart_block5_m_8_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3905 mbk_sig1532 mbk_sig1526 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3906 heart_block5_m_8_0_dff_s mbk_sig1533 mbk_sig1532 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3907 vssi mbk_sig1535 heart_block5_m_8_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3908 vssi heart_block5_m_8_0_dff_m mbk_sig1526 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3909 heart_block5_m_8_0_dff_m heart_block5_ck8 mbk_sig1529 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3910 mbk_sig1533 heart_block5_ck8 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3911 vssi heart_block5_m_8_0_dff_s mbk_sig1535 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3912 heart_block5_s08 heart_block5_m_8_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3913 mbk_sig1529 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3914 mbk_sig1528 heart_block5_s22 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3915 heart_block5_b22s heart_block5_b2 mbk_sig1528 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3916 mbk_sig1524 heart_block5_s15 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3917 heart_block5_a15s heart_block5_a5 mbk_sig1524 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3918 vssi mbk_sig1521 heart_block5_oa431s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3919 mbk_sig1521 heart_block5_a16s mbk_sig1519 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3920 mbk_sig1519 heart_block5_a17s mbk_sig1520 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3921 mbk_sig1520 heart_block5_a18s mbk_sig1518 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3922 mbk_sig1518 heart_block5_a15s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3923 mbk_sig1515 heart_block5_s01 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3924 heart_block5_b01s heart_block5_b1 mbk_sig1515 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3925 vssi mbk_sig1514 heart_block5_ck4 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3926 mbk_sig1514 heart_block5_enable mbk_sig1516 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3927 mbk_sig1516 heart_block5_b4 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3928 mbk_sig1512 heart_block5_s24 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3929 heart_block5_a24s heart_block5_a4 mbk_sig1512 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3930 mbk_sig1508 heart_block5_s28 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3931 heart_block5_b28s heart_block5_b8 mbk_sig1508 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3932 vssi mbk_sig1506 heart_block5_ob441s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3933 mbk_sig1506 heart_block5_b12s mbk_sig1509 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3934 mbk_sig1509 heart_block5_b13s mbk_sig1510 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3935 mbk_sig1510 heart_block5_b14s mbk_sig1504 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3936 mbk_sig1504 heart_block5_b11s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3937 mbk_sig1505 heart_block5_s14 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3938 heart_block5_a14s heart_block5_a4 mbk_sig1505 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3939 mbk_sig1503 heart_block5_s14 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3940 heart_block5_b14s heart_block5_b4 mbk_sig1503 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3941 mbk_sig1500 heart_block5_s31 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3942 heart_block5_a31s heart_block5_a1 mbk_sig1500 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3943 vssi mbk_sig1498 heart_block5_m_4_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3944 mbk_sig1496 mbk_sig1498 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3945 heart_block5_m_4_1_dff_s mbk_sig1497 mbk_sig1496 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3946 vssi mbk_sig1501 heart_block5_m_4_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3947 vssi heart_block5_m_4_1_dff_m mbk_sig1498 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3948 heart_block5_m_4_1_dff_m heart_block5_ck4 mbk_sig1493 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3949 mbk_sig1497 heart_block5_ck4 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3950 vssi heart_block5_m_4_1_dff_s mbk_sig1501 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3951 heart_block5_s14 heart_block5_m_4_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3952 mbk_sig1493 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3953 vssi mbk_sig1491 heart_block5_oa443s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3954 mbk_sig1491 heart_block5_a32s mbk_sig1495 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3955 mbk_sig1495 heart_block5_a33s mbk_sig1490 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3956 mbk_sig1490 heart_block5_a34s mbk_sig1489 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3957 mbk_sig1489 heart_block5_a31s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3958 vssi mbk_sig1481 heart_block5_m_4_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3959 mbk_sig1486 mbk_sig1481 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3960 heart_block5_m_4_3_dff_s mbk_sig1488 mbk_sig1486 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3961 vssi mbk_sig1487 heart_block5_m_4_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M3962 vssi heart_block5_m_4_3_dff_m mbk_sig1481 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3963 heart_block5_m_4_3_dff_m heart_block5_ck4 mbk_sig1483 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3964 mbk_sig1488 heart_block5_ck4 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M3965 vssi heart_block5_m_4_3_dff_s mbk_sig1487 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M3966 heart_block5_s34 heart_block5_m_4_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3967 mbk_sig1483 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3968 mbk_sig1477 heart_block5_s34 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3969 heart_block5_b34s heart_block5_b4 mbk_sig1477 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3970 mbk_sig1478 heart_block5_s32 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3971 heart_block5_b32s heart_block5_b2 mbk_sig1478 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3972 mbk_sig1475 heart_block5_s32 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3973 heart_block5_a32s heart_block5_a2 mbk_sig1475 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3974 mbk_sig1474 heart_block5_s12 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3975 heart_block5_b12s heart_block5_b2 mbk_sig1474 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3976 mbk_sig1473 heart_block5_s03 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3977 heart_block5_a03s heart_block5_a3 mbk_sig1473 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3978 mbk_sig1446 heart_block3_na22 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3979 heart_block3_cout2 heart_block3_gb2 mbk_sig1446 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3980 mbk_sig1444 heart_block3_cout1 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3981 heart_block3_na22 heart_block3_not2 mbk_sig1444 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3982 heart_block3_no43 heart_block3_cout2 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3983 vssi heart_block3_n4 heart_block3_no43 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3984 heart_block3_no33 heart_block3_pb3 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3985 vssi heart_block3_n3 heart_block3_no33 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3986 vssi ii_5 heart_block3_ni5 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M3987 mbk_sig1436 ii_5 mbk_sig1434 vsse TN L=0.18U W=1.98U AS=0.7128P 
+ AD=0.7128P PS=4.68U PD=4.68U 
M3988 vssi ii_3 mbk_sig1436 vsse TN L=0.18U W=1.98U AS=0.7128P AD=0.7128P 
+ PS=4.68U PD=4.68U 
M3989 vssi ii_5 mbk_sig1435 vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3990 mbk_sig1435 ii_3 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M3991 heart_block3_nn0 mbk_sig1434 mbk_sig1435 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3992 mbk_sig1429 heart_block3_no20 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3993 vssi heart_block3_no30 mbk_sig1429 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3994 mbk_sig1432 heart_block3_no30 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M3995 heart_block3_x20 heart_block3_no20 mbk_sig1432 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M3996 vssi mbk_sig1429 heart_block3_x20 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M3997 vssi heart_block3_g ngc vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M3998 heart_block3_pb1 heart_block3_x11 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M3999 vssi heart_block3_x01 heart_block3_pb1 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4000 mbk_sig1427 heart_block3_x11 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4001 heart_block3_gb1 heart_block3_x01 mbk_sig1427 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4002 mbk_sig1423 heart_block4_decaln vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4003 mbk_sig1422 heart_block4_ni7 mbk_sig1423 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4004 mbk_sig1426 heart_block4_ni6 mbk_sig1422 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4005 vssi mbk_sig1426 heart_block4_selalu vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4006 mbk_sig1415 mbk_sig1413 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4007 mbk_sig1414 heart_block4_shacc3 mbk_sig1415 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4008 vssi heart_block4_test_mode mbk_sig1413 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4009 vssi mbk_sig1421 heart_block4_m3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4010 heart_block4_m3_dff_s mbk_sig1417 mbk_sig1420 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4011 mbk_sig1410 heart_q_2 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M4012 mbk_sig1414 heart_block4_test_mode mbk_sig1410 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4013 heart_q_3 heart_block4_m3_dff_s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4014 vssi heart_block4_m3_dff_s mbk_sig1421 vsse TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M4015 mbk_sig1420 mbk_sig1418 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4016 vssi mbk_sig1418 heart_block4_m3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4017 heart_block4_m3_dff_m heart_block4_ckin mbk_sig1414 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4018 vssi heart_block4_m3_dff_m mbk_sig1418 vsse TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M4019 mbk_sig1417 heart_block4_ckin vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4020 vssi mbk_sig1409 heart_block5_a214sh vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4021 mbk_sig1409 heart_block2_a26ms_i0 mbk_sig1411 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4022 mbk_sig1411 heart_block5_decaldra vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4023 vssi mbk_sig1407 heart_block5_a29sh vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4024 mbk_sig1407 heart_block2_a25ms_i0 mbk_sig1408 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4025 mbk_sig1408 heart_block5_decalgra vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4026 mbk_sig1399 mbk_sig1397 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4027 mbk_sig1398 heart_block4_shacc0 mbk_sig1399 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4028 vssi heart_block4_test_mode mbk_sig1397 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4029 vssi mbk_sig1406 heart_block4_m0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4030 heart_block4_m0_dff_s mbk_sig1402 mbk_sig1404 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4031 mbk_sig1391 scini vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M4032 mbk_sig1398 heart_block4_test_mode mbk_sig1391 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4033 heart_q_0 heart_block4_m0_dff_s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4034 vssi heart_block4_m0_dff_s mbk_sig1406 vsse TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M4035 mbk_sig1404 mbk_sig1403 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4036 vssi mbk_sig1403 heart_block4_m0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4037 heart_block4_m0_dff_m heart_block4_ckin mbk_sig1398 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4038 vssi heart_block4_m0_dff_m mbk_sig1403 vsse TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
M4039 mbk_sig1402 heart_block4_ckin vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4040 vssi mbk_sig1389 heart_block4_shacc3 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4041 mbk_sig1389 heart_block4_a218s vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4042 vssi heart_block4_a217s mbk_sig1389 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4043 mbk_sig1389 heart_block4_a216s vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4044 vssi noei oec vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
M4045 vssi mbk_sig1387 heart_block4_a218s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4046 mbk_sig1387 heart_block4_insh2 mbk_sig1388 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4047 mbk_sig1388 heart_block4_decalga vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4048 vssi mbk_sig1385 heart_block4_a214s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4049 mbk_sig1385 heart_q_0 mbk_sig1386 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4050 mbk_sig1386 ii_8 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4051 vssi mbk_sig1384 scoutc vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4052 mbk_sig1384 heart_block4_test_mode mbk_sig1383 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4053 mbk_sig1383 heart_q_3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4054 mbk_sig1378 heart_block4_a210s vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4055 vssi heart_block4_a214s mbk_sig1378 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4056 vssi mbk_sig1378 heart_block4_insh0 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4057 mbk_sig1380 heart_block5_s16 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4058 heart_block5_b16s heart_block5_b6 mbk_sig1380 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4059 vssi ii_8 heart_block5_decalnr vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4060 mbk_sig1376 heart_block5_s23 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4061 heart_block5_a23s heart_block5_a3 mbk_sig1376 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4062 mbk_sig1374 heart_block5_s36 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4063 heart_block5_a36s heart_block5_a6 mbk_sig1374 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4064 vssi mbk_sig1371 heart_block5_oa442s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4065 mbk_sig1371 heart_block5_a22s mbk_sig1369 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4066 mbk_sig1369 heart_block5_a23s mbk_sig1368 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4067 mbk_sig1368 heart_block5_a24s mbk_sig1370 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4068 mbk_sig1370 heart_block5_a21s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4069 mbk_sig1361 heart_block5_s06 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4070 heart_block5_b06s heart_block5_b6 mbk_sig1361 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4071 vssi mbk_sig1360 heart_block5_b9 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4072 mbk_sig1360 heart_block5_nb1 mbk_sig1362 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4073 mbk_sig1362 heart_block5_nb2 mbk_sig1363 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4074 mbk_sig1363 heart_b_3 mbk_sig1364 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4075 mbk_sig1364 heart_block5_nb0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4076 mbk_sig1358 heart_block5_s07 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4077 heart_block5_b07s heart_block5_b7 mbk_sig1358 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4078 vssi mbk_sig1356 heart_block5_oa430s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4079 mbk_sig1356 heart_block5_a06s mbk_sig1354 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4080 mbk_sig1354 heart_block5_a07s mbk_sig1355 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4081 mbk_sig1355 heart_block5_a08s mbk_sig1357 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4082 mbk_sig1357 heart_block5_a05s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4083 vssi mbk_sig1350 heart_block5_ob430s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4084 mbk_sig1350 heart_block5_b06s mbk_sig1351 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4085 mbk_sig1351 heart_block5_b07s mbk_sig1352 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4086 mbk_sig1352 heart_block5_b08s mbk_sig1353 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4087 mbk_sig1353 heart_block5_b05s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4088 mbk_sig1349 heart_block5_s05 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4089 heart_block5_b05s heart_block5_b5 mbk_sig1349 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4090 vssi mbk_sig1343 heart_block5_m_7_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4091 mbk_sig1347 mbk_sig1343 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4092 heart_block5_m_7_0_dff_s mbk_sig1345 mbk_sig1347 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4093 vssi mbk_sig1348 heart_block5_m_7_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4094 vssi heart_block5_m_7_0_dff_m mbk_sig1343 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4095 heart_block5_m_7_0_dff_m heart_block5_ck7 mbk_sig1342 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4096 mbk_sig1345 heart_block5_ck7 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4097 vssi heart_block5_m_7_0_dff_s mbk_sig1348 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4098 heart_block5_s07 heart_block5_m_7_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4099 mbk_sig1342 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4100 mbk_sig1341 heart_block5_s22 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4101 heart_block5_a22s heart_block5_a2 mbk_sig1341 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4102 mbk_sig1338 heart_block5_s07 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4103 heart_block5_a07s heart_block5_a7 mbk_sig1338 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4104 mbk_sig1339 heart_block5_s11 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4105 heart_block5_a11s heart_block5_a1 mbk_sig1339 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4106 mbk_sig1335 heart_block5_s05 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4107 heart_block5_a05s heart_block5_a5 mbk_sig1335 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4108 vssi mbk_sig1333 heart_block5_oa441s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4109 mbk_sig1333 heart_block5_a12s mbk_sig1336 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4110 mbk_sig1336 heart_block5_a13s mbk_sig1337 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4111 mbk_sig1337 heart_block5_a14s mbk_sig1331 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4112 mbk_sig1331 heart_block5_a11s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4113 mbk_sig1332 heart_block5_s13 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4114 heart_block5_a13s heart_block5_a3 mbk_sig1332 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4115 vssi mbk_sig1325 heart_block5_m_3_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4116 mbk_sig1326 mbk_sig1325 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4117 heart_block5_m_3_1_dff_s mbk_sig1328 mbk_sig1326 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4118 vssi mbk_sig1330 heart_block5_m_3_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4119 vssi heart_block5_m_3_1_dff_m mbk_sig1325 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4120 heart_block5_m_3_1_dff_m heart_block5_ck3 mbk_sig1322 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4121 mbk_sig1328 heart_block5_ck3 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4122 vssi heart_block5_m_3_1_dff_s mbk_sig1330 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4123 heart_block5_s13 heart_block5_m_3_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4124 mbk_sig1322 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4125 mbk_sig1324 heart_block5_s13 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4126 heart_block5_b13s heart_block5_b3 mbk_sig1324 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4127 mbk_sig1319 heart_block5_s01 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4128 heart_block5_a01s heart_block5_a1 mbk_sig1319 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4129 vssi mbk_sig1317 heart_block5_oa433s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4130 mbk_sig1317 heart_block5_a36s mbk_sig1320 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4131 mbk_sig1320 heart_block5_a37s mbk_sig1316 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4132 mbk_sig1316 heart_block5_a38s mbk_sig1315 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4133 mbk_sig1315 heart_block5_a35s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4134 vssi mbk_sig1312 heart_block5_ob440s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4135 mbk_sig1312 heart_block5_b02s mbk_sig1311 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4136 mbk_sig1311 heart_block5_b03s mbk_sig1309 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4137 mbk_sig1309 heart_block5_b04s mbk_sig1310 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4138 mbk_sig1310 heart_block5_b01s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4139 mbk_sig1306 heart_block5_s02 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4140 heart_block5_b02s heart_block5_b2 mbk_sig1306 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4141 mbk_sig1307 heart_block5_s35 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4142 heart_block5_a35s heart_block5_a5 mbk_sig1307 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4143 mbk_sig1303 heart_block5_s03 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4144 heart_block5_b03s heart_block5_b3 mbk_sig1303 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4145 vssi mbk_sig1296 heart_block5_m_2_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4146 mbk_sig1300 mbk_sig1296 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4147 heart_block5_m_2_2_dff_s mbk_sig1302 mbk_sig1300 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4148 vssi mbk_sig1301 heart_block5_m_2_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4149 vssi heart_block5_m_2_2_dff_m mbk_sig1296 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4150 heart_block5_m_2_2_dff_m heart_block5_ck2 mbk_sig1298 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4151 mbk_sig1302 heart_block5_ck2 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4152 vssi heart_block5_m_2_2_dff_s mbk_sig1301 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4153 heart_block5_s22 heart_block5_m_2_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4154 mbk_sig1298 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4155 mbk_sig1290 heart_block5_s34 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4156 heart_block5_a34s heart_block5_a4 mbk_sig1290 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4157 vssi mbk_sig1288 heart_block5_oa440s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4158 mbk_sig1288 heart_block5_a02s mbk_sig1291 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4159 mbk_sig1291 heart_block5_a03s mbk_sig1292 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4160 mbk_sig1292 heart_block5_a04s mbk_sig1286 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4161 mbk_sig1286 heart_block5_a01s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4162 vssi mbk_sig1280 heart_block5_m_3_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4163 mbk_sig1283 mbk_sig1280 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4164 heart_block5_m_3_0_dff_s mbk_sig1285 mbk_sig1283 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4165 vssi mbk_sig1284 heart_block5_m_3_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4166 vssi heart_block5_m_3_0_dff_m mbk_sig1280 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4167 heart_block5_m_3_0_dff_m heart_block5_ck3 mbk_sig1279 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4168 mbk_sig1285 heart_block5_ck3 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4169 vssi heart_block5_m_3_0_dff_s mbk_sig1284 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4170 heart_block5_s03 heart_block5_m_3_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4171 mbk_sig1279 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4172 vssi heart_block3_pb2 heart_block3_not2 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4173 vssi heart_block5_decalgra mbk_sig1220 vsse TN L=0.18U W=1.62U 
+ AS=0.5832P AD=0.5832P PS=3.96U PD=3.96U 
M4174 vssi mbk_sig1220 decalgrc vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M4175 decalgrc mbk_sig1220 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M4176 vssi heart_block3_pb0 heart_block3_not0 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4177 heart_block3_no31_csh heart_block3_pb3 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4178 vssi heart_block3_pb2 heart_block3_no31_csh vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4179 heart_block3_no31_csh heart_block3_gb1 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4180 heart_block3_no32_csh heart_block3_ngb3 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4181 vssi heart_block3_no31_csh heart_block3_no32_csh vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4182 heart_block3_no32_csh heart_block3_no2_csh vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4183 vssi heart_block3_gb3 heart_block3_ngb3 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4184 mbk_sig1218 ii_5 mbk_sig1216 vsse TN L=0.18U W=1.98U AS=0.7128P 
+ AD=0.7128P PS=4.68U PD=4.68U 
M4185 vssi ii_4 mbk_sig1218 vsse TN L=0.18U W=1.98U AS=0.7128P AD=0.7128P 
+ PS=4.68U PD=4.68U 
M4186 vssi ii_5 mbk_sig1217 vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M4187 mbk_sig1217 ii_4 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M4188 heart_block3_nn1 mbk_sig1216 mbk_sig1217 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4189 heart_block3_no22 heart_block3_gb2 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4190 vssi heart_block3_n2 heart_block3_no22 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4191 heart_block3_no32 heart_block3_pb2 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4192 vssi heart_block3_n3 heart_block3_no32 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4193 heart_block3_no20 heart_block3_gb0 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4194 vssi heart_block3_n2 heart_block3_no20 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4195 vssi heart_block3_nn0 heart_block3_n0 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4196 heart_block3_no30_csh heart_block3_pb1 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4197 vssi heart_block3_pb2 heart_block3_no30_csh vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4198 heart_block3_no30_csh heart_block3_pb3 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4199 mbk_sig1209 heart_block3_no22 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4200 vssi heart_block3_no32 mbk_sig1209 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4201 mbk_sig1211 heart_block3_no32 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4202 heart_block3_x22 heart_block3_no22 mbk_sig1211 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4203 vssi mbk_sig1209 heart_block3_x22 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4204 vssi mbk_sig1208 heart_block5_a213sh vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4205 mbk_sig1208 heart_block2_a25ms_i0 mbk_sig1207 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4206 mbk_sig1207 heart_block5_decalnr vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4207 vssi mbk_sig1205 heart_block5_shram0 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4208 mbk_sig1205 heart_block5_a214sh vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4209 vssi heart_block5_a213sh mbk_sig1205 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4210 mbk_sig1205 heart_block5_a212sh vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4211 vssi mbk_sig1204 heart_block5_a211sh vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4212 mbk_sig1204 heart_block2_a27ms_i0 mbk_sig1203 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4213 mbk_sig1203 heart_block5_decaldra vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4214 vssi mbk_sig1202 heart_block5_shram1 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4215 mbk_sig1202 heart_block5_a211sh vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4216 vssi heart_block5_a210sh mbk_sig1202 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4217 mbk_sig1202 heart_block5_a29sh vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4218 vssi mbk_sig1199 heart_block5_a210sh vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4219 mbk_sig1199 heart_block2_a26ms_i0 mbk_sig1200 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4220 mbk_sig1200 heart_block5_decalnr vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4221 vssi mbk_sig1197 heart_block5_a212sh vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4222 mbk_sig1197 r0i mbk_sig1198 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4223 mbk_sig1198 heart_block5_decalgra vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4224 vssi mbk_sig1194 heart_block5_a24sh vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4225 mbk_sig1194 heart_block2_a28ms_i0 mbk_sig1195 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4226 mbk_sig1195 heart_block5_decalnr vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4227 mbk_sig1192 ii_8 vssi vsse TN L=0.18U W=0.72U AS=0.2592P AD=0.2592P 
+ PS=2.16U PD=2.16U 
M4228 vssi heart_block4_ni7 mbk_sig1192 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4229 vssi mbk_sig1192 heart_block4_o21s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4230 vssi mbk_sig1191 heart_block5_decalgra vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4231 mbk_sig1191 ii_8 mbk_sig1193 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4232 mbk_sig1193 ii_7 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4233 vssi mbk_sig1190 heart_block5_shram3 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4234 mbk_sig1190 heart_block5_a25sh vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4235 vssi heart_block5_a24sh mbk_sig1190 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4236 mbk_sig1190 heart_block5_a23sh vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4237 vssi ii_7 heart_block4_ni7 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4238 vssi mbk_sig1186 heart_block5_a23sh vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4239 mbk_sig1186 heart_block2_a27ms_i0 mbk_sig1189 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4240 mbk_sig1189 heart_block5_decalgra vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4241 mbk_sig1185 heart_block5_s313 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4242 heart_block5_b313s heart_block5_b13 mbk_sig1185 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4243 mbk_sig1182 heart_block5_s36 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4244 heart_block5_b36s heart_block5_b6 mbk_sig1182 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4245 vssi mbk_sig1181 heart_block5_a25sh vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4246 mbk_sig1181 r3i mbk_sig1183 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4247 mbk_sig1183 heart_block5_decaldra vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4248 vssi mbk_sig1178 heart_block5_m_7_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4249 mbk_sig1176 mbk_sig1178 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4250 heart_block5_m_7_2_dff_s mbk_sig1177 mbk_sig1176 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4251 vssi mbk_sig1180 heart_block5_m_7_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4252 vssi heart_block5_m_7_2_dff_m mbk_sig1178 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4253 heart_block5_m_7_2_dff_m heart_block5_ck7 mbk_sig1174 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4254 mbk_sig1177 heart_block5_ck7 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4255 vssi heart_block5_m_7_2_dff_s mbk_sig1180 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4256 heart_block5_s27 heart_block5_m_7_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4257 mbk_sig1174 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4258 vssi mbk_sig1172 heart_block5_ck6 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4259 mbk_sig1172 heart_block5_enable mbk_sig1171 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4260 mbk_sig1171 heart_block5_b6 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4261 mbk_sig1169 heart_block5_s06 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4262 heart_block5_a06s heart_block5_a6 mbk_sig1169 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4263 vssi mbk_sig1162 heart_block5_m_6_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4264 mbk_sig1166 mbk_sig1162 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4265 heart_block5_m_6_1_dff_s mbk_sig1168 mbk_sig1166 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4266 vssi mbk_sig1167 heart_block5_m_6_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4267 vssi heart_block5_m_6_1_dff_m mbk_sig1162 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4268 heart_block5_m_6_1_dff_m heart_block5_ck6 mbk_sig1164 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4269 mbk_sig1168 heart_block5_ck6 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4270 vssi heart_block5_m_6_1_dff_s mbk_sig1167 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4271 heart_block5_s16 heart_block5_m_6_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4272 mbk_sig1164 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4273 vssi mbk_sig1159 heart_block5_oa432s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4274 mbk_sig1159 heart_block5_a26s mbk_sig1157 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4275 mbk_sig1157 heart_block5_a27s mbk_sig1158 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4276 mbk_sig1158 heart_block5_a28s mbk_sig1160 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4277 mbk_sig1160 heart_block5_a25s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4278 mbk_sig1156 heart_block5_s26 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4279 heart_block5_a26s heart_block5_a6 mbk_sig1156 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4280 mbk_sig1155 heart_block5_s27 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4281 heart_block5_a27s heart_block5_a7 mbk_sig1155 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4282 mbk_sig1153 heart_block5_s08 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4283 heart_block5_a08s heart_block5_a8 mbk_sig1153 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4284 mbk_sig1145 heart_block5_s16 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4285 heart_block5_a16s heart_block5_a6 mbk_sig1145 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4286 mbk_sig1147 heart_block5_s08 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4287 heart_block5_b08s heart_block5_b8 mbk_sig1147 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4288 vssi mbk_sig1138 heart_block5_m_5_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4289 mbk_sig1142 mbk_sig1138 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4290 heart_block5_m_5_0_dff_s mbk_sig1140 mbk_sig1142 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4291 vssi mbk_sig1144 heart_block5_m_5_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4292 vssi heart_block5_m_5_0_dff_m mbk_sig1138 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4293 heart_block5_m_5_0_dff_m heart_block5_ck5 mbk_sig1137 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4294 mbk_sig1140 heart_block5_ck5 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4295 vssi heart_block5_m_5_0_dff_s mbk_sig1144 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4296 heart_block5_s05 heart_block5_m_5_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4297 mbk_sig1137 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4298 mbk_sig1135 heart_block5_s35 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4299 heart_block5_b35s heart_block5_b5 mbk_sig1135 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4300 mbk_sig1132 heart_block5_s25 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4301 heart_block5_a25s heart_block5_a5 mbk_sig1132 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4302 vssi mbk_sig1127 heart_block5_m_11_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4303 mbk_sig1130 mbk_sig1127 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4304 heart_block5_m_11_3_dff_s mbk_sig1131 mbk_sig1130 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4305 vssi mbk_sig1133 heart_block5_m_11_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4306 vssi heart_block5_m_11_3_dff_m mbk_sig1127 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4307 heart_block5_m_11_3_dff_m heart_block5_ck11 mbk_sig1125 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4308 mbk_sig1131 heart_block5_ck11 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4309 vssi heart_block5_m_11_3_dff_s mbk_sig1133 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4310 heart_block5_s311 heart_block5_m_11_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4311 mbk_sig1125 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4312 vssi mbk_sig1118 heart_block5_m_5_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4313 mbk_sig1122 mbk_sig1118 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4314 heart_block5_m_5_3_dff_s mbk_sig1124 mbk_sig1122 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4315 vssi mbk_sig1123 heart_block5_m_5_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4316 vssi heart_block5_m_5_3_dff_m mbk_sig1118 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4317 heart_block5_m_5_3_dff_m heart_block5_ck5 mbk_sig1117 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4318 mbk_sig1124 heart_block5_ck5 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4319 vssi heart_block5_m_5_3_dff_s mbk_sig1123 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4320 heart_block5_s35 heart_block5_m_5_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4321 mbk_sig1117 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4322 vssi mbk_sig1111 heart_block5_m_2_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4323 mbk_sig1115 mbk_sig1111 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4324 heart_block5_m_2_0_dff_s mbk_sig1113 mbk_sig1115 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4325 vssi mbk_sig1116 heart_block5_m_2_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4326 vssi heart_block5_m_2_0_dff_m mbk_sig1111 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4327 heart_block5_m_2_0_dff_m heart_block5_ck2 mbk_sig1110 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4328 mbk_sig1113 heart_block5_ck2 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4329 vssi heart_block5_m_2_0_dff_s mbk_sig1116 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4330 heart_block5_s02 heart_block5_m_2_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4331 mbk_sig1110 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4332 vssi mbk_sig1107 heart_block5_m_2_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4333 mbk_sig1105 mbk_sig1107 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4334 heart_block5_m_2_1_dff_s mbk_sig1106 mbk_sig1105 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4335 vssi mbk_sig1109 heart_block5_m_2_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4336 vssi heart_block5_m_2_1_dff_m mbk_sig1107 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4337 heart_block5_m_2_1_dff_m heart_block5_ck2 mbk_sig1101 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4338 mbk_sig1106 heart_block5_ck2 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4339 vssi heart_block5_m_2_1_dff_s mbk_sig1109 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4340 heart_block5_s12 heart_block5_m_2_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4341 mbk_sig1101 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4342 mbk_sig1102 heart_block5_s12 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4343 heart_block5_a12s heart_block5_a2 mbk_sig1102 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4344 mbk_sig1098 heart_block5_s310 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4345 heart_block5_b310s heart_block5_b10 mbk_sig1098 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4346 vssi mbk_sig1097 heart_block5_ck10 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4347 mbk_sig1097 heart_block5_enable mbk_sig1099 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4348 mbk_sig1099 heart_block5_b10 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4349 vssi mbk_sig1090 heart_block5_m_10_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4350 mbk_sig1094 mbk_sig1090 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4351 heart_block5_m_10_3_dff_s mbk_sig1095 mbk_sig1094 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4352 vssi mbk_sig1096 heart_block5_m_10_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4353 vssi heart_block5_m_10_3_dff_m mbk_sig1090 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4354 heart_block5_m_10_3_dff_m heart_block5_ck10 mbk_sig1092 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4355 mbk_sig1095 heart_block5_ck10 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4356 vssi heart_block5_m_10_3_dff_s mbk_sig1096 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4357 heart_block5_s310 heart_block5_m_10_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4358 mbk_sig1092 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4359 mbk_sig1087 heart_block5_s02 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4360 heart_block5_a02s heart_block5_a2 mbk_sig1087 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4361 mbk_sig1086 heart_block5_s010 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4362 heart_block5_a010s heart_block5_a10 mbk_sig1086 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4363 mbk_sig1055 heart_block3_x10 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4364 heart_block3_gb0 heart_block3_x00 mbk_sig1055 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4365 mbk_sig1053 heart_block3_cout2 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4366 heart_block3_na23 heart_block3_not3 mbk_sig1053 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4367 mbk_sig1054 heart_block3_na23 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4368 heart_block3_couta heart_block3_gb3 mbk_sig1054 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4369 heart_block3_no30 heart_block3_pb0 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4370 vssi heart_block3_n3 heart_block3_no30 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4371 vssi mbk_sig1050 heart_s_1 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4372 mbk_sig1050 heart_block1_srq1 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4373 vssi heart_block1_sra1 mbk_sig1050 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4374 mbk_sig1050 heart_block1_srb1 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4375 mbk_sig1049 heart_s_1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4376 vssi heart_block3_n1 mbk_sig1049 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4377 mbk_sig1047 heart_block3_n1 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4378 heart_block3_x11 heart_s_1 mbk_sig1047 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4379 vssi mbk_sig1049 heart_block3_x11 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4380 mbk_sig1046 heart_block3_cout2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4381 vssi heart_block3_couta mbk_sig1046 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4382 mbk_sig1045 heart_block3_couta vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4383 ovrc heart_block3_cout2 mbk_sig1045 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4384 vssi mbk_sig1046 ovrc vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4385 vssi mbk_sig1042 heart_block1_srq1 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4386 mbk_sig1042 heart_q_1 mbk_sig1041 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4387 mbk_sig1041 heart_block1_selqs vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4388 heart_block3_no2_csh heart_block3_pb3 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4389 vssi heart_block3_gb2 heart_block3_no2_csh vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4390 vssi heart_block3_gb0 heart_block3_ngb0 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4391 vssi heart_block3_p npc vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4392 vssi mbk_sig1037 coutc vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4393 mbk_sig1037 heart_block3_couta mbk_sig1036 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4394 mbk_sig1036 heart_block3_flag vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4395 vssi heart_block3_nprop heart_block3_propf vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4396 vssi heart_block5_decaldra mbk_sig1035 vsse TN L=0.18U W=1.62U 
+ AS=0.5832P AD=0.5832P PS=3.96U PD=3.96U 
M4397 vssi mbk_sig1035 decaldrc vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M4398 decaldrc mbk_sig1035 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M4399 vssi mbk_sig1034 heart_block3_p vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4400 mbk_sig1034 heart_block3_propf mbk_sig1033 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4401 mbk_sig1033 heart_block3_flag vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4402 vssi ii_7 heart_block5_ni7 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4403 vssi mbk_sig1030 heart_block2_syalu3 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4404 mbk_sig1030 heart_block2_a28ms_i0 mbk_sig1029 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4405 mbk_sig1029 heart_block2_selaluy vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4406 vssi mbk_sig1028 heart_block5_decaldra vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4407 mbk_sig1028 ii_8 mbk_sig1027 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4408 mbk_sig1027 heart_block5_ni7 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4409 mbk_sig1023 heart_block2_syra3 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4410 vssi heart_block2_syalu3 mbk_sig1023 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4411 vssi mbk_sig1023 yc_3 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4412 vssi mbk_sig1022 s0c vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4413 mbk_sig1022 heart_block5_decaldra mbk_sig1024 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4414 mbk_sig1024 heart_block2_a25ms_i0 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4415 vssi mbk_sig1020 heart_block1_srq0 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4416 mbk_sig1020 heart_q_0 mbk_sig1019 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4417 mbk_sig1019 heart_block1_selqs vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4418 vssi mbk_sig1016 heart_block4_decalga vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4419 mbk_sig1016 ii_8 mbk_sig1018 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4420 mbk_sig1018 ii_7 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4421 vssi mbk_sig1013 heart_block1_srb3 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4422 mbk_sig1013 heart_rb_3 mbk_sig1014 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4423 mbk_sig1014 heart_block1_selbs vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4424 vssi mbk_sig1012 heart_block5_ck16 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4425 mbk_sig1012 heart_block5_enable mbk_sig1015 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4426 mbk_sig1015 heart_block5_b16 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4427 vssi mbk_sig1011 heart_block5_ck13 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4428 mbk_sig1011 heart_block5_enable mbk_sig1010 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4429 mbk_sig1010 heart_block5_b13 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4430 mbk_sig1009 heart_block5_s113 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4431 heart_block5_b113s heart_block5_b13 mbk_sig1009 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4432 mbk_sig1006 heart_block5_s116 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4433 heart_block5_b116s heart_block5_b16 mbk_sig1006 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4434 vssi mbk_sig1002 heart_block5_m_6_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4435 mbk_sig1003 mbk_sig1002 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4436 heart_block5_m_6_0_dff_s mbk_sig1004 mbk_sig1003 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4437 vssi mbk_sig1008 heart_block5_m_6_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4438 vssi heart_block5_m_6_0_dff_m mbk_sig1002 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4439 heart_block5_m_6_0_dff_m heart_block5_ck6 mbk_sig1000 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4440 mbk_sig1004 heart_block5_ck6 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4441 vssi heart_block5_m_6_0_dff_s mbk_sig1008 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4442 heart_block5_s06 heart_block5_m_6_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4443 mbk_sig1000 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4444 mbk_sig1001 heart_block5_s316 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4445 heart_block5_b316s heart_block5_b16 mbk_sig1001 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4446 vssi mbk_sig994 heart_block5_ob413s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4447 mbk_sig994 heart_block5_b314s mbk_sig996 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4448 mbk_sig996 heart_block5_b315s mbk_sig997 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4449 mbk_sig997 heart_block5_b316s mbk_sig998 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4450 mbk_sig998 heart_block5_b313s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4451 vssi mbk_sig990 heart_block5_m_16_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4452 mbk_sig991 mbk_sig990 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4453 heart_block5_m_16_3_dff_s mbk_sig989 mbk_sig991 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4454 vssi mbk_sig993 heart_block5_m_16_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4455 vssi heart_block5_m_16_3_dff_m mbk_sig990 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4456 heart_block5_m_16_3_dff_m heart_block5_ck16 mbk_sig987 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4457 mbk_sig989 heart_block5_ck16 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4458 vssi heart_block5_m_16_3_dff_s mbk_sig993 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4459 heart_block5_s316 heart_block5_m_16_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4460 mbk_sig987 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4461 mbk_sig982 heart_block5_ob442s vssi vsse TN L=0.18U W=4.32U AS=1.5552P 
+ AD=1.5552P PS=9.36U PD=9.36U 
M4462 mbk_sig986 heart_block5_ob432s mbk_sig982 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4463 mbk_sig985 heart_block5_ob422s mbk_sig986 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4464 heart_rb_2 heart_block5_ob412s mbk_sig985 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4465 mbk_sig981 heart_block5_s315 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4466 heart_block5_b315s heart_block5_b15 mbk_sig981 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4467 vssi mbk_sig974 heart_block5_ob433s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4468 mbk_sig974 heart_block5_b36s mbk_sig975 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4469 mbk_sig975 heart_block5_b37s mbk_sig976 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4470 mbk_sig976 heart_block5_b38s mbk_sig977 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4471 mbk_sig977 heart_block5_b35s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4472 vssi mbk_sig971 heart_block5_m_7_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4473 mbk_sig969 mbk_sig971 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4474 heart_block5_m_7_3_dff_s mbk_sig970 mbk_sig969 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4475 vssi mbk_sig973 heart_block5_m_7_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4476 vssi heart_block5_m_7_3_dff_m mbk_sig971 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4477 heart_block5_m_7_3_dff_m heart_block5_ck7 mbk_sig967 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4478 mbk_sig970 heart_block5_ck7 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4479 vssi heart_block5_m_7_3_dff_s mbk_sig973 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4480 heart_block5_s37 heart_block5_m_7_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4481 mbk_sig967 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4482 mbk_sig962 heart_block5_ob443s vssi vsse TN L=0.18U W=4.32U AS=1.5552P 
+ AD=1.5552P PS=9.36U PD=9.36U 
M4483 mbk_sig963 heart_block5_ob433s mbk_sig962 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4484 mbk_sig966 heart_block5_ob423s mbk_sig963 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4485 heart_rb_3 heart_block5_ob413s mbk_sig966 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4486 vssi mbk_sig955 heart_block5_m_11_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4487 mbk_sig958 mbk_sig955 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4488 heart_block5_m_11_2_dff_s mbk_sig960 mbk_sig958 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4489 vssi mbk_sig961 heart_block5_m_11_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4490 vssi heart_block5_m_11_2_dff_m mbk_sig955 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4491 heart_block5_m_11_2_dff_m heart_block5_ck11 mbk_sig957 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4492 mbk_sig960 heart_block5_ck11 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4493 vssi heart_block5_m_11_2_dff_s mbk_sig961 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4494 heart_block5_s211 heart_block5_m_11_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4495 mbk_sig957 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4496 mbk_sig954 heart_block5_s211 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4497 heart_block5_b211s heart_block5_b11 mbk_sig954 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4498 vssi mbk_sig952 heart_block5_a3 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4499 mbk_sig952 heart_a_1 mbk_sig953 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4500 mbk_sig953 heart_block5_na2 mbk_sig950 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4501 mbk_sig950 heart_block5_na3 mbk_sig951 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4502 mbk_sig951 heart_block5_na0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4503 vssi mbk_sig948 heart_block5_a5 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4504 mbk_sig948 heart_block5_na1 mbk_sig946 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4505 mbk_sig946 heart_a_2 mbk_sig947 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4506 mbk_sig947 heart_block5_na3 mbk_sig945 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4507 mbk_sig945 heart_block5_na0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4508 mbk_sig941 heart_block5_s37 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4509 heart_block5_a37s heart_block5_a7 mbk_sig941 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4510 mbk_sig942 heart_block5_s29 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4511 heart_block5_b29s heart_block5_b9 mbk_sig942 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4512 vssi mbk_sig937 heart_block5_ob422s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4513 mbk_sig937 heart_block5_b210s mbk_sig938 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4514 mbk_sig938 heart_block5_b211s mbk_sig939 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4515 mbk_sig939 heart_block5_b212s mbk_sig940 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4516 mbk_sig940 heart_block5_b29s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4517 vssi mbk_sig933 heart_block5_a7 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4518 mbk_sig933 heart_a_1 mbk_sig934 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4519 mbk_sig934 heart_a_2 mbk_sig935 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4520 mbk_sig935 heart_block5_na3 mbk_sig936 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4521 mbk_sig936 heart_block5_na0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4522 mbk_sig932 heart_block5_s210 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4523 heart_block5_b210s heart_block5_b10 mbk_sig932 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4524 mbk_sig930 heart_block5_s311 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4525 heart_block5_b311s heart_block5_b11 mbk_sig930 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4526 vssi mbk_sig927 heart_block5_a4 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4527 mbk_sig927 heart_a_1 mbk_sig928 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4528 mbk_sig928 heart_block5_na2 mbk_sig929 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4529 mbk_sig929 heart_block5_na3 mbk_sig926 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4530 mbk_sig926 heart_a_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M4531 mbk_sig925 heart_block5_s311 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4532 heart_block5_a311s heart_block5_a11 mbk_sig925 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4533 vssi mbk_sig918 heart_block5_ob423s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4534 mbk_sig918 heart_block5_b310s mbk_sig919 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4535 mbk_sig919 heart_block5_b311s mbk_sig920 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4536 mbk_sig920 heart_block5_b312s mbk_sig921 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4537 mbk_sig921 heart_block5_b39s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4538 vssi mbk_sig915 heart_block5_m_10_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4539 mbk_sig913 mbk_sig915 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4540 heart_block5_m_10_0_dff_s mbk_sig914 mbk_sig913 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4541 vssi mbk_sig917 heart_block5_m_10_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4542 vssi heart_block5_m_10_0_dff_m mbk_sig915 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4543 heart_block5_m_10_0_dff_m heart_block5_ck10 mbk_sig911 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4544 mbk_sig914 heart_block5_ck10 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4545 vssi heart_block5_m_10_0_dff_s mbk_sig917 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4546 heart_block5_s010 heart_block5_m_10_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4547 mbk_sig911 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4548 vssi mbk_sig906 heart_block5_m_10_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4549 mbk_sig907 mbk_sig906 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4550 heart_block5_m_10_1_dff_s mbk_sig908 mbk_sig907 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4551 vssi mbk_sig910 heart_block5_m_10_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4552 vssi heart_block5_m_10_1_dff_m mbk_sig906 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4553 heart_block5_m_10_1_dff_m heart_block5_ck10 mbk_sig905 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4554 mbk_sig908 heart_block5_ck10 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4555 vssi heart_block5_m_10_1_dff_s mbk_sig910 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4556 heart_block5_s110 heart_block5_m_10_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4557 mbk_sig905 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4558 mbk_sig866 heart_r_0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4559 vssi heart_block3_n0 mbk_sig866 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4560 mbk_sig869 heart_block3_n0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4561 heart_block3_x00 heart_r_0 mbk_sig869 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4562 vssi mbk_sig866 heart_block3_x00 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4563 heart_block3_pb0 heart_block3_x10 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4564 vssi heart_block3_x00 heart_block3_pb0 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4565 vssi heart_block3_pb3 heart_block3_not3 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4566 vssi mbk_sig861 heart_block3_ngen vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4567 mbk_sig861 heart_block3_na_csh mbk_sig862 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4568 mbk_sig862 heart_block3_no32_csh vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4569 mbk_sig858 heart_block3_no30_csh vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4570 heart_block3_na_csh heart_block3_ngb0 mbk_sig858 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4571 heart_block3_pb2 heart_block3_x12 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4572 vssi heart_block3_x02 heart_block3_pb2 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4573 mbk_sig853 heart_r_3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4574 vssi heart_block3_n0 mbk_sig853 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4575 mbk_sig852 heart_block3_n0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4576 heart_block3_x03 heart_r_3 mbk_sig852 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4577 vssi mbk_sig853 heart_block3_x03 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4578 heart_block3_pb3 heart_block3_x13 vssi vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4579 vssi heart_block3_x03 heart_block3_pb3 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4580 mbk_sig848 heart_block3_x13 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4581 heart_block3_gb3 heart_block3_x03 mbk_sig848 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4582 vssi heart_block3_ngen heart_block3_genf vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4583 vssi mbk_sig844 heart_block3_g vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4584 mbk_sig844 heart_block3_genf mbk_sig845 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4585 mbk_sig845 heart_block3_flag vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4586 mbk_sig841 heart_block3_no30_csh vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4587 heart_block3_nprop heart_block3_npb0 mbk_sig841 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4588 mbk_sig837 heart_s_3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4589 vssi heart_block3_n1 mbk_sig837 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4590 mbk_sig842 heart_block3_n1 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4591 heart_block3_x13 heart_s_3 mbk_sig842 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4592 vssi mbk_sig837 heart_block3_x13 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4593 vssi mbk_sig832 heart_s_3 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4594 mbk_sig832 heart_block1_srq3 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4595 vssi heart_block1_sra3 mbk_sig832 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4596 mbk_sig832 heart_block1_srb3 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4597 vssi mbk_sig830 heart_block1_srq3 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4598 mbk_sig830 heart_q_3 mbk_sig831 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4599 mbk_sig831 heart_block1_selqs vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4600 vssi mbk_sig824 heart_block5_m_13_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4601 mbk_sig828 mbk_sig824 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4602 heart_block5_m_13_0_dff_s mbk_sig826 mbk_sig828 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4603 vssi mbk_sig829 heart_block5_m_13_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4604 vssi heart_block5_m_13_0_dff_m mbk_sig824 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4605 heart_block5_m_13_0_dff_m heart_block5_ck13 mbk_sig822 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4606 mbk_sig826 heart_block5_ck13 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4607 vssi heart_block5_m_13_0_dff_s mbk_sig829 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4608 heart_block5_s013 heart_block5_m_13_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4609 mbk_sig822 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4610 vssi mbk_sig815 heart_block5_m_13_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4611 mbk_sig820 mbk_sig815 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4612 heart_block5_m_13_2_dff_s mbk_sig821 mbk_sig820 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4613 vssi mbk_sig823 heart_block5_m_13_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4614 vssi heart_block5_m_13_2_dff_m mbk_sig815 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4615 heart_block5_m_13_2_dff_m heart_block5_ck13 mbk_sig818 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4616 mbk_sig821 heart_block5_ck13 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4617 vssi heart_block5_m_13_2_dff_s mbk_sig823 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4618 heart_block5_s213 heart_block5_m_13_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4619 mbk_sig818 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4620 mbk_sig817 heart_block5_s213 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4621 heart_block5_a213s heart_block5_a13 mbk_sig817 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4622 vssi mbk_sig812 heart_block5_m_16_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4623 mbk_sig810 mbk_sig812 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4624 heart_block5_m_16_1_dff_s mbk_sig811 mbk_sig810 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4625 vssi mbk_sig814 heart_block5_m_16_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4626 vssi heart_block5_m_16_1_dff_m mbk_sig812 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4627 heart_block5_m_16_1_dff_m heart_block5_ck16 mbk_sig808 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4628 mbk_sig811 heart_block5_ck16 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4629 vssi heart_block5_m_16_1_dff_s mbk_sig814 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4630 heart_block5_s116 heart_block5_m_16_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4631 mbk_sig808 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4632 mbk_sig809 heart_block5_s214 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4633 heart_block5_b214s heart_block5_b14 mbk_sig809 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4634 mbk_sig805 heart_block5_s113 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4635 heart_block5_a113s heart_block5_a13 mbk_sig805 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4636 mbk_sig806 heart_block5_s213 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4637 heart_block5_b213s heart_block5_b13 mbk_sig806 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4638 vssi mbk_sig801 heart_block5_m_6_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4639 mbk_sig799 mbk_sig801 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4640 heart_block5_m_6_2_dff_s mbk_sig800 mbk_sig799 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4641 vssi mbk_sig804 heart_block5_m_6_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4642 vssi heart_block5_m_6_2_dff_m mbk_sig801 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4643 heart_block5_m_6_2_dff_m heart_block5_ck6 mbk_sig796 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4644 mbk_sig800 heart_block5_ck6 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4645 vssi heart_block5_m_6_2_dff_s mbk_sig804 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4646 heart_block5_s26 heart_block5_m_6_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4647 mbk_sig796 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4648 mbk_sig797 heart_block5_s216 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4649 heart_block5_b216s heart_block5_b16 mbk_sig797 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4650 vssi mbk_sig793 heart_block5_ob412s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4651 mbk_sig793 heart_block5_b214s mbk_sig791 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4652 mbk_sig791 heart_block5_b215s mbk_sig792 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4653 mbk_sig792 heart_block5_b216s mbk_sig794 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4654 mbk_sig794 heart_block5_b213s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4655 mbk_sig788 heart_block5_s216 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4656 heart_block5_a216s heart_block5_a16 mbk_sig788 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4657 vssi mbk_sig787 heart_block5_oa412s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4658 mbk_sig787 heart_block5_a214s mbk_sig789 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4659 mbk_sig789 heart_block5_a215s mbk_sig786 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4660 mbk_sig786 heart_block5_a216s mbk_sig785 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4661 mbk_sig785 heart_block5_a213s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4662 mbk_sig707 heart_block5_ob440s vssi vsse TN L=0.18U W=4.32U AS=1.5552P 
+ AD=1.5552P PS=9.36U PD=9.36U 
M4663 mbk_sig708 heart_block5_ob430s mbk_sig707 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4664 mbk_sig709 heart_block5_ob420s mbk_sig708 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4665 heart_rb_0 heart_block5_ob410s mbk_sig709 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4666 mbk_sig782 heart_block5_s115 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4667 heart_block5_b115s heart_block5_b15 mbk_sig782 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4668 vssi mbk_sig779 heart_block5_ob411s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4669 mbk_sig779 heart_block5_b114s mbk_sig783 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4670 mbk_sig783 heart_block5_b115s mbk_sig784 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4671 mbk_sig784 heart_block5_b116s mbk_sig778 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4672 mbk_sig778 heart_block5_b113s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4673 mbk_sig702 heart_block5_oa440s vssi vsse TN L=0.18U W=4.32U AS=1.5552P 
+ AD=1.5552P PS=9.36U PD=9.36U 
M4674 mbk_sig703 heart_block5_oa430s mbk_sig702 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4675 mbk_sig706 heart_block5_oa420s mbk_sig703 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4676 heart_ra_0 heart_block5_oa410s mbk_sig706 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4677 mbk_sig772 heart_block5_s37 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4678 heart_block5_b37s heart_block5_b7 mbk_sig772 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4679 vssi mbk_sig773 heart_block5_ck15 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4680 mbk_sig773 heart_block5_enable mbk_sig774 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4681 mbk_sig774 heart_block5_b15 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4682 vssi mbk_sig768 heart_block5_a8 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4683 mbk_sig768 heart_a_1 mbk_sig769 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4684 mbk_sig769 heart_a_2 mbk_sig770 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4685 mbk_sig770 heart_block5_na3 mbk_sig771 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4686 mbk_sig771 heart_a_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M4687 vssi mbk_sig764 heart_block5_m_15_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4688 mbk_sig762 mbk_sig764 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4689 heart_block5_m_15_1_dff_s mbk_sig763 mbk_sig762 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4690 vssi mbk_sig767 heart_block5_m_15_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4691 vssi heart_block5_m_15_1_dff_m mbk_sig764 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4692 heart_block5_m_15_1_dff_m heart_block5_ck15 mbk_sig759 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4693 mbk_sig763 heart_block5_ck15 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4694 vssi heart_block5_m_15_1_dff_s mbk_sig767 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4695 heart_block5_s115 heart_block5_m_15_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4696 mbk_sig759 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4697 vssi mbk_sig758 heart_block5_ck11 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4698 mbk_sig758 heart_block5_enable mbk_sig761 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4699 mbk_sig761 heart_block5_b11 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4700 vssi mbk_sig755 heart_block5_m_9_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4701 mbk_sig753 mbk_sig755 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4702 heart_block5_m_9_3_dff_s mbk_sig754 mbk_sig753 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4703 vssi mbk_sig757 heart_block5_m_9_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4704 vssi heart_block5_m_9_3_dff_m mbk_sig755 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4705 heart_block5_m_9_3_dff_m heart_block5_ck9 mbk_sig750 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4706 mbk_sig754 heart_block5_ck9 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4707 vssi heart_block5_m_9_3_dff_s mbk_sig757 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4708 heart_block5_s39 heart_block5_m_9_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4709 mbk_sig750 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4710 vssi mbk_sig749 heart_block5_a1 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4711 mbk_sig749 heart_block5_na1 mbk_sig752 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4712 mbk_sig752 heart_block5_na2 mbk_sig747 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4713 mbk_sig747 heart_block5_na3 mbk_sig746 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4714 mbk_sig746 heart_block5_na0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4715 vssi mbk_sig738 heart_block5_m_10_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4716 mbk_sig743 mbk_sig738 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4717 heart_block5_m_10_2_dff_s mbk_sig745 mbk_sig743 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4718 vssi mbk_sig744 heart_block5_m_10_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4719 vssi heart_block5_m_10_2_dff_m mbk_sig738 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4720 heart_block5_m_10_2_dff_m heart_block5_ck10 mbk_sig740 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4721 mbk_sig745 heart_block5_ck10 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4722 vssi heart_block5_m_10_2_dff_s mbk_sig744 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4723 heart_block5_s210 heart_block5_m_10_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4724 mbk_sig740 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4725 vssi mbk_sig736 heart_block5_a13 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4726 mbk_sig736 heart_block5_na1 mbk_sig734 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4727 mbk_sig734 heart_a_2 mbk_sig735 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4728 mbk_sig735 heart_a_3 mbk_sig737 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4729 mbk_sig737 heart_block5_na0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4730 mbk_sig733 heart_block5_s39 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4731 heart_block5_b39s heart_block5_b9 mbk_sig733 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4732 vssi heart_a_1 heart_block5_na1 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4733 mbk_sig730 heart_block5_s210 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4734 heart_block5_a210s heart_block5_a10 mbk_sig730 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4735 vssi mbk_sig729 heart_block5_a2 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4736 mbk_sig729 heart_block5_na1 mbk_sig727 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4737 mbk_sig727 heart_block5_na2 mbk_sig728 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4738 mbk_sig728 heart_block5_na3 mbk_sig726 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4739 mbk_sig726 heart_a_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M4740 mbk_sig722 heart_block5_s312 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4741 heart_block5_b312s heart_block5_b12 mbk_sig722 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4742 vssi mbk_sig721 heart_block5_a10 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4743 mbk_sig721 heart_block5_na1 mbk_sig723 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4744 mbk_sig723 heart_block5_na2 mbk_sig720 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4745 mbk_sig720 heart_a_3 mbk_sig719 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4746 mbk_sig719 heart_a_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M4747 mbk_sig717 heart_block5_s010 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4748 heart_block5_b010s heart_block5_b10 mbk_sig717 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4749 vssi heart_a_0 heart_block5_na0 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4750 mbk_sig667 heart_s_2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4751 vssi heart_block3_n1 mbk_sig667 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4752 mbk_sig666 heart_block3_n1 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4753 heart_block3_x12 heart_s_2 mbk_sig666 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4754 vssi mbk_sig667 heart_block3_x12 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4755 vssi heart_block3_nn1 heart_block3_n1 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4756 vssi mbk_sig663 heart_s_0 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4757 mbk_sig663 heart_block1_srq0 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4758 vssi heart_block1_sra0 mbk_sig663 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4759 mbk_sig663 heart_block1_srb0 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4760 mbk_sig662 heart_s_0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4761 vssi heart_block3_n1 mbk_sig662 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4762 mbk_sig661 heart_block3_n1 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4763 heart_block3_x10 heart_s_0 mbk_sig661 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4764 vssi mbk_sig662 heart_block3_x10 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4765 vssi heart_block3_pb0 heart_block3_npb0 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4766 vssi mbk_sig656 heart_block1_sra0 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4767 mbk_sig656 heart_ra_0 mbk_sig655 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4768 mbk_sig655 heart_block1_selas vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4769 vssi mbk_sig654 heart_block4_ckin vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4770 mbk_sig654 cko mbk_sig653 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4771 mbk_sig653 heart_block4_w vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4772 mbk_sig650 heart_block3_x12 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4773 heart_block3_gb2 heart_block3_x02 mbk_sig650 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4774 mbk_sig648 heart_block4_test_mode vssi vsse TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
M4775 vssi heart_block4_a231s mbk_sig648 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4776 vssi mbk_sig648 heart_block4_w vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4777 vssi mbk_sig646 heart_fonc_mode vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4778 mbk_sig646 fonci mbk_sig647 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4779 mbk_sig647 heart_block4_n15s vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4780 vssi ii_6 heart_block4_ni6 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4781 vssi mbk_sig642 heart_block4_a231s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4782 mbk_sig642 heart_fonc_mode mbk_sig643 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4783 mbk_sig643 heart_block4_waccu vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4784 vssi mbk_sig641 heart_block4_waccu vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4785 mbk_sig641 heart_block4_o21s mbk_sig644 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4786 mbk_sig644 heart_block4_ni6 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4787 vssi fonci heart_block4_n14s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4788 vssi mbk_sig639 heart_block2_syra3 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4789 mbk_sig639 heart_ra_3 mbk_sig638 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4790 mbk_sig638 heart_block2_selray vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4791 vssi mbk_sig634 heart_block2_syalu2 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4792 mbk_sig634 heart_block2_a27ms_i0 mbk_sig635 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4793 mbk_sig635 heart_block2_selaluy vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4794 mbk_sig631 heart_block5_s313 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4795 heart_block5_a313s heart_block5_a13 mbk_sig631 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4796 vssi mbk_sig630 heart_block2_syalu0 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4797 mbk_sig630 heart_block2_a25ms_i0 mbk_sig632 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4798 mbk_sig632 heart_block2_selaluy vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4799 vssi mbk_sig628 heart_block2_syra0 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4800 mbk_sig628 heart_ra_0 mbk_sig629 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4801 mbk_sig629 heart_block2_selray vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4802 mbk_sig624 heart_block2_syra0 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4803 vssi heart_block2_syalu0 mbk_sig624 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4804 vssi mbk_sig624 yc_0 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4805 vssi mbk_sig623 heart_block1_srb2 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4806 mbk_sig623 heart_rb_2 mbk_sig625 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4807 mbk_sig625 heart_block1_selbs vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4808 vssi mbk_sig621 heart_block1_srb0 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4809 mbk_sig621 heart_rb_0 mbk_sig620 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4810 mbk_sig620 heart_block1_selbs vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4811 vssi mbk_sig612 heart_block5_m_13_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4812 mbk_sig617 mbk_sig612 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4813 heart_block5_m_13_1_dff_s mbk_sig614 mbk_sig617 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4814 vssi mbk_sig619 heart_block5_m_13_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4815 vssi heart_block5_m_13_1_dff_m mbk_sig612 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4816 heart_block5_m_13_1_dff_m heart_block5_ck13 mbk_sig609 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4817 mbk_sig614 heart_block5_ck13 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4818 vssi heart_block5_m_13_1_dff_s mbk_sig619 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4819 heart_block5_s113 heart_block5_m_13_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4820 mbk_sig609 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4821 vssi mbk_sig610 heart_block1_srb1 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4822 mbk_sig610 heart_rb_1 mbk_sig611 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4823 mbk_sig611 heart_block1_selbs vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4824 mbk_sig606 heart_block5_s013 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4825 heart_block5_a013s heart_block5_a13 mbk_sig606 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4826 vssi mbk_sig605 heart_block5_ob410s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4827 mbk_sig605 heart_block5_b014s mbk_sig602 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4828 mbk_sig602 heart_block5_b015s mbk_sig603 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4829 mbk_sig603 heart_block5_b016s mbk_sig601 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4830 mbk_sig601 heart_block5_b013s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4831 vssi mbk_sig593 heart_block5_m_16_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4832 mbk_sig597 mbk_sig593 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4833 heart_block5_m_16_2_dff_s mbk_sig595 mbk_sig597 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4834 vssi mbk_sig599 heart_block5_m_16_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4835 vssi heart_block5_m_16_2_dff_m mbk_sig593 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4836 heart_block5_m_16_2_dff_m heart_block5_ck16 mbk_sig596 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4837 mbk_sig595 heart_block5_ck16 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4838 vssi heart_block5_m_16_2_dff_s mbk_sig599 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4839 heart_block5_s216 heart_block5_m_16_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4840 mbk_sig596 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4841 mbk_sig591 heart_block5_s214 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4842 heart_block5_a214s heart_block5_a14 mbk_sig591 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4843 vssi mbk_sig589 heart_block5_oa413s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4844 mbk_sig589 heart_block5_a314s mbk_sig590 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4845 mbk_sig590 heart_block5_a315s mbk_sig587 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4846 mbk_sig587 heart_block5_a316s mbk_sig586 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4847 mbk_sig586 heart_block5_a313s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4848 mbk_sig588 heart_block5_s316 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4849 heart_block5_a316s heart_block5_a16 mbk_sig588 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4850 mbk_sig582 heart_block5_s013 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4851 heart_block5_b013s heart_block5_b13 mbk_sig582 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4852 mbk_sig579 heart_block5_s315 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4853 heart_block5_a315s heart_block5_a15 mbk_sig579 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4854 mbk_sig580 heart_block5_s115 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4855 heart_block5_a115s heart_block5_a15 mbk_sig580 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4856 mbk_sig575 heart_block5_s215 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4857 heart_block5_b215s heart_block5_b15 mbk_sig575 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4858 mbk_sig570 heart_block5_ob441s vssi vsse TN L=0.18U W=4.32U AS=1.5552P 
+ AD=1.5552P PS=9.36U PD=9.36U 
M4859 mbk_sig571 heart_block5_ob431s mbk_sig570 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4860 mbk_sig576 heart_block5_ob421s mbk_sig571 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4861 heart_rb_1 heart_block5_ob411s mbk_sig576 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4862 vssi mbk_sig569 heart_block5_ck9 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4863 mbk_sig569 heart_block5_enable mbk_sig572 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4864 mbk_sig572 heart_block5_b9 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4865 vssi mbk_sig566 heart_block5_a16 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4866 mbk_sig566 heart_a_1 mbk_sig567 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4867 mbk_sig567 heart_a_2 mbk_sig568 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4868 mbk_sig568 heart_a_3 mbk_sig564 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4869 mbk_sig564 heart_a_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M4870 mbk_sig560 heart_block5_oa441s vssi vsse TN L=0.18U W=4.32U AS=1.5552P 
+ AD=1.5552P PS=9.36U PD=9.36U 
M4871 mbk_sig561 heart_block5_oa431s mbk_sig560 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4872 mbk_sig565 heart_block5_oa421s mbk_sig561 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4873 heart_ra_1 heart_block5_oa411s mbk_sig565 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4874 vssi mbk_sig553 heart_block5_m_15_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4875 mbk_sig556 mbk_sig553 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4876 heart_block5_m_15_2_dff_s mbk_sig558 mbk_sig556 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4877 vssi mbk_sig559 heart_block5_m_15_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4878 vssi heart_block5_m_15_2_dff_m mbk_sig553 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4879 heart_block5_m_15_2_dff_m heart_block5_ck15 mbk_sig555 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4880 mbk_sig558 heart_block5_ck15 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4881 vssi heart_block5_m_15_2_dff_s mbk_sig559 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4882 heart_block5_s215 heart_block5_m_15_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4883 mbk_sig555 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4884 vssi mbk_sig546 heart_block5_m_15_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4885 mbk_sig549 mbk_sig546 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4886 heart_block5_m_15_3_dff_s mbk_sig548 mbk_sig549 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4887 vssi mbk_sig552 heart_block5_m_15_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4888 vssi heart_block5_m_15_3_dff_m mbk_sig546 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4889 heart_block5_m_15_3_dff_m heart_block5_ck15 mbk_sig543 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4890 mbk_sig548 heart_block5_ck15 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4891 vssi heart_block5_m_15_3_dff_s mbk_sig552 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4892 heart_block5_s315 heart_block5_m_15_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4893 mbk_sig543 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4894 vssi mbk_sig542 heart_block5_m_9_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4895 mbk_sig540 mbk_sig542 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4896 heart_block5_m_9_2_dff_s mbk_sig541 mbk_sig540 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4897 vssi mbk_sig545 heart_block5_m_9_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4898 vssi heart_block5_m_9_2_dff_m mbk_sig542 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4899 heart_block5_m_9_2_dff_m heart_block5_ck9 mbk_sig539 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4900 mbk_sig541 heart_block5_ck9 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4901 vssi heart_block5_m_9_2_dff_s mbk_sig545 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4902 heart_block5_s29 heart_block5_m_9_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4903 mbk_sig539 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4904 vssi mbk_sig536 heart_block5_a6 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4905 mbk_sig536 heart_block5_na1 mbk_sig538 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4906 mbk_sig538 heart_a_2 mbk_sig533 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4907 mbk_sig533 heart_block5_na3 mbk_sig534 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4908 mbk_sig534 heart_a_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M4909 vssi heart_a_3 heart_block5_na3 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4910 vssi mbk_sig528 heart_block5_a14 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4911 mbk_sig528 heart_block5_na1 mbk_sig530 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4912 mbk_sig530 heart_a_2 mbk_sig531 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4913 mbk_sig531 heart_a_3 mbk_sig532 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4914 mbk_sig532 heart_a_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M4915 mbk_sig523 heart_block5_oa443s vssi vsse TN L=0.18U W=4.32U AS=1.5552P 
+ AD=1.5552P PS=9.36U PD=9.36U 
M4916 mbk_sig527 heart_block5_oa433s mbk_sig523 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4917 mbk_sig526 heart_block5_oa423s mbk_sig527 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4918 heart_ra_3 heart_block5_oa413s mbk_sig526 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M4919 mbk_sig522 heart_block5_s312 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4920 heart_block5_a312s heart_block5_a12 mbk_sig522 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4921 vssi mbk_sig517 heart_block5_oa423s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4922 mbk_sig517 heart_block5_a310s mbk_sig518 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4923 mbk_sig518 heart_block5_a311s mbk_sig519 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4924 mbk_sig519 heart_block5_a312s mbk_sig520 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4925 mbk_sig520 heart_block5_a39s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4926 mbk_sig515 heart_block5_s39 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4927 heart_block5_a39s heart_block5_a9 mbk_sig515 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4928 vssi mbk_sig514 heart_block5_a11 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4929 mbk_sig514 heart_a_1 mbk_sig511 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4930 mbk_sig511 heart_block5_na2 mbk_sig512 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4931 mbk_sig512 heart_a_3 mbk_sig513 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4932 mbk_sig513 heart_block5_na0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4933 mbk_sig508 heart_block5_s212 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4934 heart_block5_b212s heart_block5_b12 mbk_sig508 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4935 vssi mbk_sig502 heart_block5_m_2_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4936 mbk_sig504 mbk_sig502 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4937 heart_block5_m_2_3_dff_s mbk_sig505 mbk_sig504 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4938 vssi mbk_sig507 heart_block5_m_2_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4939 vssi heart_block5_m_2_3_dff_m mbk_sig502 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4940 heart_block5_m_2_3_dff_m heart_block5_ck2 mbk_sig501 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4941 mbk_sig505 heart_block5_ck2 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4942 vssi heart_block5_m_2_3_dff_s mbk_sig507 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4943 heart_block5_s32 heart_block5_m_2_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M4944 mbk_sig501 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4945 mbk_sig465 heart_block1_ssa0 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4946 vssi heart_block1_ssd0 mbk_sig465 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4947 vssi mbk_sig465 heart_r_0 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4948 vssi heart_block2_selray heart_block2_selaluy vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4949 mbk_sig463 heart_block2_syra1 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4950 vssi heart_block2_syalu1 mbk_sig463 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4951 vssi mbk_sig463 yc_1 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4952 vssi mbk_sig461 heart_block2_syra1 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4953 mbk_sig461 heart_ra_1 mbk_sig462 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4954 mbk_sig462 heart_block2_selray vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4955 vssi mbk_sig458 heart_block2_syalu1 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4956 mbk_sig458 heart_block2_a26ms_i0 mbk_sig457 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4957 mbk_sig457 heart_block2_selaluy vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4958 vssi mbk_sig455 heart_block1_ssa0 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4959 mbk_sig455 heart_ra_0 mbk_sig454 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4960 mbk_sig454 heart_block1_selar vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4961 vssi mbk_sig453 heart_block5_enable vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4962 mbk_sig453 cko mbk_sig452 vsse TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
M4963 mbk_sig452 heart_block5_wram vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M4964 vssi mbk_sig450 heart_block1_sra1 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4965 mbk_sig450 heart_ra_1 mbk_sig451 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4966 mbk_sig451 heart_block1_selas vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4967 vssi mbk_sig446 heart_block5_wram vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4968 mbk_sig446 heart_fonc_mode mbk_sig448 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4969 mbk_sig448 heart_block5_o21s vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4970 mbk_sig443 heart_r_2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4971 vssi heart_block3_n0 mbk_sig443 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4972 mbk_sig445 heart_block3_n0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4973 heart_block3_x02 heart_r_2 mbk_sig445 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M4974 vssi mbk_sig443 heart_block3_x02 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4975 vssi mbk_sig440 heart_block1_sra3 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4976 mbk_sig440 heart_ra_3 mbk_sig441 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4977 mbk_sig441 heart_block1_selas vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4978 mbk_sig437 ii_8 vssi vsse TN L=0.18U W=0.72U AS=0.2592P AD=0.2592P 
+ PS=2.16U PD=2.16U 
M4979 vssi ii_7 mbk_sig437 vsse TN L=0.18U W=0.72U AS=0.2592P AD=0.2592P 
+ PS=2.16U PD=2.16U 
M4980 vssi mbk_sig437 heart_block5_o21s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4981 vssi mbk_sig436 heart_block1_srq2 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4982 mbk_sig436 heart_q_2 mbk_sig438 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4983 mbk_sig438 heart_block1_selqs vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4984 vssi mbk_sig433 heart_block1_ssa3 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4985 mbk_sig433 heart_ra_3 mbk_sig434 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4986 mbk_sig434 heart_block1_selar vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4987 vssi mbk_sig430 heart_s_2 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4988 mbk_sig430 heart_block1_srq2 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4989 vssi heart_block1_sra2 mbk_sig430 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4990 mbk_sig430 heart_block1_srb2 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M4991 vssi mbk_sig428 heart_block1_sra2 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4992 mbk_sig428 heart_ra_2 mbk_sig431 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4993 mbk_sig431 heart_block1_selas vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M4994 vssi mbk_sig424 heart_block5_m_13_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4995 mbk_sig422 mbk_sig424 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M4996 heart_block5_m_13_3_dff_s mbk_sig423 mbk_sig422 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M4997 vssi mbk_sig426 heart_block5_m_13_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M4998 vssi heart_block5_m_13_3_dff_m mbk_sig424 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M4999 heart_block5_m_13_3_dff_m heart_block5_ck13 mbk_sig419 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5000 mbk_sig423 heart_block5_ck13 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M5001 vssi heart_block5_m_13_3_dff_s mbk_sig426 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5002 heart_block5_s313 heart_block5_m_13_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5003 mbk_sig419 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5004 vssi mbk_sig416 heart_block4_test_mode vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5005 mbk_sig416 testi mbk_sig420 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5006 mbk_sig420 heart_block4_n14s vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5007 vssi testi heart_block4_n15s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5008 vssi mbk_sig405 heart_block5_m_16_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5009 mbk_sig410 mbk_sig405 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5010 heart_block5_m_16_0_dff_s mbk_sig412 mbk_sig410 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5011 vssi mbk_sig411 heart_block5_m_16_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5012 vssi heart_block5_m_16_0_dff_m mbk_sig405 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5013 heart_block5_m_16_0_dff_m heart_block5_ck16 mbk_sig407 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5014 mbk_sig412 heart_block5_ck16 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M5015 vssi heart_block5_m_16_0_dff_s mbk_sig411 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5016 heart_block5_s016 heart_block5_m_16_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5017 mbk_sig407 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5018 mbk_sig402 heart_block5_s016 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5019 heart_block5_b016s heart_block5_b16 mbk_sig402 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5020 mbk_sig403 heart_block5_s116 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5021 heart_block5_a116s heart_block5_a16 mbk_sig403 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5022 mbk_sig397 heart_block5_s016 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5023 heart_block5_a016s heart_block5_a16 mbk_sig397 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5024 vssi mbk_sig396 heart_block5_oa411s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5025 mbk_sig396 heart_block5_a114s mbk_sig392 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5026 mbk_sig392 heart_block5_a115s mbk_sig390 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5027 mbk_sig390 heart_block5_a116s mbk_sig391 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5028 mbk_sig391 heart_block5_a113s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5029 vssi mbk_sig383 heart_block5_m_14_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5030 mbk_sig387 mbk_sig383 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5031 heart_block5_m_14_2_dff_s mbk_sig385 mbk_sig387 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5032 vssi mbk_sig388 heart_block5_m_14_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5033 vssi heart_block5_m_14_2_dff_m mbk_sig383 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5034 heart_block5_m_14_2_dff_m heart_block5_ck14 mbk_sig382 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5035 mbk_sig385 heart_block5_ck14 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M5036 vssi heart_block5_m_14_2_dff_s mbk_sig388 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5037 heart_block5_s214 heart_block5_m_14_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5038 mbk_sig382 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5039 vssi mbk_sig381 heart_block5_ck14 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5040 mbk_sig381 heart_block5_enable mbk_sig380 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5041 mbk_sig380 heart_block5_b14 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5042 mbk_sig377 heart_block5_s314 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5043 heart_block5_a314s heart_block5_a14 mbk_sig377 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5044 vssi mbk_sig375 heart_block5_m_9_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5045 mbk_sig373 mbk_sig375 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5046 heart_block5_m_9_0_dff_s mbk_sig374 mbk_sig373 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5047 vssi mbk_sig378 heart_block5_m_9_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5048 vssi heart_block5_m_9_0_dff_m mbk_sig375 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5049 heart_block5_m_9_0_dff_m heart_block5_ck9 mbk_sig370 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5050 mbk_sig374 heart_block5_ck9 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M5051 vssi heart_block5_m_9_0_dff_s mbk_sig378 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5052 heart_block5_s09 heart_block5_m_9_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5053 mbk_sig370 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5054 vssi mbk_sig369 heart_block5_oa410s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5055 mbk_sig369 heart_block5_a014s mbk_sig372 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5056 mbk_sig372 heart_block5_a015s mbk_sig367 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5057 mbk_sig367 heart_block5_a016s mbk_sig366 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5058 mbk_sig366 heart_block5_a013s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5059 mbk_sig363 heart_block5_s114 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5060 heart_block5_a114s heart_block5_a14 mbk_sig363 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5061 vssi heart_a_2 heart_block5_na2 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5062 vssi mbk_sig356 heart_block5_m_9_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5063 mbk_sig361 mbk_sig356 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5064 heart_block5_m_9_1_dff_s mbk_sig358 mbk_sig361 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5065 vssi mbk_sig362 heart_block5_m_9_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5066 vssi heart_block5_m_9_1_dff_m mbk_sig356 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5067 heart_block5_m_9_1_dff_m heart_block5_ck9 mbk_sig355 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5068 mbk_sig358 heart_block5_ck9 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M5069 vssi heart_block5_m_9_1_dff_s mbk_sig362 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5070 heart_block5_s19 heart_block5_m_9_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5071 mbk_sig355 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5072 mbk_sig353 heart_block5_s09 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5073 heart_block5_b09s heart_block5_b9 mbk_sig353 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5074 mbk_sig349 heart_block5_s215 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5075 heart_block5_a215s heart_block5_a15 mbk_sig349 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5076 mbk_sig350 heart_block5_s19 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5077 heart_block5_b19s heart_block5_b9 mbk_sig350 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5078 vssi mbk_sig343 heart_block5_m_11_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5079 mbk_sig347 mbk_sig343 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5080 heart_block5_m_11_1_dff_s mbk_sig345 mbk_sig347 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5081 vssi mbk_sig348 heart_block5_m_11_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5082 vssi heart_block5_m_11_1_dff_m mbk_sig343 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5083 heart_block5_m_11_1_dff_m heart_block5_ck11 mbk_sig342 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5084 mbk_sig345 heart_block5_ck11 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M5085 vssi heart_block5_m_11_1_dff_s mbk_sig348 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5086 heart_block5_s111 heart_block5_m_11_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5087 mbk_sig342 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5088 vssi mbk_sig338 heart_block5_ob421s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5089 mbk_sig338 heart_block5_b110s mbk_sig339 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5090 mbk_sig339 heart_block5_b111s mbk_sig340 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5091 mbk_sig340 heart_block5_b112s mbk_sig341 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5092 mbk_sig341 heart_block5_b19s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5093 vssi mbk_sig332 heart_block5_a15 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5094 mbk_sig332 heart_a_1 mbk_sig335 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5095 mbk_sig335 heart_a_2 mbk_sig334 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5096 mbk_sig334 heart_a_3 mbk_sig336 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5097 mbk_sig336 heart_block5_na0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5098 mbk_sig330 heart_block5_s211 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5099 heart_block5_a211s heart_block5_a11 mbk_sig330 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5100 vssi mbk_sig326 heart_block5_a9 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5101 mbk_sig326 heart_block5_na1 mbk_sig324 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5102 mbk_sig324 heart_block5_na2 mbk_sig325 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5103 mbk_sig325 heart_a_3 mbk_sig327 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5104 mbk_sig327 heart_block5_na0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5105 mbk_sig323 heart_block5_s011 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5106 heart_block5_a011s heart_block5_a11 mbk_sig323 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5107 vssi mbk_sig321 heart_block5_oa420s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5108 mbk_sig321 heart_block5_a010s mbk_sig320 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5109 mbk_sig320 heart_block5_a011s mbk_sig318 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5110 mbk_sig318 heart_block5_a012s mbk_sig319 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5111 mbk_sig319 heart_block5_a09s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5112 mbk_sig315 heart_block5_s19 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5113 heart_block5_a19s heart_block5_a9 mbk_sig315 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5114 mbk_sig316 heart_block5_s09 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5115 heart_block5_a09s heart_block5_a9 mbk_sig316 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5116 vssi mbk_sig309 heart_block5_a12 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5117 mbk_sig309 heart_a_1 mbk_sig307 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5118 mbk_sig307 heart_block5_na2 mbk_sig308 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5119 mbk_sig308 heart_a_3 mbk_sig310 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5120 mbk_sig310 heart_a_0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
M5121 vssi mbk_sig303 heart_block5_oa421s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5122 mbk_sig303 heart_block5_a110s mbk_sig304 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5123 mbk_sig304 heart_block5_a111s mbk_sig305 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5124 mbk_sig305 heart_block5_a112s mbk_sig306 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5125 mbk_sig306 heart_block5_a19s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5126 vssi mbk_sig299 heart_block5_m_12_2_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5127 mbk_sig297 mbk_sig299 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5128 heart_block5_m_12_2_dff_s mbk_sig298 mbk_sig297 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5129 vssi mbk_sig302 heart_block5_m_12_2_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5130 vssi heart_block5_m_12_2_dff_m mbk_sig299 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5131 heart_block5_m_12_2_dff_m heart_block5_ck12 mbk_sig293 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5132 mbk_sig298 heart_block5_ck12 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M5133 vssi heart_block5_m_12_2_dff_s mbk_sig302 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5134 heart_block5_s212 heart_block5_m_12_2_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5135 mbk_sig293 heart_block5_shram2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5136 mbk_sig294 heart_block5_s310 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5137 heart_block5_a310s heart_block5_a10 mbk_sig294 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5138 mbk_sig289 heart_block5_s110 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5139 heart_block5_b110s heart_block5_b10 mbk_sig289 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5140 mbk_sig286 heart_block5_s012 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5141 heart_block5_a012s heart_block5_a12 mbk_sig286 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5142 mbk_sig285 heart_block5_s110 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5143 heart_block5_a110s heart_block5_a10 mbk_sig285 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5144 vssi mbk_sig264 heart_block1_ssd0 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5145 mbk_sig264 heart_d_0 mbk_sig263 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5146 mbk_sig263 heart_block1_seldr vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5147 vssi ii_2 heart_block1_ni2 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5148 vssi mbk_sig262 heart_block1_selas vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5149 mbk_sig262 heart_block1_ni1 mbk_sig260 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5150 mbk_sig260 ii_2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5151 vssi mbk_sig259 heart_block1_selar vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5152 mbk_sig259 heart_block1_ni2 mbk_sig261 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5153 mbk_sig261 heart_block1_ni1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5154 vssi ii_1 heart_block1_ni1 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5155 mbk_sig257 heart_block1_ssa3 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M5156 vssi heart_block1_ssd3 mbk_sig257 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M5157 vssi mbk_sig257 heart_r_3 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5158 vssi mbk_sig256 heart_block1_seldr vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5159 mbk_sig256 heart_block1_o22s mbk_sig255 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5160 mbk_sig255 ii_2 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5161 vssi mbk_sig254 heart_block1_ssd2 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5162 mbk_sig254 heart_d_2 mbk_sig253 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5163 mbk_sig253 heart_block1_seldr vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5164 mbk_sig251 heart_block1_ssa2 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M5165 vssi heart_block1_ssd2 mbk_sig251 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M5166 vssi mbk_sig251 heart_r_2 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5167 mbk_sig247 heart_r_1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5168 vssi heart_block3_n0 mbk_sig247 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5169 mbk_sig249 heart_block3_n0 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5170 heart_block3_x01 heart_r_1 mbk_sig249 vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5171 vssi mbk_sig247 heart_block3_x01 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5172 mbk_sig244 ii_1 vssi vsse TN L=0.18U W=0.72U AS=0.2592P AD=0.2592P 
+ PS=2.16U PD=2.16U 
M5173 vssi ii_0 mbk_sig244 vsse TN L=0.18U W=0.72U AS=0.2592P AD=0.2592P 
+ PS=2.16U PD=2.16U 
M5174 vssi mbk_sig244 heart_block1_o22s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5175 vssi mbk_sig243 heart_block2_syra2 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5176 mbk_sig243 heart_ra_2 mbk_sig245 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5177 mbk_sig245 heart_block2_selray vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5178 mbk_sig241 heart_block2_syra2 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M5179 vssi heart_block2_syalu2 mbk_sig241 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M5180 vssi mbk_sig241 yc_2 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5181 mbk_sig239 ii_1 vssi vsse TN L=0.18U W=0.72U AS=0.2592P AD=0.2592P 
+ PS=2.16U PD=2.16U 
M5182 vssi heart_block1_ni2 mbk_sig239 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M5183 vssi mbk_sig239 heart_block1_o21s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5184 vssi mbk_sig238 heart_block1_ssa2 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5185 mbk_sig238 heart_ra_2 mbk_sig237 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5186 mbk_sig237 heart_block1_selar vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5187 vssi mbk_sig236 heart_block1_ssd3 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5188 mbk_sig236 heart_d_3 mbk_sig235 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5189 mbk_sig235 heart_block1_seldr vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5190 vssi ii_6 heart_block2_ni6 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5191 mbk_sig232 ii_7 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5192 mbk_sig233 heart_block2_ni6 mbk_sig232 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5193 mbk_sig234 heart_block2_ni8 mbk_sig233 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5194 vssi mbk_sig234 heart_block2_selray vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5195 vssi ii_8 heart_block2_ni8 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5196 vssi mbk_sig230 heart_block1_ssa1 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5197 mbk_sig230 heart_ra_1 mbk_sig231 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5198 mbk_sig231 heart_block1_selar vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5199 mbk_sig228 heart_block1_ssa1 vssi vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M5200 vssi heart_block1_ssd1 mbk_sig228 vsse TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
M5201 vssi mbk_sig228 heart_r_1 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5202 vssi mbk_sig227 heart_block1_ssd1 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5203 mbk_sig227 heart_d_1 mbk_sig226 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5204 mbk_sig226 heart_block1_seldr vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5205 vssi mbk_sig224 heart_block1_selqs vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5206 mbk_sig224 heart_block1_o21s mbk_sig225 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5207 mbk_sig225 heart_block1_ni0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5208 vssi ii_0 heart_block1_ni0 vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5209 vssi mbk_sig223 heart_block1_selbs vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5210 mbk_sig223 heart_block1_ni2 mbk_sig221 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5211 mbk_sig221 ii_0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5212 mbk_sig222 heart_block5_s014 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5213 heart_block5_a014s heart_block5_a14 mbk_sig222 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5214 mbk_sig220 heart_block5_s014 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5215 heart_block5_b014s heart_block5_b14 mbk_sig220 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5216 vssi mbk_sig147 heart_block5_m_14_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5217 mbk_sig218 mbk_sig147 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5218 heart_block5_m_14_0_dff_s mbk_sig219 mbk_sig218 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5219 vssi mbk_sig149 heart_block5_m_14_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5220 vssi heart_block5_m_14_0_dff_m mbk_sig147 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5221 heart_block5_m_14_0_dff_m heart_block5_ck14 mbk_sig217 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5222 mbk_sig219 heart_block5_ck14 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M5223 vssi heart_block5_m_14_0_dff_s mbk_sig149 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5224 heart_block5_s014 heart_block5_m_14_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5225 mbk_sig217 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5226 vssi mbk_sig143 heart_block5_m_14_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5227 mbk_sig216 mbk_sig143 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5228 heart_block5_m_14_1_dff_s mbk_sig215 mbk_sig216 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5229 vssi mbk_sig145 heart_block5_m_14_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5230 vssi heart_block5_m_14_1_dff_m mbk_sig143 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5231 heart_block5_m_14_1_dff_m heart_block5_ck14 mbk_sig214 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5232 mbk_sig215 heart_block5_ck14 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M5233 vssi heart_block5_m_14_1_dff_s mbk_sig145 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5234 heart_block5_s114 heart_block5_m_14_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5235 mbk_sig214 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5236 mbk_sig213 heart_block5_s015 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5237 heart_block5_b015s heart_block5_b15 mbk_sig213 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5238 mbk_sig212 heart_block5_s314 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5239 heart_block5_b314s heart_block5_b14 mbk_sig212 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5240 mbk_sig211 heart_block5_s015 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5241 heart_block5_a015s heart_block5_a15 mbk_sig211 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5242 mbk_sig131 heart_block5_oa442s vssi vsse TN L=0.18U W=4.32U AS=1.5552P 
+ AD=1.5552P PS=9.36U PD=9.36U 
M5243 mbk_sig130 heart_block5_oa432s mbk_sig131 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M5244 mbk_sig132 heart_block5_oa422s mbk_sig130 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M5245 heart_ra_2 heart_block5_oa412s mbk_sig132 vsse TN L=0.18U W=4.32U 
+ AS=1.5552P AD=1.5552P PS=9.36U PD=9.36U 
M5246 vssi mbk_sig125 heart_block5_m_14_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5247 mbk_sig210 mbk_sig125 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5248 heart_block5_m_14_3_dff_s mbk_sig209 mbk_sig210 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5249 vssi mbk_sig128 heart_block5_m_14_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5250 vssi heart_block5_m_14_3_dff_m mbk_sig125 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5251 heart_block5_m_14_3_dff_m heart_block5_ck14 mbk_sig208 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5252 mbk_sig209 heart_block5_ck14 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M5253 vssi heart_block5_m_14_3_dff_s mbk_sig128 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5254 heart_block5_s314 heart_block5_m_14_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5255 mbk_sig208 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5256 mbk_sig207 heart_block5_s011 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5257 heart_block5_b011s heart_block5_b11 mbk_sig207 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5258 mbk_sig206 heart_block5_s114 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5259 heart_block5_b114s heart_block5_b14 mbk_sig206 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5260 vssi mbk_sig115 heart_block5_m_15_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5261 mbk_sig204 mbk_sig115 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5262 heart_block5_m_15_0_dff_s mbk_sig205 mbk_sig204 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5263 vssi mbk_sig119 heart_block5_m_15_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5264 vssi heart_block5_m_15_0_dff_m mbk_sig115 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5265 heart_block5_m_15_0_dff_m heart_block5_ck15 mbk_sig203 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5266 mbk_sig205 heart_block5_ck15 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M5267 vssi heart_block5_m_15_0_dff_s mbk_sig119 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5268 heart_block5_s015 heart_block5_m_15_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5269 mbk_sig203 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5270 vssi mbk_sig110 heart_block5_m_11_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5271 mbk_sig201 mbk_sig110 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5272 heart_block5_m_11_0_dff_s mbk_sig202 mbk_sig201 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5273 vssi mbk_sig113 heart_block5_m_11_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5274 vssi heart_block5_m_11_0_dff_m mbk_sig110 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5275 heart_block5_m_11_0_dff_m heart_block5_ck11 mbk_sig200 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5276 mbk_sig202 heart_block5_ck11 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M5277 vssi heart_block5_m_11_0_dff_s mbk_sig113 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5278 heart_block5_s011 heart_block5_m_11_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5279 mbk_sig200 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5280 mbk_sig199 heart_block5_s111 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5281 heart_block5_b111s heart_block5_b11 mbk_sig199 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5282 vssi mbk_sig105 heart_block5_ob420s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5283 mbk_sig105 heart_block5_b010s mbk_sig104 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5284 mbk_sig104 heart_block5_b011s mbk_sig99 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5285 mbk_sig99 heart_block5_b012s mbk_sig98 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5286 mbk_sig98 heart_block5_b09s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5287 vssi mbk_sig94 heart_block5_m_12_3_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5288 mbk_sig197 mbk_sig94 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5289 heart_block5_m_12_3_dff_s mbk_sig198 mbk_sig197 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5290 vssi mbk_sig97 heart_block5_m_12_3_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5291 vssi heart_block5_m_12_3_dff_m mbk_sig94 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5292 heart_block5_m_12_3_dff_m heart_block5_ck12 mbk_sig196 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5293 mbk_sig198 heart_block5_ck12 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M5294 vssi heart_block5_m_12_3_dff_s mbk_sig97 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5295 heart_block5_s312 heart_block5_m_12_3_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5296 mbk_sig196 heart_block5_shram3 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5297 vssi mbk_sig88 heart_block5_oa422s vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5298 mbk_sig88 heart_block5_a210s mbk_sig87 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5299 mbk_sig87 heart_block5_a211s mbk_sig89 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5300 mbk_sig89 heart_block5_a212s mbk_sig90 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5301 mbk_sig90 heart_block5_a29s vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5302 mbk_sig195 heart_block5_s29 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5303 heart_block5_a29s heart_block5_a9 mbk_sig195 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5304 vssi mbk_sig79 heart_block5_m_12_0_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5305 mbk_sig193 mbk_sig79 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5306 heart_block5_m_12_0_dff_s mbk_sig194 mbk_sig193 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5307 vssi mbk_sig82 heart_block5_m_12_0_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5308 vssi heart_block5_m_12_0_dff_m mbk_sig79 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5309 heart_block5_m_12_0_dff_m heart_block5_ck12 mbk_sig192 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5310 mbk_sig194 heart_block5_ck12 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M5311 vssi heart_block5_m_12_0_dff_s mbk_sig82 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5312 heart_block5_s012 heart_block5_m_12_0_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5313 mbk_sig192 heart_block5_shram0 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5314 mbk_sig190 heart_block5_s012 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5315 heart_block5_b012s heart_block5_b12 mbk_sig190 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5316 mbk_sig191 heart_block5_s111 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5317 heart_block5_a111s heart_block5_a11 mbk_sig191 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5318 mbk_sig188 heart_block5_s112 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5319 heart_block5_a112s heart_block5_a12 mbk_sig188 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5320 mbk_sig189 heart_block5_s112 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5321 heart_block5_b112s heart_block5_b12 mbk_sig189 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5322 vssi mbk_sig67 heart_block5_m_12_1_dff_m vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5323 mbk_sig186 mbk_sig67 vssi vsse TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
M5324 heart_block5_m_12_1_dff_s mbk_sig187 mbk_sig186 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5325 vssi mbk_sig69 heart_block5_m_12_1_dff_s vsse TN L=1.26U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
M5326 vssi heart_block5_m_12_1_dff_m mbk_sig67 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5327 heart_block5_m_12_1_dff_m heart_block5_ck12 mbk_sig184 vsse TN L=0.18U 
+ W=1.08U AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5328 mbk_sig187 heart_block5_ck12 vssi vsse TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
M5329 vssi heart_block5_m_12_1_dff_s mbk_sig69 vsse TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
M5330 heart_block5_s112 heart_block5_m_12_1_dff_s vssi vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
M5331 mbk_sig184 heart_block5_shram1 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5332 vssi mbk_sig183 heart_block5_ck12 vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5333 mbk_sig183 heart_block5_enable mbk_sig185 vsse TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
M5334 mbk_sig185 heart_block5_b12 vssi vsse TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
M5335 mbk_sig182 heart_block5_s212 vssi vsse TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
M5336 heart_block5_a212s heart_block5_a12 mbk_sig182 vsse TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
C0 zero vsse 1.80526e-13

C1 y_3 vsse 1.80958e-13

C2 y_2 vsse 1.80958e-13

C3 y_1 vsse 1.80958e-13

C4 y_0 vsse 1.80959e-13

C5 vssi vsse 2.37451e-12

C6 mbk_sig1970 vsse 1.33164e-16
C7 mbk_sig1964 vsse 1.33164e-16
C8 mbk_sig1807 vsse 1.33164e-16
C9 mbk_sig1801 vsse 3.68064e-16
C10 mbk_sig1629 vsse 1.33164e-16
C11 mbk_sig1625 vsse 1.33164e-16
C12 mbk_sig1617 vsse 1.33164e-16
C13 mbk_sig1605 vsse 3.68064e-16
C14 mbk_sig1433 vsse 1.33164e-16
C15 mbk_sig1412 vsse 3.68064e-16
C16 mbk_sig1392 vsse 3.68064e-16
C17 mbk_sig1233 vsse 1.33164e-16
C18 mbk_sig1062 vsse 1.33164e-16
C19 mbk_sig1060 vsse 1.33164e-16
C20 mbk_sig868 vsse 1.33164e-16
C21 mbk_sig855 vsse 1.33164e-16
C22 mbk_sig839 vsse 1.33164e-16
C23 mbk_sig679 vsse 1.33164e-16
C24 mbk_sig674 vsse 1.33164e-16
C25 mbk_sig474 vsse 1.33164e-16
C26 mbk_sig250 vsse 1.33164e-16
C27 mbk_sig55 vsse 1.57322e-14
C28 mbk_sig178 vsse 2.19348e-15
C29 mbk_sig179 vsse 1.7321e-15
C30 mbk_sig467 vsse 1.57322e-14
C31 mbk_sig478 vsse 2.19348e-15
C32 mbk_sig479 vsse 1.7321e-15
C33 mbk_sig682 vsse 1.57322e-14
C34 mbk_sig687 vsse 2.19348e-15
C35 mbk_sig686 vsse 1.7321e-15
C36 mbk_sig871 vsse 1.57322e-14
C37 mbk_sig878 vsse 2.19348e-15
C38 mbk_sig879 vsse 1.7321e-15
C39 mbk_sig1066 vsse 3.23806e-15
C40 mbk_sig1271 vsse 3.23806e-15
C41 mbk_sig1466 vsse 3.23806e-15
C42 mbk_sig1636 vsse 2.06712e-15
C43 mbk_sig1647 vsse 1.7321e-15
C44 mbk_sig1646 vsse 2.19348e-15
C45 mbk_sig1639 vsse 1.33446e-14
C46 mbk_sig1638 vsse 1.19673e-14
C47 mbk_sig1653 vsse 2.04962e-15
C48 mbk_sig1652 vsse 2.4394e-15
C49 mbk_sig1815 vsse 2.06712e-15
C50 mbk_sig1827 vsse 1.7321e-15
C51 mbk_sig1826 vsse 2.19348e-15
C52 mbk_sig1818 vsse 1.33446e-14
C53 mbk_sig1817 vsse 1.19673e-14
C54 mbk_sig1836 vsse 2.04962e-15
C55 mbk_sig1835 vsse 2.4394e-15
C56 mbk_sig44 vsse 3.23806e-15
C57 mbk_sig57 vsse 1.57322e-14
C58 mbk_sig265 vsse 2.19348e-15
C59 mbk_sig180 vsse 1.7321e-15
C60 mbk_sig469 vsse 1.57322e-14
C61 mbk_sig480 vsse 2.19348e-15
C62 mbk_sig481 vsse 1.7321e-15
C63 mbk_sig671 vsse 2.06712e-15
C64 mbk_sig683 vsse 1.7321e-15
C65 mbk_sig688 vsse 2.19348e-15
C66 mbk_sig669 vsse 1.33446e-14
C67 mbk_sig670 vsse 1.19673e-14
C68 mbk_sig689 vsse 2.04962e-15
C69 mbk_sig690 vsse 2.4394e-15
C70 mbk_sig876 vsse 2.06712e-15
C71 mbk_sig881 vsse 1.7321e-15
C72 mbk_sig880 vsse 2.19348e-15
C73 mbk_sig873 vsse 1.33446e-14
C74 mbk_sig874 vsse 1.19673e-14
C75 mbk_sig884 vsse 2.04962e-15
C76 mbk_sig885 vsse 2.4394e-15
C77 mbk_sig1223 vsse 2.04962e-15
C78 mbk_sig1076 vsse 1.19673e-14
C79 mbk_sig1084 vsse 2.19348e-15
C80 mbk_sig1224 vsse 2.4394e-15
C81 mbk_sig1075 vsse 1.33704e-14
C82 mbk_sig1085 vsse 1.7321e-15
C83 mbk_sig1260 vsse 2.04962e-15
C84 mbk_sig1248 vsse 1.19673e-14
C85 mbk_sig1251 vsse 2.19348e-15
C86 mbk_sig1261 vsse 2.4394e-15
C87 mbk_sig1247 vsse 1.33704e-14
C88 mbk_sig1250 vsse 1.7321e-15
C89 mbk_sig1458 vsse 2.04962e-15
C90 mbk_sig1449 vsse 1.19673e-14
C91 mbk_sig1454 vsse 2.19348e-15
C92 mbk_sig1459 vsse 2.4394e-15
C93 mbk_sig1448 vsse 1.33704e-14
C94 mbk_sig1450 vsse 1.7321e-15
C95 mbk_sig1640 vsse 2.04962e-15
C96 mbk_sig1633 vsse 1.19673e-14
C97 mbk_sig1634 vsse 2.19348e-15
C98 mbk_sig1641 vsse 2.4394e-15
C99 mbk_sig1632 vsse 1.33704e-14
C100 mbk_sig1635 vsse 1.7321e-15
C101 mbk_sig1975 vsse 3.23806e-15
C102 mbk_sig13 vsse 1.57322e-14
C103 mbk_sig16 vsse 2.19348e-15
C104 mbk_sig17 vsse 1.7321e-15
C105 mbk_sig20 vsse 3.23806e-15
C106 mbk_sig22 vsse 3.23806e-15
C107 mbk_sig24 vsse 3.23806e-15
C108 mbk_sig40 vsse 2.14942e-15
C109 mbk_sig26 vsse 3.23806e-15
C110 mbk_sig28 vsse 3.23806e-15
C111 mbk_sig30 vsse 3.23806e-15
C112 mbk_sig32 vsse 3.23806e-15
C113 mbk_sig34 vsse 3.23806e-15
C114 mbk_sig36 vsse 3.23806e-15
C115 ck_log_log_ck vsse 1.49339e-13
C116 mbk_sig38 vsse 9.29916e-15
C117 mbk_sig1976 vsse 3.23806e-15
C118 mbk_sig1977 vsse 3.23806e-15
C119 mbk_sig1978 vsse 3.23806e-15
C120 mbk_sig1979 vsse 3.23806e-15
C121 mbk_sig1980 vsse 3.23806e-15
C122 mbk_sig1981 vsse 3.23806e-15
C123 mbk_sig1982 vsse 3.23806e-15
C124 mbk_sig1983 vsse 3.23806e-15
C125 mbk_sig1984 vsse 3.23806e-15
C126 mbk_sig1985 vsse 3.23806e-15
C127 mbk_sig1986 vsse 3.23806e-15
C128 mbk_sig1987 vsse 3.23806e-15
C129 heart_block3_no31 vsse 2.51748e-15
C130 mbk_sig1967 vsse 7.91856e-16
C131 heart_block3_no21 vsse 2.46046e-15
C132 mbk_sig1965 vsse 5.68296e-16
C133 heart_block3_x21 vsse 3.44639e-15
C134 mbk_sig1961 vsse 7.91856e-16
C135 mbk_sig1959 vsse 6.57072e-16
C136 decalgc vsse 5.88044e-15
C137 mbk_sig1958 vsse 5.51448e-16
C138 heart_block4_a29s vsse 3.23741e-15
C139 mbk_sig1955 vsse 5.51448e-16
C140 heart_block3_fb1 vsse 4.06134e-15
C141 mbk_sig1953 vsse 5.51448e-16
C142 mbk_sig1952 vsse 5.51448e-16
C143 mbk_sig1949 vsse 5.51448e-16
C144 heart_block4_a221s vsse 3.56011e-15
C145 heart_block4_a219s vsse 2.50873e-15
C146 mbk_sig1946 vsse 7.12152e-16
C147 heart_block4_a220s vsse 2.76372e-15
C148 mbk_sig1945 vsse 5.51448e-16
C149 heart_block4_a28s vsse 3.45708e-15
C150 heart_block4_a212s vsse 3.39941e-15
C151 mbk_sig1942 vsse 5.68296e-16
C152 mbk_sig1940 vsse 5.51448e-16
C153 q0i vsse 1.03542e-14
C154 mbk_sig1939 vsse 5.51448e-16
C155 mbk_sig1936 vsse 5.51448e-16
C156 f3c vsse 8.93349e-15
C157 mbk_sig1935 vsse 5.51448e-16
C158 heart_block4_insh1 vsse 7.6532e-15
C159 mbk_sig1933 vsse 5.51448e-16
C160 mbk_sig1929 vsse 3.00996e-16
C161 mbk_sig1925 vsse 1.35108e-15
C162 heart_block5_m_1_2_dff_m vsse 5.32008e-16
C163 mbk_sig1930 vsse 6.73272e-16
C164 mbk_sig1931 vsse 7.51032e-16
C165 heart_block5_m_1_2_dff_s vsse 5.89032e-16
C166 mbk_sig1927 vsse 2.26476e-16
C167 heart_block4_a227s vsse 2.98469e-15
C168 heart_block4_a225s vsse 2.88976e-15
C169 mbk_sig1922 vsse 7.12152e-16
C170 mbk_sig1921 vsse 5.51448e-16
C171 mbk_sig1919 vsse 7.75008e-16
C172 mbk_sig1914 vsse 7.75008e-16
C173 heart_block4_a226s vsse 2.6568e-15
C174 mbk_sig1911 vsse 5.51448e-16
C175 mbk_sig1909 vsse 7.75008e-16
C176 mbk_sig1905 vsse 7.75008e-16
C177 mbk_sig1900 vsse 7.75008e-16
C178 mbk_sig1894 vsse 7.75008e-16
C179 mbk_sig1890 vsse 7.75008e-16
C180 mbk_sig1887 vsse 3.00996e-16
C181 mbk_sig1883 vsse 1.35108e-15
C182 heart_block5_m_8_1_dff_m vsse 5.32008e-16
C183 mbk_sig1885 vsse 6.73272e-16
C184 mbk_sig1888 vsse 7.51032e-16
C185 heart_block5_m_8_1_dff_s vsse 5.89032e-16
C186 mbk_sig1881 vsse 2.26476e-16
C187 heart_block5_s18 vsse 3.84232e-15
C188 mbk_sig1880 vsse 7.75008e-16
C189 mbk_sig1876 vsse 5.51448e-16
C190 mbk_sig1874 vsse 5.51448e-16
C191 mbk_sig1870 vsse 3.00996e-16
C192 mbk_sig1866 vsse 1.35108e-15
C193 heart_block5_m_8_2_dff_m vsse 5.32008e-16
C194 mbk_sig1872 vsse 6.73272e-16
C195 mbk_sig1871 vsse 7.51032e-16
C196 heart_block5_m_8_2_dff_s vsse 5.89032e-16
C197 mbk_sig1868 vsse 2.26476e-16
C198 mbk_sig1862 vsse 3.00996e-16
C199 mbk_sig1857 vsse 1.35108e-15
C200 heart_block5_m_5_1_dff_m vsse 5.32008e-16
C201 mbk_sig1863 vsse 6.73272e-16
C202 mbk_sig1865 vsse 7.51032e-16
C203 heart_block5_m_5_1_dff_s vsse 5.89032e-16
C204 mbk_sig1860 vsse 2.26476e-16
C205 mbk_sig1852 vsse 3.00996e-16
C206 mbk_sig1854 vsse 1.35108e-15
C207 heart_block5_m_4_0_dff_m vsse 5.32008e-16
C208 mbk_sig1853 vsse 6.73272e-16
C209 mbk_sig1856 vsse 7.51032e-16
C210 heart_block5_m_4_0_dff_s vsse 5.89032e-16
C211 mbk_sig1851 vsse 2.26476e-16
C212 mbk_sig1848 vsse 3.00996e-16
C213 mbk_sig1844 vsse 1.35108e-15
C214 heart_block5_m_8_3_dff_m vsse 5.32008e-16
C215 mbk_sig1846 vsse 6.73272e-16
C216 mbk_sig1849 vsse 7.51032e-16
C217 heart_block5_m_8_3_dff_s vsse 5.89032e-16
C218 mbk_sig1843 vsse 2.26476e-16
C219 mbk_sig1841 vsse 5.51448e-16
C220 mbk_sig1838 vsse 5.51448e-16
C221 heart_block3_not1 vsse 1.74215e-15
C222 heart_block3_cout0 vsse 4.11577e-15
C223 heart_block3_no41 vsse 3.41366e-15
C224 heart_block3_na21 vsse 3.05078e-15
C225 heart_block4_a213s vsse 3.12725e-15
C226 mbk_sig1779 vsse 5.51448e-16
C227 heart_block3_na1_csb vsse 1.78783e-15
C228 zeroc vsse 1.36762e-14
C229 heart_block3_na0_csb vsse 2.8201e-15
C230 mbk_sig1805 vsse 7.91856e-16
C231 mbk_sig1774 vsse 5.51448e-16
C232 heart_block3_no42 vsse 3.05014e-15
C233 mbk_sig1773 vsse 5.51448e-16
C234 heart_block3_flag1 vsse 3.97548e-15
C235 mbk_sig1765 vsse 6.4476e-16
C236 mbk_sig1772 vsse 7.2414e-16
C237 heart_block4_m1_dff_s vsse 5.66676e-16
C238 mbk_sig1770 vsse 2.84472e-16
C239 mbk_sig1764 vsse 7.40988e-16
C240 mbk_sig1769 vsse 1.33164e-15
C241 heart_block4_m1_dff_m vsse 5.51124e-16
C242 mbk_sig1768 vsse 6.82992e-16
C243 heart_block4_shacc1 vsse 2.11669e-15
C244 heart_block4_a224s vsse 4.0811e-15
C245 heart_block4_a223s vsse 2.5907e-15
C246 mbk_sig1762 vsse 7.12152e-16
C247 heart_block4_a222s vsse 1.88665e-15
C248 mbk_sig1757 vsse 5.51448e-16
C249 heart_block5_a26sh vsse 3.37381e-15
C250 mbk_sig1756 vsse 7.12152e-16
C251 mbk_sig1754 vsse 5.51448e-16
C252 heart_block4_a27s vsse 1.95242e-15
C253 heart_block4_insh3 vsse 6.03061e-15
C254 mbk_sig1752 vsse 5.68296e-16
C255 mbk_sig1751 vsse 5.51448e-16
C256 mbk_sig1748 vsse 3.00996e-16
C257 mbk_sig1746 vsse 1.35108e-15
C258 heart_block5_m_1_1_dff_m vsse 5.32008e-16
C259 mbk_sig1749 vsse 6.73272e-16
C260 mbk_sig1750 vsse 7.51032e-16
C261 heart_block5_m_1_1_dff_s vsse 5.89032e-16
C262 mbk_sig1745 vsse 2.26476e-16
C263 f0c vsse 9.81509e-15
C264 mbk_sig1743 vsse 5.51448e-16
C265 mbk_sig1739 vsse 7.75008e-16
C266 mbk_sig1735 vsse 7.75008e-16
C267 heart_b_2 vsse 1.63878e-14
C268 mbk_sig1728 vsse 7.75008e-16
C269 mbk_sig1724 vsse 7.75008e-16
C270 heart_block5_b18s vsse 3.05143e-15
C271 mbk_sig1721 vsse 7.75008e-16
C272 mbk_sig1716 vsse 3.00996e-16
C273 mbk_sig1714 vsse 1.35108e-15
C274 heart_block5_m_1_0_dff_m vsse 5.32008e-16
C275 mbk_sig1717 vsse 6.73272e-16
C276 mbk_sig1718 vsse 7.51032e-16
C277 heart_block5_m_1_0_dff_s vsse 5.89032e-16
C278 mbk_sig1713 vsse 2.26476e-16
C279 heart_block5_b17s vsse 2.84602e-15
C280 mbk_sig1704 vsse 7.75008e-16
C281 heart_b_0 vsse 2.33459e-14
C282 mbk_sig1698 vsse 7.75008e-16
C283 heart_block5_nb3 vsse 1.59325e-14
C284 mbk_sig1694 vsse 3.00996e-16
C285 mbk_sig1692 vsse 1.35108e-15
C286 heart_block5_m_5_2_dff_m vsse 5.32008e-16
C287 mbk_sig1695 vsse 6.73272e-16
C288 mbk_sig1696 vsse 7.51032e-16
C289 heart_block5_m_5_2_dff_s vsse 5.89032e-16
C290 mbk_sig1691 vsse 2.26476e-16
C291 heart_block5_s38 vsse 4.55771e-15
C292 mbk_sig1685 vsse 3.00996e-16
C293 mbk_sig1683 vsse 1.35108e-15
C294 heart_block5_m_4_2_dff_m vsse 5.32008e-16
C295 mbk_sig1680 vsse 6.73272e-16
C296 mbk_sig1686 vsse 7.51032e-16
C297 heart_block5_m_4_2_dff_s vsse 5.89032e-16
C298 mbk_sig1682 vsse 2.26476e-16
C299 mbk_sig1679 vsse 5.51448e-16
C300 heart_block5_s04 vsse 3.64597e-15
C301 mbk_sig1671 vsse 3.00996e-16
C302 mbk_sig1673 vsse 1.35108e-15
C303 heart_block5_m_1_3_dff_m vsse 5.32008e-16
C304 heart_block5_ck1 vsse 1.32466e-14
C305 mbk_sig1672 vsse 6.73272e-16
C306 mbk_sig1675 vsse 7.51032e-16
C307 heart_block5_m_1_3_dff_s vsse 5.89032e-16
C308 mbk_sig1666 vsse 2.26476e-16
C309 mbk_sig1664 vsse 7.75008e-16
C310 heart_block5_b33s vsse 3.04819e-15
C311 heart_block5_b31s vsse 2.56608e-15
C312 mbk_sig1658 vsse 3.00996e-16
C313 mbk_sig1656 vsse 1.35108e-15
C314 heart_block5_m_3_3_dff_m vsse 5.32008e-16
C315 mbk_sig1659 vsse 6.73272e-16
C316 mbk_sig1660 vsse 7.51032e-16
C317 heart_block5_m_3_3_dff_s vsse 5.89032e-16
C318 heart_block5_s33 vsse 3.57097e-15
C319 mbk_sig1655 vsse 2.26476e-16
C320 heart_block3_nn3 vsse 4.50376e-15
C321 mbk_sig1626 vsse 7.91856e-16
C322 heart_block3_x23 vsse 2.52104e-15
C323 mbk_sig1623 vsse 7.91856e-16
C324 heart_block3_na20 vsse 3.13049e-15
C325 heart_block3_no23 vsse 2.6393e-15
C326 cini vsse 2.83228e-14
C327 heart_block3_no40 vsse 3.19594e-15
C328 mbk_sig1614 vsse 7.91856e-16
C329 signec vsse 1.69619e-14
C330 heart_block3_signea vsse 6.6893e-15
C331 heart_block4_shacc2 vsse 4.06652e-15
C332 mbk_sig1602 vsse 6.4476e-16
C333 mbk_sig1612 vsse 7.2414e-16
C334 heart_block4_m2_dff_s vsse 5.66676e-16
C335 mbk_sig1610 vsse 2.84472e-16
C336 mbk_sig1603 vsse 7.40988e-16
C337 mbk_sig1609 vsse 1.33164e-15
C338 heart_block4_m2_dff_m vsse 5.51124e-16
C339 mbk_sig1608 vsse 6.82992e-16
C340 heart_block5_a27sh vsse 3.47328e-15
C341 mbk_sig1597 vsse 5.51448e-16
C342 heart_block3_fb0 vsse 7.07648e-15
C343 heart_block3_fb2 vsse 5.13054e-15
C344 mbk_sig1594 vsse 3.00996e-16
C345 mbk_sig1590 vsse 1.35108e-15
C346 heart_block5_m_3_2_dff_m vsse 5.32008e-16
C347 mbk_sig1592 vsse 6.73272e-16
C348 mbk_sig1595 vsse 7.51032e-16
C349 heart_block5_m_3_2_dff_s vsse 5.89032e-16
C350 mbk_sig1587 vsse 2.26476e-16
C351 mbk_sig1588 vsse 5.51448e-16
C352 s3c vsse 1.80479e-14
C353 mbk_sig1586 vsse 5.51448e-16
C354 heart_block5_a28sh vsse 2.77279e-15
C355 mbk_sig1584 vsse 5.51448e-16
C356 q3i vsse 1.21518e-14
C357 mbk_sig1580 vsse 5.51448e-16
C358 mbk_sig1577 vsse 3.00996e-16
C359 mbk_sig1573 vsse 1.35108e-15
C360 heart_block5_m_6_3_dff_m vsse 5.32008e-16
C361 mbk_sig1578 vsse 6.73272e-16
C362 mbk_sig1579 vsse 7.51032e-16
C363 heart_block5_m_6_3_dff_s vsse 5.89032e-16
C364 mbk_sig1575 vsse 2.26476e-16
C365 heart_block4_a211s vsse 3.29443e-15
C366 mbk_sig1572 vsse 5.51448e-16
C367 heart_block4_decalda vsse 1.21301e-14
C368 mbk_sig1567 vsse 6.57072e-16
C369 decaldc vsse 1.21152e-14
C370 heart_block5_s21 vsse 6.65998e-15
C371 heart_block5_b26s vsse 3.25944e-15
C372 mbk_sig1558 vsse 7.75008e-16
C373 heart_block5_b27s vsse 3.52836e-15
C374 heart_block5_b25s vsse 4.26514e-15
C375 mbk_sig1554 vsse 5.51448e-16
C376 mbk_sig1549 vsse 7.75008e-16
C377 heart_block5_b23s vsse 4.82695e-15
C378 heart_block5_b24s vsse 4.2917e-15
C379 heart_block5_b21s vsse 5.12827e-15
C380 heart_b_1 vsse 2.14559e-14
C381 mbk_sig1546 vsse 7.75008e-16
C382 heart_block5_b15s vsse 2.63412e-15
C383 mbk_sig1540 vsse 3.00996e-16
C384 mbk_sig1536 vsse 1.35108e-15
C385 heart_block5_m_7_1_dff_m vsse 5.32008e-16
C386 mbk_sig1538 vsse 6.73272e-16
C387 mbk_sig1542 vsse 7.51032e-16
C388 heart_block5_m_7_1_dff_s vsse 5.89032e-16
C389 heart_block5_s17 vsse 5.03593e-15
C390 mbk_sig1534 vsse 2.26476e-16
C391 mbk_sig1532 vsse 3.00996e-16
C392 mbk_sig1526 vsse 1.35108e-15
C393 heart_block5_m_8_0_dff_m vsse 5.32008e-16
C394 heart_block5_ck8 vsse 1.10654e-14
C395 mbk_sig1533 vsse 6.73272e-16
C396 mbk_sig1535 vsse 7.51032e-16
C397 heart_block5_m_8_0_dff_s vsse 5.89032e-16
C398 mbk_sig1529 vsse 2.26476e-16
C399 heart_block5_b22s vsse 3.97483e-15
C400 heart_block5_s15 vsse 7.90333e-15
C401 mbk_sig1521 vsse 7.75008e-16
C402 heart_block5_a17s vsse 2.5447e-15
C403 heart_block5_a18s vsse 4.69606e-15
C404 heart_block5_a15s vsse 2.4961e-15
C405 heart_block5_b1 vsse 1.64333e-14
C406 mbk_sig1514 vsse 5.51448e-16
C407 heart_block5_s24 vsse 4.54604e-15
C408 heart_block5_s28 vsse 5.18449e-15
C409 heart_block5_b28s vsse 4.92739e-15
C410 mbk_sig1506 vsse 7.75008e-16
C411 heart_block5_b11s vsse 5.62982e-15
C412 heart_block5_b14s vsse 2.93285e-15
C413 heart_block5_s31 vsse 3.98309e-15
C414 mbk_sig1496 vsse 3.00996e-16
C415 mbk_sig1498 vsse 1.35108e-15
C416 heart_block5_m_4_1_dff_m vsse 5.32008e-16
C417 mbk_sig1497 vsse 6.73272e-16
C418 mbk_sig1501 vsse 7.51032e-16
C419 heart_block5_m_4_1_dff_s vsse 5.89032e-16
C420 heart_block5_s14 vsse 4.07365e-15
C421 mbk_sig1493 vsse 2.26476e-16
C422 mbk_sig1491 vsse 7.75008e-16
C423 heart_block5_a33s vsse 4.76086e-15
C424 heart_block5_a31s vsse 2.48832e-15
C425 mbk_sig1486 vsse 3.00996e-16
C426 mbk_sig1481 vsse 1.35108e-15
C427 heart_block5_m_4_3_dff_m vsse 5.32008e-16
C428 heart_block5_ck4 vsse 9.80375e-15
C429 mbk_sig1488 vsse 6.73272e-16
C430 mbk_sig1487 vsse 7.51032e-16
C431 heart_block5_m_4_3_dff_s vsse 5.89032e-16
C432 mbk_sig1483 vsse 2.26476e-16
C433 heart_block5_b4 vsse 1.32801e-14
C434 heart_block5_b34s vsse 2.54794e-15
C435 heart_block5_b32s vsse 2.7715e-15
C436 heart_block5_a32s vsse 3.14863e-15
C437 heart_block5_b12s vsse 4.25671e-15
C438 heart_block3_cout1 vsse 9.18491e-15
C439 heart_block3_na22 vsse 2.0885e-15
C440 heart_block3_no43 vsse 2.74298e-15
C441 heart_block3_n4 vsse 9.83e-15
C442 heart_block3_no33 vsse 3.03264e-15
C443 heart_block3_ni5 vsse 1.06755e-14
C444 ii_3 vsse 2.6145e-14
C445 mbk_sig1435 vsse 1.33164e-16
C446 mbk_sig1434 vsse 7.17012e-16
C447 heart_block3_x20 vsse 3.49304e-15
C448 mbk_sig1429 vsse 7.91856e-16
C449 ngc vsse 2.17707e-14
C450 heart_block4_decaln vsse 1.90224e-14
C451 heart_block4_selalu vsse 1.16851e-14
C452 mbk_sig1426 vsse 6.42492e-16
C453 mbk_sig1413 vsse 6.4476e-16
C454 mbk_sig1421 vsse 7.2414e-16
C455 heart_block4_m3_dff_s vsse 5.66676e-16
C456 mbk_sig1420 vsse 2.84472e-16
C457 mbk_sig1414 vsse 7.40988e-16
C458 mbk_sig1418 vsse 1.33164e-15
C459 heart_block4_m3_dff_m vsse 5.51124e-16
C460 mbk_sig1417 vsse 6.82992e-16
C461 mbk_sig1409 vsse 5.51448e-16
C462 mbk_sig1407 vsse 5.51448e-16
C463 heart_block4_shacc0 vsse 1.1444e-14
C464 mbk_sig1397 vsse 6.4476e-16
C465 scini vsse 1.04986e-14
C466 mbk_sig1406 vsse 7.2414e-16
C467 heart_block4_m0_dff_s vsse 5.66676e-16
C468 mbk_sig1404 vsse 2.84472e-16
C469 mbk_sig1398 vsse 7.40988e-16
C470 mbk_sig1403 vsse 1.33164e-15
C471 heart_block4_m0_dff_m vsse 5.51124e-16
C472 mbk_sig1402 vsse 6.82992e-16
C473 heart_block4_shacc3 vsse 3.12368e-15
C474 heart_block4_a217s vsse 1.14806e-14
C475 heart_block4_a216s vsse 2.64676e-15
C476 mbk_sig1389 vsse 7.12152e-16
C477 oec vsse 2.31843e-14
C478 noei vsse 1.78767e-14
C479 heart_block4_a218s vsse 2.82334e-15
C480 heart_block4_insh2 vsse 1.49926e-14
C481 mbk_sig1387 vsse 5.51448e-16
C482 mbk_sig1385 vsse 5.51448e-16
C483 scoutc vsse 2.34082e-14
C484 mbk_sig1384 vsse 5.51448e-16
C485 heart_block4_a210s vsse 3.80894e-15
C486 heart_block4_a214s vsse 2.79677e-15
C487 heart_block4_insh0 vsse 1.69217e-14
C488 mbk_sig1378 vsse 5.68296e-16
C489 heart_block5_b16s vsse 6.68477e-15
C490 heart_block5_s23 vsse 5.936e-15
C491 mbk_sig1371 vsse 7.75008e-16
C492 heart_block5_a23s vsse 2.69633e-15
C493 heart_block5_a24s vsse 6.71587e-15
C494 heart_block5_a21s vsse 2.91211e-15
C495 heart_block5_nb1 vsse 2.01927e-14
C496 mbk_sig1360 vsse 7.75008e-16
C497 heart_block5_nb2 vsse 1.65917e-14
C498 heart_b_3 vsse 2.41406e-14
C499 heart_block5_nb0 vsse 1.69755e-14
C500 mbk_sig1356 vsse 7.75008e-16
C501 heart_block5_b06s vsse 4.23533e-15
C502 mbk_sig1350 vsse 7.75008e-16
C503 heart_block5_b07s vsse 2.20838e-15
C504 heart_block5_b05s vsse 2.05092e-15
C505 mbk_sig1347 vsse 3.00996e-16
C506 mbk_sig1343 vsse 1.35108e-15
C507 heart_block5_m_7_0_dff_m vsse 5.32008e-16
C508 mbk_sig1345 vsse 6.73272e-16
C509 mbk_sig1348 vsse 7.51032e-16
C510 heart_block5_m_7_0_dff_s vsse 5.89032e-16
C511 mbk_sig1342 vsse 2.26476e-16
C512 heart_block5_a22s vsse 5.75942e-15
C513 heart_block5_s07 vsse 5.00288e-15
C514 heart_block5_a07s vsse 4.06879e-15
C515 heart_block5_s11 vsse 1.14881e-14
C516 heart_block5_a05s vsse 4.16988e-15
C517 mbk_sig1333 vsse 7.75008e-16
C518 heart_block5_a14s vsse 3.69878e-15
C519 heart_block5_a11s vsse 2.86351e-15
C520 heart_block5_a13s vsse 2.2181e-15
C521 mbk_sig1326 vsse 3.00996e-16
C522 mbk_sig1325 vsse 1.35108e-15
C523 heart_block5_m_3_1_dff_m vsse 5.32008e-16
C524 mbk_sig1328 vsse 6.73272e-16
C525 mbk_sig1330 vsse 7.51032e-16
C526 heart_block5_m_3_1_dff_s vsse 5.89032e-16
C527 mbk_sig1322 vsse 2.26476e-16
C528 heart_block5_s13 vsse 3.61487e-15
C529 heart_block5_b13s vsse 2.62246e-15
C530 heart_block5_s01 vsse 6.8816e-15
C531 heart_block5_a36s vsse 7.01525e-15
C532 mbk_sig1317 vsse 7.75008e-16
C533 heart_block5_a38s vsse 1.06194e-14
C534 mbk_sig1312 vsse 7.75008e-16
C535 heart_block5_b04s vsse 6.50981e-15
C536 heart_block5_b01s vsse 3.82968e-15
C537 heart_block5_b2 vsse 1.70068e-14
C538 heart_block5_b02s vsse 2.88814e-15
C539 heart_block5_a35s vsse 2.84213e-15
C540 heart_block5_b3 vsse 2.09539e-14
C541 heart_block5_b03s vsse 2.71966e-15
C542 mbk_sig1300 vsse 3.00996e-16
C543 mbk_sig1296 vsse 1.35108e-15
C544 heart_block5_m_2_2_dff_m vsse 5.32008e-16
C545 mbk_sig1302 vsse 6.73272e-16
C546 mbk_sig1301 vsse 7.51032e-16
C547 heart_block5_m_2_2_dff_s vsse 5.89032e-16
C548 heart_block5_s22 vsse 5.96516e-15
C549 mbk_sig1298 vsse 2.26476e-16
C550 heart_block5_s34 vsse 3.99784e-15
C551 heart_block5_a34s vsse 3.0281e-15
C552 mbk_sig1288 vsse 7.75008e-16
C553 heart_block5_a03s vsse 3.20371e-15
C554 heart_block5_a04s vsse 8.16026e-15
C555 heart_block5_a01s vsse 3.87245e-15
C556 mbk_sig1283 vsse 3.00996e-16
C557 mbk_sig1280 vsse 1.35108e-15
C558 heart_block5_m_3_0_dff_m vsse 5.32008e-16
C559 heart_block5_ck3 vsse 2.64052e-14
C560 mbk_sig1285 vsse 6.73272e-16
C561 mbk_sig1284 vsse 7.51032e-16
C562 heart_block5_m_3_0_dff_s vsse 5.89032e-16
C563 heart_block5_s03 vsse 4.7696e-15
C564 mbk_sig1279 vsse 2.26476e-16
C565 heart_block3_not2 vsse 3.07573e-15
C566 mbk_sig1220 vsse 6.57072e-16
C567 decalgrc vsse 1.81762e-14
C568 heart_block3_not0 vsse 6.1628e-15
C569 heart_block3_gb1 vsse 1.16974e-14
C570 heart_block3_no31_csh vsse 2.1883e-15
C571 heart_block3_ngb3 vsse 2.12058e-15
C572 ii_5 vsse 2.38595e-14
C573 ii_4 vsse 2.96873e-14
C574 mbk_sig1217 vsse 1.33164e-16
C575 mbk_sig1216 vsse 7.17012e-16
C576 heart_block3_no20 vsse 3.99427e-15
C577 heart_block3_n2 vsse 1.06761e-14
C578 heart_block3_nn0 vsse 4.32022e-15
C579 heart_block3_pb1 vsse 1.11728e-14
C580 heart_block3_no32 vsse 3.06569e-15
C581 heart_block3_no22 vsse 3.65407e-15
C582 heart_block3_x22 vsse 1.02407e-14
C583 mbk_sig1209 vsse 7.91856e-16
C584 mbk_sig1208 vsse 5.51448e-16
C585 heart_block5_a214sh vsse 3.23352e-15
C586 heart_block5_a213sh vsse 1.72951e-15
C587 mbk_sig1205 vsse 7.12152e-16
C588 mbk_sig1204 vsse 5.51448e-16
C589 heart_block5_a211sh vsse 1.65499e-15
C590 heart_block5_a29sh vsse 3.02972e-15
C591 mbk_sig1202 vsse 7.12152e-16
C592 heart_block5_a210sh vsse 1.86365e-15
C593 mbk_sig1199 vsse 5.51448e-16
C594 heart_block5_a212sh vsse 2.46791e-15
C595 r0i vsse 1.76011e-14
C596 mbk_sig1197 vsse 5.51448e-16
C597 mbk_sig1194 vsse 5.51448e-16
C598 heart_block5_decalnr vsse 1.21165e-14
C599 mbk_sig1192 vsse 5.68296e-16
C600 mbk_sig1191 vsse 5.51448e-16
C601 heart_block5_a24sh vsse 2.39825e-15
C602 mbk_sig1190 vsse 7.12152e-16
C603 heart_block4_ni7 vsse 1.79169e-14
C604 heart_block5_a23sh vsse 2.75368e-15
C605 mbk_sig1186 vsse 5.51448e-16
C606 heart_block5_decalgra vsse 1.64932e-14
C607 heart_block5_s36 vsse 6.85049e-15
C608 heart_block5_a25sh vsse 3.73702e-15
C609 r3i vsse 1.47801e-14
C610 mbk_sig1181 vsse 5.51448e-16
C611 mbk_sig1176 vsse 3.00996e-16
C612 mbk_sig1178 vsse 1.35108e-15
C613 heart_block5_m_7_2_dff_m vsse 5.32008e-16
C614 mbk_sig1177 vsse 6.73272e-16
C615 mbk_sig1180 vsse 7.51032e-16
C616 heart_block5_m_7_2_dff_s vsse 5.89032e-16
C617 mbk_sig1174 vsse 2.26476e-16
C618 mbk_sig1172 vsse 5.51448e-16
C619 heart_block5_b6 vsse 1.25616e-14
C620 heart_block5_a06s vsse 3.45578e-15
C621 mbk_sig1166 vsse 3.00996e-16
C622 mbk_sig1162 vsse 1.35108e-15
C623 heart_block5_m_6_1_dff_m vsse 5.32008e-16
C624 mbk_sig1168 vsse 6.73272e-16
C625 mbk_sig1167 vsse 7.51032e-16
C626 heart_block5_m_6_1_dff_s vsse 5.89032e-16
C627 mbk_sig1164 vsse 2.26476e-16
C628 mbk_sig1159 vsse 7.75008e-16
C629 heart_block5_a28s vsse 1.43364e-14
C630 heart_block5_a26s vsse 2.73262e-15
C631 heart_block5_s27 vsse 1.04586e-14
C632 heart_block5_a27s vsse 3.67416e-15
C633 heart_block5_a08s vsse 3.67934e-15
C634 heart_block5_s16 vsse 7.46204e-15
C635 heart_block5_a16s vsse 8.79984e-15
C636 heart_block5_s08 vsse 9.39827e-15
C637 heart_block5_b8 vsse 3.4703e-14
C638 heart_block5_b08s vsse 3.67934e-15
C639 mbk_sig1142 vsse 3.00996e-16
C640 mbk_sig1138 vsse 1.35108e-15
C641 heart_block5_m_5_0_dff_m vsse 5.32008e-16
C642 mbk_sig1140 vsse 6.73272e-16
C643 mbk_sig1144 vsse 7.51032e-16
C644 heart_block5_m_5_0_dff_s vsse 5.89032e-16
C645 heart_block5_s05 vsse 4.98928e-15
C646 mbk_sig1137 vsse 2.26476e-16
C647 heart_block5_b5 vsse 1.32051e-14
C648 heart_block5_s25 vsse 1.41716e-14
C649 heart_block5_a25s vsse 4.3254e-15
C650 mbk_sig1130 vsse 3.00996e-16
C651 mbk_sig1127 vsse 1.35108e-15
C652 heart_block5_m_11_3_dff_m vsse 5.32008e-16
C653 mbk_sig1131 vsse 6.73272e-16
C654 mbk_sig1133 vsse 7.51032e-16
C655 heart_block5_m_11_3_dff_s vsse 5.89032e-16
C656 mbk_sig1125 vsse 2.26476e-16
C657 mbk_sig1122 vsse 3.00996e-16
C658 mbk_sig1118 vsse 1.35108e-15
C659 heart_block5_m_5_3_dff_m vsse 5.32008e-16
C660 heart_block5_ck5 vsse 2.32096e-14
C661 mbk_sig1124 vsse 6.73272e-16
C662 mbk_sig1123 vsse 7.51032e-16
C663 heart_block5_m_5_3_dff_s vsse 5.89032e-16
C664 heart_block5_s35 vsse 5.95544e-15
C665 mbk_sig1117 vsse 2.26476e-16
C666 mbk_sig1115 vsse 3.00996e-16
C667 mbk_sig1111 vsse 1.35108e-15
C668 heart_block5_m_2_0_dff_m vsse 5.32008e-16
C669 mbk_sig1113 vsse 6.73272e-16
C670 mbk_sig1116 vsse 7.51032e-16
C671 heart_block5_m_2_0_dff_s vsse 5.89032e-16
C672 mbk_sig1110 vsse 2.26476e-16
C673 mbk_sig1105 vsse 3.00996e-16
C674 mbk_sig1107 vsse 1.35108e-15
C675 heart_block5_m_2_1_dff_m vsse 5.32008e-16
C676 mbk_sig1106 vsse 6.73272e-16
C677 mbk_sig1109 vsse 7.51032e-16
C678 heart_block5_m_2_1_dff_s vsse 5.89032e-16
C679 mbk_sig1101 vsse 2.26476e-16
C680 heart_block5_s12 vsse 1.78185e-14
C681 heart_block5_a12s vsse 5.3784e-15
C682 mbk_sig1097 vsse 5.51448e-16
C683 mbk_sig1094 vsse 3.00996e-16
C684 mbk_sig1090 vsse 1.35108e-15
C685 heart_block5_m_10_3_dff_m vsse 5.32008e-16
C686 mbk_sig1095 vsse 6.73272e-16
C687 mbk_sig1096 vsse 7.51032e-16
C688 heart_block5_m_10_3_dff_s vsse 5.89032e-16
C689 mbk_sig1092 vsse 2.26476e-16
C690 heart_block5_s02 vsse 6.2626e-15
C691 heart_block5_a02s vsse 3.54521e-15
C692 heart_block3_na23 vsse 2.02241e-15
C693 heart_block3_no30 vsse 6.21108e-15
C694 heart_block3_n3 vsse 1.42772e-14
C695 mbk_sig1050 vsse 7.12152e-16
C696 heart_s_1 vsse 2.4125e-15
C697 heart_block3_x11 vsse 6.8965e-15
C698 mbk_sig1049 vsse 7.91856e-16
C699 heart_block3_cout2 vsse 9.39146e-15
C700 ovrc vsse 9.05693e-15
C701 mbk_sig1046 vsse 7.91856e-16
C702 heart_block1_srq1 vsse 2.78446e-15
C703 heart_q_1 vsse 1.28777e-14
C704 mbk_sig1042 vsse 5.51448e-16
C705 heart_block3_no2_csh vsse 4.19872e-15
C706 heart_block3_gb0 vsse 1.31481e-14
C707 npc vsse 1.89354e-14
C708 coutc vsse 8.94386e-15
C709 heart_block3_couta vsse 5.07967e-15
C710 mbk_sig1037 vsse 5.51448e-16
C711 mbk_sig1035 vsse 6.57072e-16
C712 decaldrc vsse 1.53953e-14
C713 heart_block3_p vsse 2.22361e-15
C714 heart_block3_propf vsse 2.27156e-15
C715 mbk_sig1034 vsse 5.51448e-16
C716 heart_block2_a28ms_i0 vsse 1.52857e-14
C717 mbk_sig1030 vsse 5.51448e-16
C718 mbk_sig1028 vsse 5.51448e-16
C719 heart_block5_ni7 vsse 2.05254e-15
C720 heart_block2_syalu3 vsse 1.78589e-15
C721 yc_3 vsse 1.81707e-14
C722 mbk_sig1023 vsse 5.68296e-16
C723 s0c vsse 1.47104e-14
C724 heart_block5_decaldra vsse 1.51285e-14
C725 mbk_sig1022 vsse 5.51448e-16
C726 heart_q_0 vsse 1.14714e-14
C727 mbk_sig1020 vsse 5.51448e-16
C728 heart_block4_decalga vsse 3.24146e-14
C729 mbk_sig1016 vsse 5.51448e-16
C730 mbk_sig1013 vsse 5.51448e-16
C731 mbk_sig1012 vsse 5.51448e-16
C732 mbk_sig1011 vsse 5.51448e-16
C733 mbk_sig1003 vsse 3.00996e-16
C734 mbk_sig1002 vsse 1.35108e-15
C735 heart_block5_m_6_0_dff_m vsse 5.32008e-16
C736 mbk_sig1004 vsse 6.73272e-16
C737 mbk_sig1008 vsse 7.51032e-16
C738 heart_block5_m_6_0_dff_s vsse 5.89032e-16
C739 heart_block5_s06 vsse 7.27623e-15
C740 mbk_sig1000 vsse 2.26476e-16
C741 mbk_sig994 vsse 7.75008e-16
C742 heart_block5_b316s vsse 2.37686e-15
C743 heart_block5_b313s vsse 3.64889e-15
C744 mbk_sig991 vsse 3.00996e-16
C745 mbk_sig990 vsse 1.35108e-15
C746 heart_block5_m_16_3_dff_m vsse 5.32008e-16
C747 mbk_sig989 vsse 6.73272e-16
C748 mbk_sig993 vsse 7.51032e-16
C749 heart_block5_m_16_3_dff_s vsse 5.89032e-16
C750 mbk_sig987 vsse 2.26476e-16
C751 heart_block5_ob442s vsse 6.7865e-15
C752 heart_block5_ob432s vsse 8.79109e-15
C753 heart_block5_b315s vsse 4.77252e-15
C754 heart_block5_b36s vsse 5.48532e-15
C755 mbk_sig974 vsse 7.75008e-16
C756 heart_block5_b38s vsse 1.45424e-14
C757 heart_block5_b35s vsse 4.02991e-15
C758 mbk_sig969 vsse 3.00996e-16
C759 mbk_sig971 vsse 1.35108e-15
C760 heart_block5_m_7_3_dff_m vsse 5.32008e-16
C761 heart_block5_ck7 vsse 1.60779e-14
C762 mbk_sig970 vsse 6.73272e-16
C763 mbk_sig973 vsse 7.51032e-16
C764 heart_block5_m_7_3_dff_s vsse 5.89032e-16
C765 mbk_sig967 vsse 2.26476e-16
C766 heart_block5_ob443s vsse 1.22783e-14
C767 heart_block5_ob433s vsse 3.18071e-15
C768 heart_block5_ob413s vsse 4.57067e-15
C769 heart_rb_3 vsse 7.73647e-15
C770 mbk_sig958 vsse 3.00996e-16
C771 mbk_sig955 vsse 1.35108e-15
C772 heart_block5_m_11_2_dff_m vsse 5.32008e-16
C773 mbk_sig960 vsse 6.73272e-16
C774 mbk_sig961 vsse 7.51032e-16
C775 heart_block5_m_11_2_dff_s vsse 5.89032e-16
C776 mbk_sig957 vsse 2.26476e-16
C777 heart_block5_a3 vsse 3.0277e-14
C778 mbk_sig952 vsse 7.75008e-16
C779 heart_block5_a5 vsse 1.08459e-14
C780 mbk_sig948 vsse 7.75008e-16
C781 heart_block5_a37s vsse 1.66659e-14
C782 heart_block5_ob422s vsse 6.12781e-15
C783 mbk_sig937 vsse 7.75008e-16
C784 heart_block5_b211s vsse 3.13373e-15
C785 heart_block5_b29s vsse 3.50698e-15
C786 heart_block5_a7 vsse 2.3576e-14
C787 mbk_sig933 vsse 7.75008e-16
C788 heart_block5_b210s vsse 3.15641e-15
C789 heart_block5_a4 vsse 3.03151e-14
C790 mbk_sig927 vsse 7.75008e-16
C791 heart_block5_s311 vsse 5.62966e-15
C792 heart_block5_ob423s vsse 4.92836e-15
C793 heart_block5_b310s vsse 2.96006e-15
C794 mbk_sig918 vsse 7.75008e-16
C795 heart_block5_b311s vsse 2.88684e-15
C796 mbk_sig913 vsse 3.00996e-16
C797 mbk_sig915 vsse 1.35108e-15
C798 heart_block5_m_10_0_dff_m vsse 5.32008e-16
C799 mbk_sig914 vsse 6.73272e-16
C800 mbk_sig917 vsse 7.51032e-16
C801 heart_block5_m_10_0_dff_s vsse 5.89032e-16
C802 mbk_sig911 vsse 2.26476e-16
C803 mbk_sig907 vsse 3.00996e-16
C804 mbk_sig906 vsse 1.35108e-15
C805 heart_block5_m_10_1_dff_m vsse 5.32008e-16
C806 mbk_sig908 vsse 6.73272e-16
C807 mbk_sig910 vsse 7.51032e-16
C808 heart_block5_m_10_1_dff_s vsse 5.89032e-16
C809 mbk_sig905 vsse 2.26476e-16
C810 mbk_sig866 vsse 7.91856e-16
C811 heart_block3_x00 vsse 3.77249e-15
C812 heart_block3_not3 vsse 3.12239e-15
C813 mbk_sig861 vsse 5.51448e-16
C814 heart_block3_no32_csh vsse 4.80686e-15
C815 heart_block3_ngb0 vsse 4.06134e-15
C816 heart_block3_na_csh vsse 2.01722e-15
C817 heart_block3_pb2 vsse 1.03072e-14
C818 mbk_sig853 vsse 7.91856e-16
C819 heart_block3_pb3 vsse 1.27844e-14
C820 heart_block3_x03 vsse 3.1496e-15
C821 heart_block3_gb3 vsse 1.15587e-14
C822 heart_block3_ngen vsse 3.53776e-15
C823 heart_block3_g vsse 1.14207e-14
C824 heart_block3_genf vsse 2.20352e-15
C825 mbk_sig844 vsse 5.51448e-16
C826 heart_block3_flag vsse 1.75822e-14
C827 heart_block3_no30_csh vsse 7.33957e-15
C828 heart_block3_nprop vsse 2.81426e-15
C829 heart_block3_x13 vsse 3.80279e-15
C830 mbk_sig837 vsse 7.91856e-16
C831 heart_s_3 vsse 3.00348e-15
C832 heart_block1_srb3 vsse 3.97062e-15
C833 mbk_sig832 vsse 7.12152e-16
C834 heart_block1_srq3 vsse 2.03407e-15
C835 heart_q_3 vsse 1.27635e-14
C836 mbk_sig830 vsse 5.51448e-16
C837 mbk_sig828 vsse 3.00996e-16
C838 mbk_sig824 vsse 1.35108e-15
C839 heart_block5_m_13_0_dff_m vsse 5.32008e-16
C840 mbk_sig826 vsse 6.73272e-16
C841 mbk_sig829 vsse 7.51032e-16
C842 heart_block5_m_13_0_dff_s vsse 5.89032e-16
C843 mbk_sig822 vsse 2.26476e-16
C844 mbk_sig820 vsse 3.00996e-16
C845 mbk_sig815 vsse 1.35108e-15
C846 heart_block5_m_13_2_dff_m vsse 5.32008e-16
C847 mbk_sig821 vsse 6.73272e-16
C848 mbk_sig823 vsse 7.51032e-16
C849 heart_block5_m_13_2_dff_s vsse 5.89032e-16
C850 mbk_sig818 vsse 2.26476e-16
C851 mbk_sig810 vsse 3.00996e-16
C852 mbk_sig812 vsse 1.35108e-15
C853 heart_block5_m_16_1_dff_m vsse 5.32008e-16
C854 mbk_sig811 vsse 6.73272e-16
C855 mbk_sig814 vsse 7.51032e-16
C856 heart_block5_m_16_1_dff_s vsse 5.89032e-16
C857 mbk_sig808 vsse 2.26476e-16
C858 heart_block5_s213 vsse 4.96984e-15
C859 mbk_sig799 vsse 3.00996e-16
C860 mbk_sig801 vsse 1.35108e-15
C861 heart_block5_m_6_2_dff_m vsse 5.32008e-16
C862 heart_block5_ck6 vsse 1.76194e-14
C863 mbk_sig800 vsse 6.73272e-16
C864 mbk_sig804 vsse 7.51032e-16
C865 heart_block5_m_6_2_dff_s vsse 5.89032e-16
C866 heart_block5_s26 vsse 1.49959e-14
C867 mbk_sig796 vsse 2.26476e-16
C868 heart_block5_ob412s vsse 2.79968e-15
C869 heart_block5_b214s vsse 3.96511e-15
C870 mbk_sig793 vsse 7.75008e-16
C871 heart_block5_b216s vsse 3.2711e-15
C872 heart_block5_b213s vsse 4.32734e-15
C873 mbk_sig787 vsse 7.75008e-16
C874 heart_block5_a216s vsse 2.45462e-15
C875 heart_block5_a213s vsse 4.7803e-15
C876 heart_block5_ob440s vsse 1.10827e-14
C877 heart_block5_ob430s vsse 8.61613e-15
C878 mbk_sig779 vsse 7.75008e-16
C879 heart_block5_b115s vsse 2.48443e-15
C880 heart_block5_b116s vsse 6.11712e-15
C881 heart_block5_b113s vsse 6.18192e-15
C882 heart_block5_oa440s vsse 1.1038e-14
C883 heart_block5_oa430s vsse 1.07176e-14
C884 heart_block5_s37 vsse 6.04681e-15
C885 heart_block5_b7 vsse 2.64215e-14
C886 heart_block5_b37s vsse 3.4992e-15
C887 mbk_sig773 vsse 5.51448e-16
C888 heart_block5_a8 vsse 4.11674e-14
C889 mbk_sig768 vsse 7.75008e-16
C890 mbk_sig762 vsse 3.00996e-16
C891 mbk_sig764 vsse 1.35108e-15
C892 heart_block5_m_15_1_dff_m vsse 5.32008e-16
C893 mbk_sig763 vsse 6.73272e-16
C894 mbk_sig767 vsse 7.51032e-16
C895 heart_block5_m_15_1_dff_s vsse 5.89032e-16
C896 mbk_sig759 vsse 2.26476e-16
C897 mbk_sig758 vsse 5.51448e-16
C898 mbk_sig753 vsse 3.00996e-16
C899 mbk_sig755 vsse 1.35108e-15
C900 heart_block5_m_9_3_dff_m vsse 5.32008e-16
C901 mbk_sig754 vsse 6.73272e-16
C902 mbk_sig757 vsse 7.51032e-16
C903 heart_block5_m_9_3_dff_s vsse 5.89032e-16
C904 mbk_sig750 vsse 2.26476e-16
C905 heart_block5_a1 vsse 3.24855e-14
C906 mbk_sig749 vsse 7.75008e-16
C907 mbk_sig743 vsse 3.00996e-16
C908 mbk_sig738 vsse 1.35108e-15
C909 heart_block5_m_10_2_dff_m vsse 5.32008e-16
C910 heart_block5_ck10 vsse 1.04266e-14
C911 mbk_sig745 vsse 6.73272e-16
C912 mbk_sig744 vsse 7.51032e-16
C913 heart_block5_m_10_2_dff_s vsse 5.89032e-16
C914 mbk_sig740 vsse 2.26476e-16
C915 mbk_sig736 vsse 7.75008e-16
C916 heart_block5_b39s vsse 2.82852e-15
C917 heart_block5_s210 vsse 4.72878e-15
C918 heart_block5_a2 vsse 3.32337e-14
C919 mbk_sig729 vsse 7.75008e-16
C920 heart_block5_b312s vsse 3.27888e-15
C921 mbk_sig721 vsse 7.75008e-16
C922 heart_block5_s010 vsse 6.65221e-15
C923 mbk_sig667 vsse 7.91856e-16
C924 heart_block3_nn1 vsse 7.17984e-15
C925 heart_block1_srq0 vsse 7.77082e-15
C926 mbk_sig663 vsse 7.12152e-16
C927 heart_block3_n1 vsse 1.17228e-14
C928 heart_s_0 vsse 2.49026e-15
C929 heart_block3_x10 vsse 5.22077e-15
C930 mbk_sig662 vsse 7.91856e-16
C931 heart_block3_npb0 vsse 3.64921e-15
C932 heart_block3_pb0 vsse 7.87126e-15
C933 heart_block1_sra0 vsse 2.7229e-15
C934 mbk_sig656 vsse 5.51448e-16
C935 heart_block4_ckin vsse 1.77648e-14
C936 mbk_sig654 vsse 5.51448e-16
C937 heart_block3_x12 vsse 5.32105e-15
C938 heart_block3_gb2 vsse 1.08939e-14
C939 heart_block4_w vsse 2.3396e-15
C940 mbk_sig648 vsse 5.68296e-16
C941 mbk_sig646 vsse 5.51448e-16
C942 heart_block4_a231s vsse 2.6879e-15
C943 mbk_sig642 vsse 5.51448e-16
C944 heart_block4_waccu vsse 2.21454e-15
C945 heart_block4_o21s vsse 1.31729e-14
C946 mbk_sig641 vsse 5.51448e-16
C947 heart_block4_ni6 vsse 1.34876e-14
C948 fonci vsse 1.19705e-14
C949 heart_block2_syra3 vsse 7.02821e-15
C950 mbk_sig639 vsse 5.51448e-16
C951 heart_block2_a27ms_i0 vsse 2.67835e-14
C952 mbk_sig634 vsse 5.51448e-16
C953 heart_block2_a25ms_i0 vsse 1.50715e-14
C954 mbk_sig630 vsse 5.51448e-16
C955 mbk_sig628 vsse 5.51448e-16
C956 heart_block2_syra0 vsse 1.64138e-15
C957 heart_block2_syalu0 vsse 2.40797e-15
C958 yc_0 vsse 1.69062e-14
C959 mbk_sig624 vsse 5.68296e-16
C960 heart_rb_2 vsse 1.4107e-14
C961 mbk_sig623 vsse 5.51448e-16
C962 heart_block1_srb0 vsse 5.4189e-15
C963 heart_rb_0 vsse 6.32124e-15
C964 mbk_sig621 vsse 5.51448e-16
C965 mbk_sig617 vsse 3.00996e-16
C966 mbk_sig612 vsse 1.35108e-15
C967 heart_block5_m_13_1_dff_m vsse 5.32008e-16
C968 mbk_sig614 vsse 6.73272e-16
C969 mbk_sig619 vsse 7.51032e-16
C970 heart_block5_m_13_1_dff_s vsse 5.89032e-16
C971 heart_block5_s113 vsse 5.93293e-15
C972 mbk_sig609 vsse 2.26476e-16
C973 heart_block1_srb1 vsse 1.03605e-14
C974 mbk_sig610 vsse 5.51448e-16
C975 heart_block5_a13 vsse 1.43424e-14
C976 heart_block5_ob410s vsse 4.802e-15
C977 mbk_sig605 vsse 7.75008e-16
C978 mbk_sig597 vsse 3.00996e-16
C979 mbk_sig593 vsse 1.35108e-15
C980 heart_block5_m_16_2_dff_m vsse 5.32008e-16
C981 mbk_sig595 vsse 6.73272e-16
C982 mbk_sig599 vsse 7.51032e-16
C983 heart_block5_m_16_2_dff_s vsse 5.89032e-16
C984 heart_block5_s216 vsse 5.35167e-15
C985 mbk_sig596 vsse 2.26476e-16
C986 heart_block5_a214s vsse 3.98455e-15
C987 mbk_sig589 vsse 7.75008e-16
C988 heart_block5_a313s vsse 5.76202e-15
C989 heart_block5_s316 vsse 7.57755e-15
C990 heart_block5_a316s vsse 2.79871e-15
C991 heart_block5_s013 vsse 7.57561e-15
C992 heart_block5_b13 vsse 2.6747e-14
C993 heart_block5_b013s vsse 4.75114e-15
C994 heart_block5_a315s vsse 2.87518e-15
C995 heart_block5_s115 vsse 5.39168e-15
C996 heart_block5_b215s vsse 3.13178e-15
C997 heart_block5_ob441s vsse 1.30054e-14
C998 heart_block5_ob431s vsse 1.32137e-14
C999 heart_block5_ob411s vsse 2.90077e-15
C1000 heart_rb_1 vsse 5.31814e-15
C1001 mbk_sig569 vsse 5.51448e-16
C1002 mbk_sig566 vsse 7.75008e-16
C1003 heart_block5_oa441s vsse 1.62207e-14
C1004 heart_block5_oa431s vsse 1.78735e-14
C1005 mbk_sig556 vsse 3.00996e-16
C1006 mbk_sig553 vsse 1.35108e-15
C1007 heart_block5_m_15_2_dff_m vsse 5.32008e-16
C1008 mbk_sig558 vsse 6.73272e-16
C1009 mbk_sig559 vsse 7.51032e-16
C1010 heart_block5_m_15_2_dff_s vsse 5.89032e-16
C1011 mbk_sig555 vsse 2.26476e-16
C1012 mbk_sig549 vsse 3.00996e-16
C1013 mbk_sig546 vsse 1.35108e-15
C1014 heart_block5_m_15_3_dff_m vsse 5.32008e-16
C1015 mbk_sig548 vsse 6.73272e-16
C1016 mbk_sig552 vsse 7.51032e-16
C1017 heart_block5_m_15_3_dff_s vsse 5.89032e-16
C1018 heart_block5_s315 vsse 8.27545e-15
C1019 mbk_sig543 vsse 2.26476e-16
C1020 mbk_sig540 vsse 3.00996e-16
C1021 mbk_sig542 vsse 1.35108e-15
C1022 heart_block5_m_9_2_dff_m vsse 5.32008e-16
C1023 mbk_sig541 vsse 6.73272e-16
C1024 mbk_sig545 vsse 7.51032e-16
C1025 heart_block5_m_9_2_dff_s vsse 5.89032e-16
C1026 mbk_sig539 vsse 2.26476e-16
C1027 heart_block5_a6 vsse 2.41226e-14
C1028 mbk_sig536 vsse 7.75008e-16
C1029 heart_block5_na3 vsse 1.58036e-14
C1030 mbk_sig528 vsse 7.75008e-16
C1031 heart_block5_oa443s vsse 2.58824e-14
C1032 heart_block5_oa433s vsse 2.10655e-14
C1033 heart_block5_oa413s vsse 5.86732e-15
C1034 heart_block5_oa423s vsse 2.5353e-15
C1035 mbk_sig517 vsse 7.75008e-16
C1036 heart_block5_a311s vsse 4.72586e-15
C1037 heart_block5_a312s vsse 2.14358e-15
C1038 heart_block5_s39 vsse 5.29448e-15
C1039 heart_block5_a39s vsse 2.05092e-15
C1040 mbk_sig514 vsse 7.75008e-16
C1041 heart_block5_b212s vsse 6.2707e-15
C1042 mbk_sig504 vsse 3.00996e-16
C1043 mbk_sig502 vsse 1.35108e-15
C1044 heart_block5_m_2_3_dff_m vsse 5.32008e-16
C1045 heart_block5_ck2 vsse 3.90608e-14
C1046 mbk_sig505 vsse 6.73272e-16
C1047 mbk_sig507 vsse 7.51032e-16
C1048 heart_block5_m_2_3_dff_s vsse 5.89032e-16
C1049 heart_block5_s32 vsse 2.76396e-14
C1050 mbk_sig501 vsse 2.26476e-16
C1051 heart_r_0 vsse 4.80622e-15
C1052 mbk_sig465 vsse 5.68296e-16
C1053 yc_1 vsse 2.30411e-14
C1054 mbk_sig463 vsse 5.68296e-16
C1055 heart_block2_syra1 vsse 2.11961e-15
C1056 mbk_sig461 vsse 5.51448e-16
C1057 heart_block2_syalu1 vsse 2.32049e-15
C1058 heart_block2_a26ms_i0 vsse 2.1909e-14
C1059 mbk_sig458 vsse 5.51448e-16
C1060 heart_block2_selaluy vsse 1.71581e-14
C1061 heart_block1_ssa0 vsse 2.63477e-15
C1062 heart_ra_0 vsse 1.33187e-14
C1063 mbk_sig455 vsse 5.51448e-16
C1064 cko vsse 1.72065e-14
C1065 mbk_sig453 vsse 5.67972e-16
C1066 heart_block1_sra1 vsse 6.62839e-15
C1067 mbk_sig450 vsse 5.51448e-16
C1068 heart_block5_wram vsse 2.33896e-15
C1069 heart_fonc_mode vsse 4.18171e-15
C1070 mbk_sig446 vsse 5.51448e-16
C1071 heart_block3_x02 vsse 4.88641e-15
C1072 mbk_sig443 vsse 7.91856e-16
C1073 heart_block1_sra3 vsse 4.72327e-15
C1074 mbk_sig440 vsse 5.51448e-16
C1075 heart_block5_o21s vsse 2.75368e-15
C1076 mbk_sig437 vsse 5.68296e-16
C1077 heart_q_2 vsse 1.83462e-14
C1078 mbk_sig436 vsse 5.51448e-16
C1079 heart_ra_3 vsse 1.38466e-14
C1080 mbk_sig433 vsse 5.51448e-16
C1081 heart_s_2 vsse 6.17998e-15
C1082 heart_block1_srq2 vsse 2.38982e-15
C1083 heart_block1_srb2 vsse 3.37381e-15
C1084 mbk_sig430 vsse 7.12152e-16
C1085 heart_block1_sra2 vsse 2.33021e-15
C1086 mbk_sig428 vsse 5.51448e-16
C1087 mbk_sig422 vsse 3.00996e-16
C1088 mbk_sig424 vsse 1.35108e-15
C1089 heart_block5_m_13_3_dff_m vsse 5.32008e-16
C1090 heart_block5_ck13 vsse 1.05822e-14
C1091 mbk_sig423 vsse 6.73272e-16
C1092 mbk_sig426 vsse 7.51032e-16
C1093 heart_block5_m_13_3_dff_s vsse 5.89032e-16
C1094 heart_block5_s313 vsse 1.02408e-14
C1095 mbk_sig419 vsse 2.26476e-16
C1096 heart_block4_test_mode vsse 2.98666e-14
C1097 mbk_sig416 vsse 5.51448e-16
C1098 heart_block4_n14s vsse 3.64079e-15
C1099 heart_block4_n15s vsse 4.4456e-15
C1100 testi vsse 1.71266e-14
C1101 mbk_sig410 vsse 3.00996e-16
C1102 mbk_sig405 vsse 1.35108e-15
C1103 heart_block5_m_16_0_dff_m vsse 5.32008e-16
C1104 heart_block5_ck16 vsse 1.3329e-14
C1105 mbk_sig412 vsse 6.73272e-16
C1106 mbk_sig411 vsse 7.51032e-16
C1107 heart_block5_m_16_0_dff_s vsse 5.89032e-16
C1108 mbk_sig407 vsse 2.26476e-16
C1109 heart_block5_b16 vsse 2.35308e-14
C1110 heart_block5_b016s vsse 2.83954e-15
C1111 heart_block5_s116 vsse 6.68525e-15
C1112 heart_block5_s016 vsse 3.25523e-15
C1113 heart_block5_a16 vsse 9.97223e-15
C1114 heart_block5_oa411s vsse 5.5796e-15
C1115 mbk_sig396 vsse 7.75008e-16
C1116 heart_block5_a115s vsse 4.91443e-15
C1117 heart_block5_a116s vsse 2.1222e-15
C1118 heart_block5_a113s vsse 4.79974e-15
C1119 mbk_sig387 vsse 3.00996e-16
C1120 mbk_sig383 vsse 1.35108e-15
C1121 heart_block5_m_14_2_dff_m vsse 5.32008e-16
C1122 mbk_sig385 vsse 6.73272e-16
C1123 mbk_sig388 vsse 7.51032e-16
C1124 heart_block5_m_14_2_dff_s vsse 5.89032e-16
C1125 heart_block5_s214 vsse 5.69381e-15
C1126 mbk_sig382 vsse 2.26476e-16
C1127 mbk_sig381 vsse 5.51448e-16
C1128 heart_block5_a314s vsse 2.39242e-15
C1129 mbk_sig373 vsse 3.00996e-16
C1130 mbk_sig375 vsse 1.35108e-15
C1131 heart_block5_m_9_0_dff_m vsse 5.32008e-16
C1132 mbk_sig374 vsse 6.73272e-16
C1133 mbk_sig378 vsse 7.51032e-16
C1134 heart_block5_m_9_0_dff_s vsse 5.89032e-16
C1135 mbk_sig370 vsse 2.26476e-16
C1136 heart_block5_oa410s vsse 4.3024e-15
C1137 mbk_sig369 vsse 7.75008e-16
C1138 heart_block5_a016s vsse 4.76993e-15
C1139 heart_block5_a013s vsse 5.27213e-15
C1140 heart_block5_a114s vsse 4.42584e-15
C1141 mbk_sig361 vsse 3.00996e-16
C1142 mbk_sig356 vsse 1.35108e-15
C1143 heart_block5_m_9_1_dff_m vsse 5.32008e-16
C1144 heart_block5_ck9 vsse 1.03119e-14
C1145 mbk_sig358 vsse 6.73272e-16
C1146 mbk_sig362 vsse 7.51032e-16
C1147 heart_block5_m_9_1_dff_s vsse 5.89032e-16
C1148 mbk_sig355 vsse 2.26476e-16
C1149 heart_block5_s215 vsse 4.33415e-15
C1150 heart_block5_a215s vsse 5.33628e-15
C1151 heart_block5_b9 vsse 2.83749e-14
C1152 mbk_sig347 vsse 3.00996e-16
C1153 mbk_sig343 vsse 1.35108e-15
C1154 heart_block5_m_11_1_dff_m vsse 5.32008e-16
C1155 mbk_sig345 vsse 6.73272e-16
C1156 mbk_sig348 vsse 7.51032e-16
C1157 heart_block5_m_11_1_dff_s vsse 5.89032e-16
C1158 mbk_sig342 vsse 2.26476e-16
C1159 heart_block5_ob421s vsse 4.41515e-15
C1160 mbk_sig338 vsse 7.75008e-16
C1161 heart_block5_b19s vsse 3.06569e-15
C1162 mbk_sig332 vsse 7.75008e-16
C1163 heart_a_2 vsse 3.90945e-14
C1164 heart_block5_s211 vsse 9.1483e-15
C1165 heart_block5_na1 vsse 1.46314e-14
C1166 mbk_sig326 vsse 7.75008e-16
C1167 heart_block5_na0 vsse 1.76245e-14
C1168 heart_block5_oa420s vsse 6.26972e-15
C1169 heart_block5_a010s vsse 1.17644e-14
C1170 mbk_sig321 vsse 7.75008e-16
C1171 heart_block5_a011s vsse 1.94011e-15
C1172 heart_block5_s19 vsse 6.15568e-15
C1173 heart_block5_s09 vsse 7.09074e-15
C1174 heart_block5_a09s vsse 2.4961e-15
C1175 heart_a_1 vsse 5.91193e-14
C1176 mbk_sig309 vsse 7.75008e-16
C1177 heart_block5_na2 vsse 1.81174e-14
C1178 heart_a_3 vsse 3.51741e-14
C1179 heart_a_0 vsse 5.89712e-14
C1180 heart_block5_oa421s vsse 5.46685e-15
C1181 mbk_sig303 vsse 7.75008e-16
C1182 heart_block5_a19s vsse 2.82074e-15
C1183 mbk_sig297 vsse 3.00996e-16
C1184 mbk_sig299 vsse 1.35108e-15
C1185 heart_block5_m_12_2_dff_m vsse 5.32008e-16
C1186 mbk_sig298 vsse 6.73272e-16
C1187 mbk_sig302 vsse 7.51032e-16
C1188 heart_block5_m_12_2_dff_s vsse 5.89032e-16
C1189 heart_block5_shram2 vsse 7.16639e-14
C1190 mbk_sig293 vsse 2.26476e-16
C1191 heart_block5_s310 vsse 2.10436e-14
C1192 heart_block5_a310s vsse 3.15252e-15
C1193 heart_block5_b10 vsse 4.97609e-14
C1194 heart_block5_b110s vsse 4.73688e-15
C1195 heart_block5_a012s vsse 3.55298e-15
C1196 heart_block5_s110 vsse 1.00464e-14
C1197 heart_block5_a10 vsse 1.08218e-14
C1198 heart_block5_a110s vsse 2.89397e-15
C1199 heart_block1_ssd0 vsse 2.68013e-15
C1200 heart_d_0 vsse 2.17493e-14
C1201 mbk_sig264 vsse 5.51448e-16
C1202 heart_block1_selas vsse 1.00281e-14
C1203 mbk_sig262 vsse 5.51448e-16
C1204 mbk_sig259 vsse 5.51448e-16
C1205 heart_block1_ni1 vsse 3.48494e-15
C1206 heart_block1_ssa3 vsse 4.12387e-15
C1207 heart_r_3 vsse 5.86181e-15
C1208 mbk_sig257 vsse 5.68296e-16
C1209 mbk_sig256 vsse 5.51448e-16
C1210 ii_2 vsse 9.61843e-15
C1211 heart_d_2 vsse 2.47803e-14
C1212 mbk_sig254 vsse 5.51448e-16
C1213 heart_block1_ssd2 vsse 1.60704e-15
C1214 heart_r_2 vsse 2.54146e-15
C1215 mbk_sig251 vsse 5.68296e-16
C1216 heart_block3_n0 vsse 1.68927e-14
C1217 heart_block3_x01 vsse 1.43692e-14
C1218 mbk_sig247 vsse 7.91856e-16
C1219 heart_block1_o22s vsse 3.40816e-15
C1220 mbk_sig244 vsse 5.68296e-16
C1221 mbk_sig243 vsse 5.51448e-16
C1222 heart_block2_syra2 vsse 1.6861e-15
C1223 heart_block2_syalu2 vsse 4.19256e-15
C1224 yc_2 vsse 2.30048e-14
C1225 mbk_sig241 vsse 5.68296e-16
C1226 ii_1 vsse 9.6889e-15
C1227 mbk_sig239 vsse 5.68296e-16
C1228 heart_block1_ssa2 vsse 3.63787e-15
C1229 mbk_sig238 vsse 5.51448e-16
C1230 heart_block1_ssd3 vsse 4.44334e-15
C1231 heart_d_3 vsse 2.76508e-14
C1232 mbk_sig236 vsse 5.51448e-16
C1233 ii_6 vsse 1.451e-14
C1234 ii_7 vsse 2.76615e-14
C1235 heart_block2_ni6 vsse 2.1964e-15
C1236 heart_block2_selray vsse 1.3441e-14
C1237 mbk_sig234 vsse 6.42492e-16
C1238 heart_block2_ni8 vsse 2.21519e-15
C1239 ii_8 vsse 4.61697e-14
C1240 heart_ra_1 vsse 1.602e-14
C1241 mbk_sig230 vsse 5.51448e-16
C1242 heart_block1_selar vsse 8.56073e-15
C1243 heart_block1_ssa1 vsse 2.29651e-15
C1244 heart_r_1 vsse 4.6818e-15
C1245 mbk_sig228 vsse 5.68296e-16
C1246 heart_block1_ssd1 vsse 2.09693e-15
C1247 heart_d_1 vsse 2.70184e-14
C1248 mbk_sig227 vsse 5.51448e-16
C1249 heart_block1_seldr vsse 9.06034e-15
C1250 heart_block1_selqs vsse 1.47384e-14
C1251 heart_block1_o21s vsse 3.07573e-15
C1252 mbk_sig224 vsse 5.51448e-16
C1253 heart_block1_ni0 vsse 1.87369e-15
C1254 heart_block1_selbs vsse 2.01058e-14
C1255 heart_block1_ni2 vsse 7.6788e-15
C1256 mbk_sig223 vsse 5.51448e-16
C1257 ii_0 vsse 1.04333e-14
C1258 heart_block5_a14 vsse 1.38155e-14
C1259 heart_block5_a014s vsse 5.19761e-15
C1260 heart_block5_b014s vsse 4.58719e-15
C1261 mbk_sig218 vsse 3.00996e-16
C1262 mbk_sig147 vsse 1.35108e-15
C1263 heart_block5_m_14_0_dff_m vsse 5.32008e-16
C1264 mbk_sig219 vsse 6.73272e-16
C1265 mbk_sig149 vsse 7.51032e-16
C1266 heart_block5_m_14_0_dff_s vsse 5.89032e-16
C1267 heart_block5_s014 vsse 2.53984e-15
C1268 mbk_sig217 vsse 2.26476e-16
C1269 mbk_sig216 vsse 3.00996e-16
C1270 mbk_sig143 vsse 1.35108e-15
C1271 heart_block5_m_14_1_dff_m vsse 5.32008e-16
C1272 mbk_sig215 vsse 6.73272e-16
C1273 mbk_sig145 vsse 7.51032e-16
C1274 heart_block5_m_14_1_dff_s vsse 5.89032e-16
C1275 mbk_sig214 vsse 2.26476e-16
C1276 heart_block5_b15 vsse 2.89329e-14
C1277 heart_block5_b015s vsse 5.67842e-15
C1278 heart_block5_b314s vsse 1.0112e-14
C1279 heart_block5_a15 vsse 1.02016e-14
C1280 heart_block5_a015s vsse 2.6244e-15
C1281 heart_block5_oa442s vsse 1.29976e-14
C1282 heart_block5_oa432s vsse 1.01713e-14
C1283 heart_block5_oa412s vsse 6.83154e-15
C1284 heart_ra_2 vsse 9.56205e-15
C1285 mbk_sig210 vsse 3.00996e-16
C1286 mbk_sig125 vsse 1.35108e-15
C1287 heart_block5_m_14_3_dff_m vsse 5.32008e-16
C1288 heart_block5_ck14 vsse 9.02923e-15
C1289 mbk_sig209 vsse 6.73272e-16
C1290 mbk_sig128 vsse 7.51032e-16
C1291 heart_block5_m_14_3_dff_s vsse 5.89032e-16
C1292 heart_block5_s314 vsse 3.93838e-15
C1293 mbk_sig208 vsse 2.26476e-16
C1294 heart_block5_s114 vsse 6.2276e-15
C1295 heart_block5_b14 vsse 2.81323e-14
C1296 heart_block5_b114s vsse 6.03547e-15
C1297 mbk_sig204 vsse 3.00996e-16
C1298 mbk_sig115 vsse 1.35108e-15
C1299 heart_block5_m_15_0_dff_m vsse 5.32008e-16
C1300 heart_block5_ck15 vsse 1.27936e-14
C1301 mbk_sig205 vsse 6.73272e-16
C1302 mbk_sig119 vsse 7.51032e-16
C1303 heart_block5_m_15_0_dff_s vsse 5.89032e-16
C1304 heart_block5_s015 vsse 4.01339e-15
C1305 mbk_sig203 vsse 2.26476e-16
C1306 mbk_sig201 vsse 3.00996e-16
C1307 mbk_sig110 vsse 1.35108e-15
C1308 heart_block5_m_11_0_dff_m vsse 5.32008e-16
C1309 heart_block5_ck11 vsse 1.38975e-14
C1310 mbk_sig202 vsse 6.73272e-16
C1311 mbk_sig113 vsse 7.51032e-16
C1312 heart_block5_m_11_0_dff_s vsse 5.89032e-16
C1313 heart_block5_s011 vsse 5.45778e-15
C1314 mbk_sig200 vsse 2.26476e-16
C1315 heart_block5_b11 vsse 3.64283e-14
C1316 heart_block5_b111s vsse 2.35613e-15
C1317 heart_block5_ob420s vsse 7.56832e-15
C1318 heart_block5_b010s vsse 8.63071e-15
C1319 mbk_sig105 vsse 7.75008e-16
C1320 heart_block5_b011s vsse 3.20371e-15
C1321 heart_block5_b09s vsse 3.54002e-15
C1322 mbk_sig197 vsse 3.00996e-16
C1323 mbk_sig94 vsse 1.35108e-15
C1324 heart_block5_m_12_3_dff_m vsse 5.32008e-16
C1325 mbk_sig198 vsse 6.73272e-16
C1326 mbk_sig97 vsse 7.51032e-16
C1327 heart_block5_m_12_3_dff_s vsse 5.89032e-16
C1328 heart_block5_s312 vsse 7.90998e-15
C1329 heart_block5_shram3 vsse 6.56894e-14
C1330 mbk_sig196 vsse 2.26476e-16
C1331 heart_block5_oa422s vsse 5.09555e-15
C1332 heart_block5_a210s vsse 6.75281e-15
C1333 mbk_sig88 vsse 7.75008e-16
C1334 heart_block5_a211s vsse 2.66911e-15
C1335 heart_block5_s29 vsse 1.13139e-14
C1336 heart_block5_a9 vsse 7.49558e-15
C1337 heart_block5_a29s vsse 1.8954e-15
C1338 mbk_sig193 vsse 3.00996e-16
C1339 mbk_sig79 vsse 1.35108e-15
C1340 heart_block5_m_12_0_dff_m vsse 5.32008e-16
C1341 mbk_sig194 vsse 6.73272e-16
C1342 mbk_sig82 vsse 7.51032e-16
C1343 heart_block5_m_12_0_dff_s vsse 5.89032e-16
C1344 heart_block5_shram0 vsse 5.97446e-14
C1345 mbk_sig192 vsse 2.26476e-16
C1346 heart_block5_s012 vsse 4.8046e-15
C1347 heart_block5_b012s vsse 3.34109e-15
C1348 heart_block5_s111 vsse 5.62772e-15
C1349 heart_block5_a11 vsse 2.10888e-14
C1350 heart_block5_a111s vsse 2.51165e-15
C1351 heart_block5_a112s vsse 2.40408e-15
C1352 heart_block5_b112s vsse 4.41612e-15
C1353 mbk_sig186 vsse 3.00996e-16
C1354 mbk_sig67 vsse 1.35108e-15
C1355 heart_block5_m_12_1_dff_m vsse 5.32008e-16
C1356 mbk_sig187 vsse 6.73272e-16
C1357 mbk_sig69 vsse 7.51032e-16
C1358 heart_block5_m_12_1_dff_s vsse 5.89032e-16
C1359 heart_block5_s112 vsse 2.65648e-15
C1360 heart_block5_shram1 vsse 6.73262e-14
C1361 mbk_sig184 vsse 2.26476e-16
C1362 heart_block5_ck12 vsse 8.1e-15
C1363 heart_block5_enable vsse 7.19909e-14
C1364 mbk_sig183 vsse 5.51448e-16
C1365 heart_block5_b12 vsse 2.53571e-14
C1366 heart_block5_s212 vsse 5.43332e-15
C1367 heart_block5_a12 vsse 7.77632e-15
C1368 vddi vsse 2.56382e-12
C1369 vdde vsse 1.96266e-12
C1370 test vsse 1.48599e-13
C1371 signe vsse 1.80526e-13
C1372 scout vsse 1.80526e-13
C1373 scin vsse 1.48599e-13
C1374 r3 vsse 1.8176e-13
C1375 r0 vsse 1.81761e-13
C1376 q3 vsse 1.81761e-13
C1377 q0 vsse 1.81761e-13
C1378 ovr vsse 1.80526e-13
C1379 np vsse 1.80526e-13
C1380 noe vsse 1.48599e-13
C1381 ng vsse 1.80526e-13
C1382 i_8 vsse 1.48599e-13
C1383 i_7 vsse 1.48599e-13
C1384 i_6 vsse 1.48599e-13
C1385 i_5 vsse 1.48599e-13
C1386 i_4 vsse 1.48599e-13
C1387 i_3 vsse 1.48599e-13
C1388 i_2 vsse 1.48599e-13
C1389 i_1 vsse 1.48599e-13
C1390 i_0 vsse 1.48594e-13
C1391 fonc vsse 1.48599e-13
C1392 d_3 vsse 1.48597e-13
C1393 d_2 vsse 1.48597e-13
C1394 d_1 vsse 1.48597e-13
C1395 d_0 vsse 1.48597e-13
C1396 cout vsse 1.80526e-13
C1397 cke vsse 1.50166e-13
C1398 cin vsse 1.48599e-13
C1399 b_3 vsse 1.48597e-13
C1400 b_2 vsse 1.48597e-13
C1401 b_1 vsse 1.48597e-13
C1402 b_0 vsse 1.48597e-13
C1403 a_3 vsse 1.48597e-13
C1404 a_2 vsse 1.48597e-13
C1405 a_1 vsse 1.48597e-13
C1406 a_0 vsse 1.48597e-13

C1407 heart_block5_a212s vsse 3.71045e-15

.ends cpu2901

