
.subckt ex_m32x32 a_0 a_1 a_2 a_3 a_4 a_5 a_6 a_7 a_8 a_9 a_10 a_11 a_12 a_13 
+ a_14 a_15 a_16 a_17 a_18 a_19 a_20 a_21 a_22 a_23 a_24 a_25 a_26 a_27 a_28 
+ a_29 a_30 a_31 b_0 b_1 b_2 b_3 b_4 b_5 b_6 b_7 b_8 b_9 b_10 b_11 b_12 b_13 
+ b_14 b_15 b_16 b_17 b_18 b_19 b_20 b_21 b_22 b_23 b_24 b_25 b_26 b_27 b_28 
+ b_29 b_30 b_31 p_0 p_1 p_2 p_3 p_4 p_5 p_6 p_7 p_8 p_9 p_10 p_11 p_12 p_13 
+ p_14 p_15 p_16 p_17 p_18 p_19 p_20 p_21 p_22 p_23 p_24 p_25 p_26 p_27 p_28 
+ p_29 p_30 p_31 p_32 p_33 p_34 p_35 p_36 p_37 p_38 p_39 p_40 p_41 p_42 p_43 
+ p_44 p_45 p_46 p_47 p_48 p_49 p_50 p_51 p_52 p_53 p_54 p_55 p_56 p_57 p_58 
+ p_59 p_60 p_61 p_62 p_63 vdd vss 
Mtr_23875 n12163 c_18_1_sum n12084 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23874 n12084 cla_cell0_0_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23873 cla_cell0_0_g n12161 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23872 vdd c_18_1_sum n12161 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23871 n12161 cla_cell0_0_a vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23870 vdd n12161 cla_cell0_0_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23869 vdd n12163 p_30 vdd TP L=0.18U W=1.98U AS=0.7128P AD=0.7128P 
+ PS=4.68U PD=4.68U 
Mtr_23868 n11787 c_18_2_sum n11785 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23867 n11785 c_18_1_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23866 cla_cell0_1_g n11783 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23865 vdd c_18_2_sum n11783 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23864 n11783 c_18_1_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23863 vdd n11783 cla_cell0_1_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23862 vdd n11787 cla_cell0_1_p vdd TP L=0.18U W=1.98U AS=0.7128P 
+ AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23861 vdd n11479 cla_cell0_2_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23860 n11479 c_18_3_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23859 vdd c_18_2_cout n11479 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23858 cla_cell0_2_g n11479 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23857 vdd n11481 cla_cell0_2_p vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23856 cla_cell0_2_pn cla_cell0_2_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23855 n11272 c_18_3_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23854 n11481 c_18_2_cout n11272 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23853 n11059 c_18_4_sum n11273 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23852 n11273 c_18_3_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23851 cla_cell0_3_g n11270 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23850 vdd c_18_4_sum n11270 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23849 n11270 c_18_3_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23848 vdd n11270 cla_cell0_3_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23847 vdd n11059 cla_cell1_3_p1 vdd TP L=0.18U W=1.98U AS=0.7128P 
+ AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23846 n10899 c_18_4_cout n10467 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23845 n10467 c_18_5_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23844 cla_cell0_4_g n10893 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23843 vdd c_18_4_cout n10893 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23842 n10893 c_18_5_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23841 vdd n10893 cla_cell0_4_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23840 vdd n10899 cla_cell3_4_p1 vdd TP L=0.18U W=1.98U AS=0.7128P 
+ AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23839 vdd n10461 cla_cell0_5_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23838 n10461 c_18_5_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23837 vdd c_18_6_sum n10461 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23836 cla_cell0_5_g n10461 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23835 vdd n10465 cla_cell1_5_p1 vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23834 cla_cell7_5_p cla_cell1_5_p1 vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23833 n10466 c_18_5_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23832 n10465 c_18_6_sum n10466 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23831 vdd n10073 cla_cell1_6_tsg vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23830 n10073 c_18_7_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23829 vdd c_18_6_cout n10073 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23828 cla_cell1_6_tsg n10073 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23827 vdd n10079 cla_cell0_6_p vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23826 cla_cell7_6_p cla_cell0_6_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23825 n9636 c_18_7_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23824 n10079 c_18_6_cout n9636 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23823 vdd n9630 cla_cell0_7_g vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_23822 n9630 c_18_7_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23821 vdd c_18_8_sum n9630 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23820 cla_cell0_7_g n9630 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_23819 vdd n9634 cla_cell0_7_p vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_23818 cla_cell0_7_pn cla_cell0_7_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23817 n9635 c_18_7_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23816 n9634 c_18_8_sum n9635 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23815 vdd n9289 cla_cell0_8_g vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_23814 n9289 c_18_9_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23813 vdd c_18_8_cout n9289 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23812 cla_cell0_8_g n9289 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_23811 vdd n9292 cla_cell0_8_p vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_23810 cla_cell7_8_p cla_cell0_8_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23809 n8868 c_18_9_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23808 n9292 c_18_8_cout n8868 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23807 n8869 c_18_10_sum n8867 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23806 n8867 c_18_9_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23805 cla_cell0_9_g n8862 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_23804 vdd c_18_10_sum n8862 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23803 n8862 c_18_9_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23802 vdd n8862 cla_cell0_9_g vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_23801 vdd n8869 cla_cell0_9_p vdd TP L=0.18U W=1.98U AS=0.7128P AD=0.7128P 
+ PS=4.68U PD=4.68U 
Mtr_23800 n8561 c_18_10_cout n8419 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23799 n8419 c_18_11_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23798 cla_cell0_10_g n8557 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23797 vdd c_18_10_cout n8557 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23796 n8557 c_18_11_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23795 vdd n8557 cla_cell0_10_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23794 vdd n8561 cla_cell0_10_p vdd TP L=0.18U W=1.98U AS=0.7128P 
+ AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23793 n8132 c_18_12_sum n8130 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23792 n8130 c_18_11_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23791 cla_cell0_11_g n8126 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23790 vdd c_18_12_sum n8126 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23789 n8126 c_18_11_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23788 vdd n8126 cla_cell0_11_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23787 vdd n8132 cla_cell0_11_p vdd TP L=0.18U W=1.98U AS=0.7128P 
+ AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23786 n7820 c_18_12_cout n7608 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23785 n7608 c_18_13_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23784 cla_cell0_12_g n7815 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23783 vdd c_18_12_cout n7815 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23782 n7815 c_18_13_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23781 vdd n7815 cla_cell0_12_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23780 vdd n7820 cla_cell0_12_p vdd TP L=0.18U W=1.98U AS=0.7128P 
+ AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23779 n7393 c_18_14_sum n7607 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23778 n7607 c_18_13_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23777 cla_cell0_13_g n7604 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23776 vdd c_18_14_sum n7604 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23775 n7604 c_18_13_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23774 vdd n7604 cla_cell0_13_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23773 vdd n7393 cla_cell0_13_p vdd TP L=0.18U W=1.98U AS=0.7128P 
+ AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23772 n7230 c_18_14_cout n6801 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23771 n6801 c_18_15_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23770 cla_cell0_14_g n7059 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23769 vdd c_18_14_cout n7059 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23768 n7059 c_18_15_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23767 vdd n7059 cla_cell0_14_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23766 vdd n7230 cla_cell0_14_p vdd TP L=0.18U W=1.98U AS=0.7128P 
+ AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23765 n6799 c_18_16_sum n6800 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23764 n6800 c_18_15_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23763 cla_cell0_15_g n6795 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23762 vdd c_18_16_sum n6795 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23761 n6795 c_18_15_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23760 vdd n6795 cla_cell0_15_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23759 vdd n6799 cla_cell1_15_p1 vdd TP L=0.18U W=1.98U AS=0.7128P 
+ AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23758 n6419 c_18_16_cout n5954 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23757 n5954 c_18_17_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23756 cla_cell1_16_sg n6415 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23755 vdd c_18_16_cout n6415 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23754 n6415 c_18_17_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23753 vdd n6415 cla_cell1_16_sg vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23752 vdd n6419 cla_cell5_16_p1 vdd TP L=0.18U W=1.98U AS=0.7128P 
+ AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23751 vdd n5946 cla_cell0_17_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23750 n5946 c_18_17_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23749 vdd c_18_18_sum n5946 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23748 cla_cell0_17_g n5946 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23747 vdd n5950 cla_cell0_17_p vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23746 cla_cell0_17_pn cla_cell0_17_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23745 n5951 c_18_17_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23744 n5950 c_18_18_sum n5951 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23743 vdd n5620 cla_cell1_18_tsg vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23742 n5620 c_18_19_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23741 vdd c_18_18_cout n5620 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23740 cla_cell1_18_tsg n5620 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23739 vdd n5625 cla_cell0_18_p vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23738 cla_cell7_18_p cla_cell0_18_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23737 n5182 c_18_19_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23736 n5625 c_18_18_cout n5182 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23735 vdd n5173 cla_cell0_19_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23734 n5173 c_18_19_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23733 vdd c_18_20_sum n5173 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23732 cla_cell0_19_g n5173 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23731 vdd n5180 cla_cell0_19_p vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23730 cla_cell0_19_pn cla_cell0_19_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23729 n5178 c_18_19_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23728 n5180 c_18_20_sum n5178 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23727 vdd n4866 cla_cell0_20_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23726 n4866 c_18_21_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23725 vdd c_18_20_cout n4866 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23724 cla_cell0_20_g n4866 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23723 vdd n4871 cla_cell0_20_p vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23722 cla_cell0_20_pn cla_cell0_20_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23721 n4730 c_18_21_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23720 n4871 c_18_20_cout n4730 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23719 vdd n4437 cla_cell0_21_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23718 n4437 c_18_21_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23717 vdd c_18_22_sum n4437 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23716 cla_cell0_21_g n4437 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23715 vdd n4441 cla_cell0_21_p vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23714 cla_cell0_21_pn cla_cell0_21_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23713 n4442 c_18_21_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23712 n4441 c_18_22_sum n4442 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23711 vdd n4122 cla_cell0_22_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23710 n4122 c_18_23_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23709 vdd c_18_22_cout n4122 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23708 cla_cell0_22_g n4122 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23707 vdd n4126 cla_cell0_22_p vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23706 cla_cell0_22_pn cla_cell0_22_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23705 n3948 c_18_23_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23704 n4126 c_18_22_cout n3948 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23703 vdd n3683 cla_cell0_23_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23702 n3683 c_18_23_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23701 vdd c_18_24_sum n3683 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23700 cla_cell0_23_g n3683 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23699 vdd n3689 cla_cell0_23_p vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23698 cla_cell0_23_pn cla_cell0_23_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23697 n3687 c_18_23_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23696 n3689 c_18_24_sum n3687 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23695 vdd n3349 cla_cell0_24_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23694 n3349 c_18_25_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23693 vdd c_18_24_cout n3349 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23692 cla_cell0_24_g n3349 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23691 vdd n3351 cla_cell0_24_p vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23690 cla_cell0_24_pn cla_cell0_24_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23689 n3098 c_18_25_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23688 n3351 c_18_24_cout n3098 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23687 vdd n3093 cla_cell0_25_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23686 n3093 c_18_25_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23685 vdd c_18_26_sum n3093 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23684 cla_cell0_25_g n3093 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23683 vdd n3097 cla_cell1_25_p1 vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23682 cla_cell0_25_pn cla_cell1_25_p1 vdd vdd TP L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23681 n3099 c_18_25_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23680 n3097 c_18_26_sum n3099 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23679 vdd n2727 cla_cell1_26_tsg vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23678 n2727 c_18_27_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23677 vdd c_18_26_cout n2727 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23676 cla_cell1_26_tsg n2727 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23675 vdd n2732 cla_cell0_26_p vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23674 cla_cell7_26_p cla_cell0_26_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23673 n2265 c_18_27_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23672 n2732 c_18_26_cout n2265 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23671 vdd n2261 cla_cell0_27_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23670 n2261 c_18_27_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23669 vdd c_18_28_sum n2261 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23668 cla_cell0_27_g n2261 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23667 vdd n2266 cla_cell0_27_p vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23666 cla_cell7_27_p cla_cell0_27_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23665 n2267 c_18_27_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23664 n2266 c_18_28_sum n2267 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23663 vdd n1896 cla_cell3_28_g1 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23662 n1896 c_18_29_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23661 vdd c_18_28_cout n1896 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23660 cla_cell3_28_g1 n1896 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23659 vdd n1899 cla_cell0_28_p vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23658 cla_cell7_28_p cla_cell0_28_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23657 n1452 c_18_29_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23656 n1899 c_18_28_cout n1452 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23655 vdd n1447 cla_cell0_29_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23654 n1447 c_18_29_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23653 vdd c_18_30_sum n1447 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23652 cla_cell0_29_g n1447 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23651 vdd n1455 cla_cell0_29_p vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23650 cla_cell0_29_pn cla_cell0_29_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23649 n1451 c_18_29_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23648 n1455 c_18_30_sum n1451 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23647 vdd n1131 cla_cell0_30_g vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23646 n1131 c_18_31_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23645 vdd c_18_30_cout n1131 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23644 cla_cell0_30_g n1131 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23643 vdd n1135 cla_cell0_30_p vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23642 cla_cell0_30_pn cla_cell0_30_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23641 n987 c_18_31_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23640 n1135 c_18_30_cout n987 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23639 vdd n689 cla_cell0_31_g vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_23638 n689 c_18_31_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23637 vdd c_18_32_sum n689 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23636 cla_cell0_31_g n689 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_23635 vdd n694 cla_cell0_31_p vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_23634 cla_cell0_31_pn cla_cell0_31_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23633 n695 c_18_31_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23632 n694 c_18_32_sum n695 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23631 vdd n394 cla_cell0_32_g vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_23630 n394 cla_cell0_32_a vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23629 vdd c_18_32_cout n394 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23628 cla_cell0_32_g n394 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_23627 vdd n398 cla_cell0_32_p vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_23626 cla_cell0_32_pn cla_cell0_32_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23625 n265 cla_cell0_32_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23624 n398 c_18_32_cout n265 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23623 n46 cla_cell0_32_a n44 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23622 n44 cla_cell0_33_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23621 cla_cell0_33_g n41 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_23620 vdd cla_cell0_32_a n41 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23619 n41 cla_cell0_33_a vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23618 vdd n41 cla_cell0_33_g vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_23617 vdd n46 cla_cell0_33_p vdd TP L=0.18U W=1.98U AS=0.7128P AD=0.7128P 
+ PS=4.68U PD=4.68U 
Mtr_23616 vdd cla_cell0_0_g n11781 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_23615 n11781 cla_cell0_1_p vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_23614 cla_cell1_1_co cla_cell0_1_g n11781 vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_23613 vdd cla_cell0_2_g cla_cell1_2_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23612 cla_cell1_2_np cla_cell0_2_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23611 cla_cell1_3_g cla_cell0_3_g n11269 vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23610 n11269 cla_cell0_3_g cla_cell1_3_g vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23609 n11269 cla_cell0_2_g vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23608 n11269 cla_cell0_2_g vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23607 vdd cla_cell1_3_p1 n11269 vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23606 n11054 cla_cell0_2_p vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23605 vdd cla_cell0_2_p n11054 vdd TP L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23604 n11054 cla_cell1_3_p1 vdd vdd TP L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23603 n11054 cla_cell1_3_p1 vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23602 cla_cell2_5_tsg cla_cell0_5_g n10462 vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23601 n10462 cla_cell0_5_g cla_cell2_5_tsg vdd TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23600 n10462 cla_cell0_4_g vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23599 n10462 cla_cell0_4_g vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23598 vdd cla_cell1_5_p1 n10462 vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23597 cla_cell2_5_tsp cla_cell3_4_p1 vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23596 vdd cla_cell3_4_p1 cla_cell2_5_tsp vdd TP L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23595 cla_cell2_5_tsp cla_cell1_5_p1 vdd vdd TP L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23594 cla_cell2_5_tsp cla_cell1_5_p1 vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23593 vdd cla_cell1_6_tsg cla_cell1_6_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23592 cla_cell1_6_np cla_cell0_6_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23591 cla_cell1_7_g cla_cell0_7_g n9632 vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23590 n9632 cla_cell0_7_g cla_cell1_7_g vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23589 n9632 cla_cell1_6_tsg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23588 n9632 cla_cell1_6_tsg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23587 cla_cell2_7_pl cla_cell0_6_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23586 vdd cla_cell0_7_p n9632 vdd TP L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_23585 cla_cell2_7_pl cla_cell0_7_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23584 vdd cla_cell0_8_g cla_cell1_8_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23583 cla_cell1_8_np cla_cell0_8_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23582 cla_cell1_9_g cla_cell0_9_g n8865 vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23581 n8865 cla_cell0_9_g cla_cell1_9_g vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23580 n8865 cla_cell0_8_g vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23579 n8865 cla_cell0_8_g vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_23578 vdd cla_cell0_9_p n8865 vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_23577 cla_cell2_9_sp cla_cell0_8_p vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23576 vdd cla_cell0_8_p cla_cell2_9_sp vdd TP L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23575 cla_cell2_9_sp cla_cell0_9_p vdd vdd TP L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23574 cla_cell2_9_sp cla_cell0_9_p vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23573 vdd cla_cell0_10_g cla_cell1_10_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23572 cla_cell1_10_np cla_cell0_10_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23571 cla_cell1_11_g cla_cell0_11_g n8128 vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23570 n8128 cla_cell0_11_g cla_cell1_11_g vdd TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23569 n8128 cla_cell0_10_g vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23568 n8128 cla_cell0_10_g vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23567 vdd cla_cell0_11_p n8128 vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23566 n8124 cla_cell0_10_p vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23565 vdd cla_cell0_10_p n8124 vdd TP L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23564 n8124 cla_cell0_11_p vdd vdd TP L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23563 n8124 cla_cell0_11_p vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23562 cla_cell1_13_g cla_cell0_13_g n7605 vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23561 n7605 cla_cell0_13_g cla_cell1_13_g vdd TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23560 n7605 cla_cell0_12_g vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23559 n7605 cla_cell0_12_g vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23558 vdd cla_cell0_13_p n7605 vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23557 cla_cell2_13_tsp cla_cell0_12_p vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23556 vdd cla_cell0_12_p cla_cell2_13_tsp vdd TP L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23555 cla_cell2_13_tsp cla_cell0_13_p vdd vdd TP L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23554 cla_cell2_13_tsp cla_cell0_13_p vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23553 vdd cla_cell0_14_g cla_cell1_14_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23552 cla_cell1_14_np cla_cell0_14_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23551 cla_cell2_15_gl cla_cell0_15_g n6796 vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23550 n6796 cla_cell0_15_g cla_cell2_15_gl vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23549 n6796 cla_cell0_14_g vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23548 n6796 cla_cell0_14_g vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23547 cla_cell2_15_pl cla_cell0_14_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23546 vdd cla_cell1_15_p1 n6796 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23545 cla_cell2_15_pl cla_cell1_15_p1 vdd vdd TP L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23544 cla_cell1_17_g cla_cell0_17_g n5948 vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23543 n5948 cla_cell0_17_g cla_cell1_17_g vdd TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23542 n5948 cla_cell1_16_sg vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23541 n5948 cla_cell1_16_sg vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23540 vdd cla_cell0_17_p n5948 vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23539 cla_cell2_17_tsp cla_cell5_16_p1 vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23538 vdd cla_cell5_16_p1 cla_cell2_17_tsp vdd TP L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23537 cla_cell2_17_tsp cla_cell0_17_p vdd vdd TP L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23536 cla_cell2_17_tsp cla_cell0_17_p vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23535 vdd cla_cell1_18_tsg cla_cell1_18_ng vdd TP L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23534 cla_cell1_18_np cla_cell0_18_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23533 cla_cell1_19_g cla_cell0_19_g n5175 vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23532 n5175 cla_cell0_19_g cla_cell1_19_g vdd TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23531 n5175 cla_cell1_18_tsg vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23530 n5175 cla_cell1_18_tsg vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23529 vdd cla_cell0_19_p n5175 vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23528 n5172 cla_cell0_18_p vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23527 vdd cla_cell0_18_p n5172 vdd TP L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23526 n5172 cla_cell0_19_p vdd vdd TP L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23525 n5172 cla_cell0_19_p vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23524 cla_cell1_21_g cla_cell0_21_g n4439 vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23523 n4439 cla_cell0_21_g cla_cell1_21_g vdd TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23522 n4439 cla_cell0_20_g vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23521 n4439 cla_cell0_20_g vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23520 vdd cla_cell0_21_p n4439 vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23519 cla_cell2_21_tsp cla_cell0_20_p vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23518 vdd cla_cell0_20_p cla_cell2_21_tsp vdd TP L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23517 cla_cell2_21_tsp cla_cell0_21_p vdd vdd TP L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23516 cla_cell2_21_tsp cla_cell0_21_p vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23515 vdd cla_cell0_22_g cla_cell1_22_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23514 cla_cell1_22_np cla_cell0_22_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23513 cla_cell1_23_g cla_cell0_23_g n3685 vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23512 n3685 cla_cell0_23_g cla_cell1_23_g vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23511 n3685 cla_cell0_22_g vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23510 n3685 cla_cell0_22_g vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23509 cla_cell2_23_pl cla_cell0_22_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23508 vdd cla_cell0_23_p n3685 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23507 cla_cell2_23_pl cla_cell0_23_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23506 vdd cla_cell0_24_g cla_cell1_24_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23505 cla_cell1_24_np cla_cell0_24_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23504 cla_cell4_25_gl cla_cell0_25_g n3094 vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23503 n3094 cla_cell0_25_g cla_cell4_25_gl vdd TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23502 n3094 cla_cell0_24_g vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23501 n3094 cla_cell0_24_g vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23500 vdd cla_cell1_25_p1 n3094 vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23499 cla_cell2_25_sp cla_cell0_24_p vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23498 vdd cla_cell0_24_p cla_cell2_25_sp vdd TP L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23497 cla_cell2_25_sp cla_cell1_25_p1 vdd vdd TP L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23496 cla_cell2_25_sp cla_cell1_25_p1 vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23495 vdd cla_cell1_26_tsg cla_cell1_26_ng vdd TP L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23494 cla_cell1_26_np cla_cell0_26_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23493 cla_cell1_27_g cla_cell0_27_g n2262 vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23492 n2262 cla_cell0_27_g cla_cell1_27_g vdd TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23491 n2262 cla_cell1_26_tsg vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23490 n2262 cla_cell1_26_tsg vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23489 vdd cla_cell0_27_p n2262 vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23488 n2260 cla_cell0_26_p vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23487 vdd cla_cell0_26_p n2260 vdd TP L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23486 n2260 cla_cell0_27_p vdd vdd TP L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23485 n2260 cla_cell0_27_p vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23484 cla_cell1_29_g cla_cell0_29_g n1449 vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23483 n1449 cla_cell0_29_g cla_cell1_29_g vdd TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23482 n1449 cla_cell3_28_g1 vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23481 n1449 cla_cell3_28_g1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23480 vdd cla_cell0_29_p n1449 vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23479 cla_cell2_29_tsp cla_cell0_28_p vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23478 vdd cla_cell0_28_p cla_cell2_29_tsp vdd TP L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23477 cla_cell2_29_tsp cla_cell0_29_p vdd vdd TP L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23476 cla_cell2_29_tsp cla_cell0_29_p vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23475 vdd cla_cell0_30_g cla_cell1_30_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23474 cla_cell1_30_np cla_cell0_30_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23473 cla_cell1_31_g cla_cell0_31_g n691 vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23472 n691 cla_cell0_31_g cla_cell1_31_g vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23471 n691 cla_cell0_30_g vdd vdd TP L=0.18U W=0.36U AS=0.1296P AD=0.1296P 
+ PS=1.44U PD=1.44U 
Mtr_23470 n691 cla_cell0_30_g vdd vdd TP L=0.18U W=0.36U AS=0.1296P AD=0.1296P 
+ PS=1.44U PD=1.44U 
Mtr_23469 cla_cell2_31_pl cla_cell0_30_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23468 vdd cla_cell0_31_p n691 vdd TP L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_23467 cla_cell2_31_pl cla_cell0_31_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23466 vdd cla_cell0_32_g cla_cell1_32_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23465 cla_cell1_32_np cla_cell0_32_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23464 cla_cell1_33_g cla_cell0_33_g n43 vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23463 n43 cla_cell0_33_g cla_cell1_33_g vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23462 n43 cla_cell0_32_g vdd vdd TP L=0.18U W=0.36U AS=0.1296P AD=0.1296P 
+ PS=1.44U PD=1.44U 
Mtr_23461 n43 cla_cell0_32_g vdd vdd TP L=0.18U W=0.36U AS=0.1296P AD=0.1296P 
+ PS=1.44U PD=1.44U 
Mtr_23460 n39 cla_cell0_32_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P AD=0.2592P 
+ PS=2.16U PD=2.16U 
Mtr_23459 vdd cla_cell0_33_p n43 vdd TP L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_23458 n39 cla_cell0_33_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P AD=0.2592P 
+ PS=2.16U PD=2.16U 
Mtr_23457 vdd cla_cell1_2_ng cla_cell7_2_g vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23456 cla_cell7_2_g cla_cell1_2_np n11268 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23455 n11268 cla_cell1_1_co vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23454 vdd n11054 n11053 vdd TP L=0.18U W=4.5U AS=1.62P AD=1.62P PS=9.72U 
+ PD=9.72U 
Mtr_23453 n11053 cla_cell1_1_co cla_cell3_4_g2 vdd TP L=0.18U W=4.5U AS=1.62P 
+ AD=1.62P PS=9.72U PD=9.72U 
Mtr_23452 cla_cell3_4_g2 cla_cell1_3_g vdd vdd TP L=0.18U W=2.34U AS=0.8424P 
+ AD=0.8424P PS=5.4U PD=5.4U 
Mtr_23451 vdd cla_cell2_5_tsg cla_cell2_5_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23450 cla_cell2_5_np cla_cell2_5_tsp vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23449 n9984 cla_cell1_6_np vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23448 cla_cell3_6_p1 cla_cell2_5_tsp n9984 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23447 vdd cla_cell1_6_np n9627 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23446 n9627 cla_cell2_5_tsg cla_cell2_6_g vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23445 cla_cell2_6_g cla_cell1_6_ng vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23444 n9533 cla_cell2_7_pl vdd vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23443 cla_cell3_7_p1 cla_cell2_5_tsp n9533 vdd TP L=0.18U W=2.52U 
+ AS=0.9072P AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23442 vdd cla_cell2_7_pl n9625 vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23441 n9625 cla_cell2_5_tsg cla_cell2_7_g vdd TP L=0.18U W=2.52U 
+ AS=0.9072P AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23440 cla_cell2_7_g cla_cell1_7_g vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23439 cla_cell2_10_p_s cla_cell2_10_sp vdd vdd TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23438 vdd cla_cell2_10_sg cla_cell2_10_g_s vdd TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23437 vdd n8124 n8546 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_23436 vdd n8553 cla_cell2_10_g1 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23435 vdd n8549 n8551 vdd TP L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_23434 vdd cla_cell2_10_sg cla_cell2_10_g2 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23433 n8121 cla_cell2_10_sp vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23432 cla_cell2_10_sg cla_cell2_10_g_s vdd vdd TP L=0.18U W=1.98U 
+ AS=0.7128P AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23431 cla_cell2_10_sp cla_cell2_10_p_s vdd vdd TP L=0.18U W=1.98U 
+ AS=0.7128P AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23430 n8418 cla_cell1_10_np vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23429 n8549 cla_cell2_9_sp n8418 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23428 vdd cla_cell1_10_np n8417 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23427 n8417 cla_cell1_9_g n8553 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23426 n8553 cla_cell1_10_ng vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23425 vdd cla_cell1_13_g cla_cell2_13_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23424 cla_cell2_13_np cla_cell2_13_tsp vdd vdd TP L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23423 n7055 cla_cell1_14_np vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23422 cla_cell3_14_p1 cla_cell2_13_tsp n7055 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23421 vdd cla_cell1_14_np n6792 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23420 n6792 cla_cell1_13_g cla_cell2_14_g vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23419 cla_cell2_14_g cla_cell1_14_ng vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23418 n6634 cla_cell2_15_pl vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23417 cla_cell3_15_p1 cla_cell2_13_tsp n6634 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23416 vdd cla_cell2_15_pl n6791 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23415 n6791 cla_cell1_13_g cla_cell2_15_g vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23414 cla_cell2_15_g cla_cell2_15_gl vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23413 vdd cla_cell1_17_g cla_cell2_17_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23412 cla_cell2_17_np cla_cell2_17_tsp vdd vdd TP L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23411 cla_cell2_18_g1 cla_cell1_18_ng vdd vdd TP L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23410 n5496 cla_cell1_17_g cla_cell2_18_g1 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23409 vdd cla_cell1_18_np n5496 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23408 cla_cell5_18_p1 cla_cell2_17_tsp n5497 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23407 n5497 cla_cell1_18_np vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23406 cla_cell2_18_sp cla_cell2_18_p_s vdd vdd TP L=0.18U W=1.98U 
+ AS=0.7128P AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23405 cla_cell2_18_sg cla_cell2_18_g_s vdd vdd TP L=0.18U W=1.98U 
+ AS=0.7128P AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23404 vdd n5172 n5611 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_23403 vdd cla_cell2_18_sg cla_cell2_18_g_s vdd TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23402 cla_cell2_18_p_s cla_cell2_18_sp vdd vdd TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23401 vdd cla_cell1_21_g cla_cell2_21_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23400 cla_cell2_21_np cla_cell2_21_tsp vdd vdd TP L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23399 n3946 cla_cell1_22_np vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23398 cla_cell3_22_p11 cla_cell2_21_tsp n3946 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23397 vdd cla_cell1_22_np n3945 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23396 n3945 cla_cell1_21_g cla_cell2_22_g vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23395 cla_cell2_22_g cla_cell1_22_ng vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23394 n3679 cla_cell2_23_pl vdd vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23393 cla_cell3_22_p21 cla_cell2_21_tsp n3679 vdd TP L=0.18U W=2.52U 
+ AS=0.9072P AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23392 vdd cla_cell2_23_pl n3680 vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23391 n3680 cla_cell1_21_g cla_cell2_23_g vdd TP L=0.18U W=2.52U 
+ AS=0.9072P AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23390 cla_cell2_23_g cla_cell1_23_g vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23389 cla_cell2_26_p_s cla_cell2_26_sp vdd vdd TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23388 vdd cla_cell2_26_sg cla_cell2_26_g_s vdd TP L=0.72U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23387 vdd n2260 n2717 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_23386 vdd n2586 cla_cell2_26_g1 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23385 vdd n2718 cla_cell4_26_pl vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23384 vdd cla_cell2_26_sg cla_cell4_27_gl vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23383 cla_cell4_27_pl cla_cell2_26_sp vdd vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23382 cla_cell2_26_sg cla_cell2_26_g_s vdd vdd TP L=0.18U W=1.98U 
+ AS=0.7128P AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23381 cla_cell2_26_sp cla_cell2_26_p_s vdd vdd TP L=0.18U W=1.98U 
+ AS=0.7128P AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23380 n2585 cla_cell1_26_np vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23379 n2718 cla_cell2_25_sp n2585 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23378 vdd cla_cell1_26_np n2258 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23377 n2258 cla_cell4_25_gl n2586 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23376 n2586 cla_cell1_26_ng vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23375 vdd cla_cell1_29_g cla_cell2_29_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23374 cla_cell2_29_np cla_cell2_29_tsp vdd vdd TP L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23373 n985 cla_cell1_30_np vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23372 cla_cell3_30_p1 cla_cell2_29_tsp n985 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23371 vdd cla_cell1_30_np n986 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23370 n986 cla_cell1_29_g cla_cell2_30_g vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23369 cla_cell2_30_g cla_cell1_30_ng vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23368 n686 cla_cell2_31_pl vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23367 cla_cell3_31_p1 cla_cell2_29_tsp n686 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23366 vdd cla_cell2_31_pl n684 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23365 n684 cla_cell1_29_g cla_cell2_31_g vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23364 cla_cell2_31_g cla_cell1_31_g vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23363 vdd cla_cell3_4_g2 n10733 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23362 n10733 cla_cell3_4_p1 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23361 cla_cell3_4_co cla_cell0_4_g n10733 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23360 vdd cla_cell3_4_g2 n10456 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23359 n10456 cla_cell2_5_np vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23358 cla_cell3_5_co cla_cell2_5_ng n10456 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23357 vdd cla_cell3_4_g2 n9983 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23356 n9983 cla_cell3_6_p1 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23355 cla_cell3_6_co cla_cell2_6_g n9983 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23354 n9624 cla_cell4_8_g2 vdd vdd TP L=0.54U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23353 n9532 cla_cell3_7_p1 vdd vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23352 cla_cell4_8_g2 n9624 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_23351 cla_cell3_12_g cla_cell0_12_g n7603 vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23350 n7603 cla_cell0_12_g cla_cell3_12_g vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23349 n7603 cla_cell2_10_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23348 n7603 cla_cell2_10_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23347 n7813 cla_cell2_10_sp vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23346 vdd cla_cell0_12_p n7603 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23345 n7813 cla_cell0_12_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23344 cla_cell3_13_g cla_cell2_13_ng n7386 vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23343 n7386 cla_cell2_13_ng cla_cell3_13_g vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23342 n7386 cla_cell2_10_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23341 n7386 cla_cell2_10_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23340 n7384 cla_cell2_10_sp vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23339 vdd cla_cell2_13_np n7386 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23338 n7384 cla_cell2_13_np vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23337 cla_cell3_14_g cla_cell2_14_g n6788 vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23336 n6788 cla_cell2_14_g cla_cell3_14_g vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23335 n6788 cla_cell2_10_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23334 n6788 cla_cell2_10_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23333 n7052 cla_cell2_10_sp vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23332 vdd cla_cell3_14_p1 n6788 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23331 n7052 cla_cell3_14_p1 vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23330 cla_cell3_15_g cla_cell2_15_g n6787 vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23329 n6787 cla_cell2_15_g cla_cell3_15_g vdd TP L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23328 n6787 cla_cell2_10_sg vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_23327 n6787 cla_cell2_10_sg vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23326 vdd cla_cell3_15_p1 n6787 vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23325 cla_cell4_15_p1 cla_cell2_10_sp vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23324 vdd cla_cell2_10_sp cla_cell4_15_p1 vdd TP L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23323 cla_cell4_15_p1 cla_cell3_15_p1 vdd vdd TP L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_23322 cla_cell4_15_p1 cla_cell3_15_p1 vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_23321 cla_cell3_20_g cla_cell0_20_g n4729 vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23320 n4729 cla_cell0_20_g cla_cell3_20_g vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23319 n4729 cla_cell2_18_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23318 n4729 cla_cell2_18_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23317 cla_cell4_20_p cla_cell2_18_sp vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23316 vdd cla_cell0_20_p n4729 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23315 cla_cell4_20_p cla_cell0_20_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23314 cla_cell3_21_g cla_cell2_21_ng n4432 vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23313 n4432 cla_cell2_21_ng cla_cell3_21_g vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23312 n4432 cla_cell2_18_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23311 n4432 cla_cell2_18_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23310 cla_cell4_21_p cla_cell2_18_sp vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23309 vdd cla_cell2_21_np n4432 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23308 cla_cell4_21_p cla_cell2_21_np vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23307 n4108 cla_cell3_22_sp vdd vdd TP L=0.72U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23306 vdd cla_cell3_22_sg n3676 vdd TP L=0.72U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23305 vdd cla_cell3_22_p21 n4105 vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_23304 n4114 cla_cell3_22_p11 vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23303 vdd n4114 cla_cell5_22_p1 vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_23302 vdd cla_cell3_22_sg cla_cell3_22_g2 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23301 cla_cell5_23_p1 cla_cell3_22_sp vdd vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23300 cla_cell3_22_sg n3676 vdd vdd TP L=0.18U W=1.98U AS=0.7128P 
+ AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23299 vdd n3676 cla_cell3_22_sg vdd TP L=0.18U W=1.98U AS=0.7128P 
+ AD=0.7128P PS=4.68U PD=4.68U 
Mtr_23298 cla_cell3_22_sp n4108 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_23297 vdd cla_cell3_22_p11 n3944 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23296 n4114 cla_cell2_18_sp vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23295 n3944 cla_cell2_18_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23294 n3944 cla_cell2_18_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23293 n3944 cla_cell2_22_g n4112 vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23292 n4112 cla_cell2_22_g n3944 vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23291 vdd n4112 cla_cell3_22_g1 vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_23290 cla_cell3_22_g1 n4112 vdd vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_23289 vdd n4114 cla_cell5_22_p1 vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_23288 cla_cell3_28_g cla_cell3_28_g1 n1771 vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23287 n1771 cla_cell3_28_g1 cla_cell3_28_g vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23286 n1771 cla_cell2_26_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23285 n1771 cla_cell2_26_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23284 cla_cell4_28_pl cla_cell2_26_sp vdd vdd TP L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23283 vdd cla_cell0_28_p n1771 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23282 cla_cell4_28_pl cla_cell0_28_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23281 cla_cell3_29_g cla_cell2_29_ng n1442 vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23280 n1442 cla_cell2_29_ng cla_cell3_29_g vdd TP L=0.18U W=0.36U 
+ AS=0.1296P AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23279 n1442 cla_cell2_26_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23278 n1442 cla_cell2_26_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23277 cla_cell4_29_pl cla_cell2_26_sp vdd vdd TP L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23276 vdd cla_cell2_29_np n1442 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23275 cla_cell4_29_pl cla_cell2_29_np vdd vdd TP L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23274 cla_cell3_30_g cla_cell2_30_g n984 vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23273 n984 cla_cell2_30_g cla_cell3_30_g vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23272 n984 cla_cell2_26_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23271 n984 cla_cell2_26_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23270 cla_cell4_30_pl cla_cell2_26_sp vdd vdd TP L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23269 vdd cla_cell3_30_p1 n984 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23268 cla_cell4_30_pl cla_cell3_30_p1 vdd vdd TP L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23267 cla_cell3_31_g cla_cell2_31_g n683 vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23266 n683 cla_cell2_31_g cla_cell3_31_g vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23265 n683 cla_cell2_26_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23264 n683 cla_cell2_26_sg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23263 cla_cell4_31_pl cla_cell2_26_sp vdd vdd TP L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23262 vdd cla_cell3_31_p1 n683 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23261 cla_cell4_31_pl cla_cell3_31_p1 vdd vdd TP L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23260 vdd cla_cell1_8_ng cla_cell7_8_g vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23259 cla_cell7_8_g cla_cell1_8_np n9183 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23258 n9183 cla_cell4_8_g2 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23257 vdd cla_cell1_9_g cla_cell7_10_co vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23256 cla_cell7_10_co cla_cell2_9_sp n8859 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23255 n8859 cla_cell4_8_g2 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23254 vdd cla_cell2_10_g1 cla_cell7_10_g vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23253 cla_cell7_10_g n8551 n8416 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23252 n8416 cla_cell4_8_g2 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23251 vdd cla_cell2_10_g2 cla_cell7_12_co vdd TP L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23250 cla_cell7_12_co n8121 n8118 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23249 n8118 cla_cell4_8_g2 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23248 vdd cla_cell3_12_g cla_cell7_12_g vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23247 cla_cell7_12_g n7813 n7602 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23246 n7602 cla_cell4_8_g2 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23245 vdd cla_cell3_13_g cla_cell7_14_co vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23244 cla_cell7_14_co n7384 n7382 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23243 n7382 cla_cell4_8_g2 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23242 vdd cla_cell3_14_g cla_cell7_14_g vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23241 cla_cell7_14_g n7052 n6784 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23240 n6784 cla_cell4_8_g2 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23239 vdd n6783 cla_cell5_16_g2 vdd TP L=0.18U W=3.96U AS=1.4256P 
+ AD=1.4256P PS=8.64U PD=8.64U 
Mtr_23238 cla_cell5_16_g2 n6783 vdd vdd TP L=0.18U W=3.96U AS=1.4256P 
+ AD=1.4256P PS=8.64U PD=8.64U 
Mtr_23237 n6632 cla_cell4_15_p1 vdd vdd TP L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_23236 n6783 cla_cell5_16_g2 vdd vdd TP L=0.54U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_23235 vdd cla_cell3_20_g cla_cell4_20_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23234 cla_cell4_20_np cla_cell4_20_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23233 vdd cla_cell3_21_g cla_cell4_21_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23232 cla_cell4_21_np cla_cell4_21_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23231 n3090 cla_cell1_24_np vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23230 cla_cell5_24_p1 cla_cell3_22_sp n3090 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23229 vdd cla_cell1_24_np n3088 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23228 n3088 cla_cell3_22_sg cla_cell4_24_g vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23227 cla_cell4_24_g cla_cell1_24_ng vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23226 n2934 cla_cell2_25_sp vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23225 cla_cell5_25_p1 cla_cell3_22_sp n2934 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23224 vdd cla_cell2_25_sp n2932 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23223 n2932 cla_cell3_22_sg cla_cell4_25_g vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23222 cla_cell4_25_g cla_cell4_25_gl vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23221 n2582 cla_cell4_26_pl vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23220 cla_cell5_26_p1 cla_cell3_22_sp n2582 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23219 vdd cla_cell4_26_pl n2254 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23218 n2254 cla_cell3_22_sg cla_cell4_26_g vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23217 cla_cell4_26_g cla_cell2_26_g1 vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23216 n2130 cla_cell4_27_pl vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23215 cla_cell5_27_p1 cla_cell3_22_sp n2130 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23214 vdd cla_cell4_27_pl n2253 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23213 n2253 cla_cell3_22_sg cla_cell4_27_g vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23212 cla_cell4_27_g cla_cell4_27_gl vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23211 n1770 cla_cell4_28_pl vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23210 cla_cell5_28_p1 cla_cell3_22_sp n1770 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23209 vdd cla_cell4_28_pl n1769 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23208 n1769 cla_cell3_22_sg cla_cell4_28_g vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23207 cla_cell4_28_g cla_cell3_28_g vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23206 n1439 cla_cell4_29_pl vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23205 cla_cell5_29_p1 cla_cell3_22_sp n1439 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23204 vdd cla_cell4_29_pl n1437 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23203 n1437 cla_cell3_22_sg cla_cell4_29_g vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23202 cla_cell4_29_g cla_cell3_29_g vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23201 n982 cla_cell4_30_pl vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23200 cla_cell5_30_p1 cla_cell3_22_sp n982 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23199 vdd cla_cell4_30_pl n983 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23198 n983 cla_cell3_22_sg cla_cell4_30_g vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23197 cla_cell4_30_g cla_cell3_30_g vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23196 n680 cla_cell4_31_pl vdd vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23195 n678 cla_cell3_22_sp n680 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23194 vdd cla_cell4_31_pl n677 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23193 n677 cla_cell3_22_sg cla_cell4_31_g vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_23192 cla_cell4_31_g cla_cell3_31_g vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_23191 vdd cla_cell5_16_g2 n6298 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23190 n6298 cla_cell5_16_p1 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23189 cla_cell5_16_co cla_cell1_16_sg n6298 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23188 vdd cla_cell5_16_g2 n5941 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23187 n5941 cla_cell2_17_np vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23186 cla_cell5_17_co cla_cell2_17_ng n5941 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23185 vdd cla_cell5_16_g2 n5495 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23184 n5495 cla_cell5_18_p1 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23183 cla_cell5_18_co cla_cell2_18_g1 n5495 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23182 vdd cla_cell5_16_g2 n5169 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23181 n5169 cla_cell2_18_sp vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23180 cla_cell5_19_co cla_cell2_18_sg n5169 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23179 vdd cla_cell5_16_g2 n4728 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23178 n4728 cla_cell4_20_np vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23177 cla_cell5_20_co cla_cell4_20_ng n4728 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23176 vdd cla_cell5_16_g2 n4427 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23175 n4427 cla_cell4_21_np vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23174 cla_cell5_21_co cla_cell4_21_ng n4427 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23173 vdd cla_cell5_16_g2 n3943 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23172 n3943 cla_cell5_22_p1 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23171 cla_cell5_22_co cla_cell3_22_g1 n3943 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23170 vdd cla_cell5_16_g2 n3673 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23169 n3673 cla_cell5_23_p1 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23168 cla_cell5_23_co cla_cell3_22_g2 n3673 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23167 vdd cla_cell5_16_g2 n3086 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23166 n3086 cla_cell5_24_p1 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23165 cla_cell5_24_co cla_cell4_24_g n3086 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23164 vdd cla_cell5_16_g2 n3085 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23163 n3085 cla_cell5_25_p1 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23162 cla_cell5_25_co cla_cell4_25_g n3085 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23161 vdd cla_cell5_16_g2 n2581 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23160 n2581 cla_cell5_26_p1 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23159 cla_cell5_26_co cla_cell4_26_g n2581 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23158 vdd cla_cell5_16_g2 n2251 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23157 n2251 cla_cell5_27_p1 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23156 cla_cell5_27_co cla_cell4_27_g n2251 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23155 vdd cla_cell5_16_g2 n1768 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23154 n1768 cla_cell5_28_p1 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23153 cla_cell5_28_co cla_cell4_28_g n1768 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23152 vdd cla_cell5_16_g2 n1436 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23151 n1436 cla_cell5_29_p1 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23150 cla_cell5_29_co cla_cell4_29_g n1436 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23149 vdd cla_cell5_16_g2 n981 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23148 n981 cla_cell5_30_p1 vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23147 cla_cell5_30_co cla_cell4_30_g n981 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23146 vdd cla_cell5_16_g2 n676 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_23145 n676 n678 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23144 cla_cell5_31_co cla_cell4_31_g n676 vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_23143 vdd cla_cell1_32_ng cla_cell7_32_g vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_23142 cla_cell7_32_g cla_cell1_32_np n264 vdd TP L=0.18U W=2.88U 
+ AS=1.0368P AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23141 n264 cla_cell5_31_co vdd vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_23140 vdd cla_cell1_33_g n38 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23139 n38 n39 n37 vdd TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P PS=6.48U 
+ PD=6.48U 
Mtr_23138 n37 cla_cell5_31_co vdd vdd TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_23137 n11779 cla_cell0_1_p n11778 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23136 n11778 cla_cell0_0_g vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23135 p_31 n11779 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23134 n11266 cla_cell1_1_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23133 n11473 cla_cell0_2_pn n11266 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23132 p_32 n11473 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23131 n11265 cla_cell1_3_p1 n11052 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23130 n11052 cla_cell7_2_g vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23129 p_33 n11265 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23128 n10455 cla_cell3_4_g2 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23127 n10887 cla_cell3_4_p1 n10455 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23126 p_34 n10887 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23125 n10453 cla_cell7_5_p n10454 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23124 n10454 cla_cell3_4_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23123 p_35 n10453 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23122 n9621 cla_cell3_5_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23121 n10061 cla_cell7_6_p n9621 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23120 p_36 n10061 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23119 n9619 cla_cell0_7_pn n9620 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23118 n9620 cla_cell3_6_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23117 p_37 n9619 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23116 n9182 cla_cell4_8_g2 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23115 n9280 cla_cell7_8_p n9182 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23114 p_38 n9280 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23113 n8857 cla_cell0_9_p n8858 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23112 n8858 cla_cell7_8_g vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_23111 p_39 n8857 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23110 n8415 cla_cell7_10_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23109 n8543 cla_cell0_10_p n8415 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23108 p_40 n8543 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23107 n8117 cla_cell0_11_p n8116 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23106 n8116 cla_cell7_10_g vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23105 p_41 n8117 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23104 n7601 cla_cell7_12_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23103 n7808 cla_cell0_12_p n7601 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23102 p_42 n7808 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23101 n7600 cla_cell0_13_p n7381 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23100 n7381 cla_cell7_12_g vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23099 p_43 n7600 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23098 n6781 cla_cell7_14_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23097 n7216 cla_cell0_14_p n6781 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23096 p_44 n7216 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23095 n6779 cla_cell1_15_p1 n6780 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23094 n6780 cla_cell7_14_g vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23093 p_45 n6779 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23092 n5940 cla_cell5_16_g2 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23091 n6405 cla_cell5_16_p1 n5940 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23090 p_46 n6405 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23089 n5938 cla_cell0_17_pn n5939 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23088 n5939 cla_cell5_16_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23087 p_47 n5938 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23086 n5167 cla_cell5_17_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23085 n5606 cla_cell7_18_p n5167 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23084 p_48 n5606 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23083 n5165 cla_cell0_19_pn n5166 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23082 n5166 cla_cell5_18_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23081 p_49 n5165 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23080 n4727 cla_cell5_19_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23079 n4854 cla_cell0_20_pn n4727 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23078 p_50 n4854 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23077 n4425 cla_cell0_21_pn n4424 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23076 n4424 cla_cell5_20_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23075 p_51 n4425 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23074 n3942 cla_cell5_21_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23073 n4102 cla_cell0_22_pn n3942 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23072 p_52 n4102 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23071 n3671 cla_cell0_23_pn n3670 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23070 n3670 cla_cell5_22_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23069 p_53 n3671 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23068 n3084 cla_cell5_23_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23067 n3523 cla_cell0_24_pn n3084 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23066 p_54 n3523 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23065 n3082 cla_cell0_25_pn n3083 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23064 n3083 cla_cell5_24_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23063 p_55 n3082 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23062 n2249 cla_cell5_25_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23061 n2710 cla_cell7_26_p n2249 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23060 p_56 n2710 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23059 n2247 cla_cell7_27_p n2248 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23058 n2248 cla_cell5_26_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23057 p_57 n2247 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23056 n1434 cla_cell5_27_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23055 n1880 cla_cell7_28_p n1434 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23054 p_58 n1880 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23053 n1432 cla_cell0_29_pn n1433 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23052 n1433 cla_cell5_28_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23051 p_59 n1432 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23050 n980 cla_cell5_29_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23049 n1111 cla_cell0_30_pn n980 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23048 p_60 n1111 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23047 n673 cla_cell0_31_pn n674 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23046 n674 cla_cell5_30_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23045 p_61 n673 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23044 n263 cla_cell5_31_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23043 n387 cla_cell0_32_pn n263 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_23042 p_62 n387 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23041 n36 cla_cell0_33_p n35 vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_23040 n35 cla_cell7_32_g vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_23039 p_63 n36 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_23038 cla_cell0_32_a n54 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23037 n52 n51 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_23036 cla_cell0_33_a n55 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_23035 n48 c_18_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_23034 vdd p_18_33_pi2j n48 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23033 n55 c_18_32_cin n48 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23032 n55 c_18_31_a n53 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_23031 n53 p_18_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23030 n54 c_18_32_cin n52 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23029 vdd n50 n51 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P PS=3.6U 
+ PD=3.6U 
Mtr_23028 n50 c_18_31_a n49 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_23027 n49 p_18_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23026 n61 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_23025 vdd p_18_33_t_s n57 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_23024 n57 p_18_1_n2j p_18_33_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23023 vdd n61 n58 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_23022 n58 n59 p_18_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_23021 n59 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_23020 vdd n409 n271 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_23019 n270 p_18_1_n2j p_18_32_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_23018 vdd p_18_32_t_s n270 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_23017 vdd a_30 n272 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_23016 n273 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_23015 n412 p_18_2_d2j n273 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_23014 n272 p_18_2_d2jbar n412 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_23013 n409 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_23012 n271 n412 p_18_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_23011 vdd c_18_31_a n266 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23010 c_18_32_sum c_18_32_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_23009 n269 n404 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_23008 c_18_32_cout n402 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_23007 n266 p_18_32_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23006 n402 c_18_32_cin n266 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23005 n402 p_18_32_pi2j n268 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23004 n268 c_18_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_23003 c_18_32_s2_s c_18_32_cin n269 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_23002 vdd c_18_32_s1_s n404 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_23001 c_18_32_s1_s p_18_32_pi2j n267 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_23000 n267 c_18_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22999 c_18_31_sum c_18_31_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22998 n705 n704 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22997 c_18_31_cout n707 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22996 n699 c_18_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22995 vdd p_18_31_pi2j n699 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22994 n707 c_18_31_cin n699 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22993 n707 c_18_31_a n706 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22992 n706 p_18_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22991 c_18_31_s2_s c_18_31_cin n705 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22990 vdd c_18_31_s1_s n704 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22989 c_18_31_s1_s c_18_31_a n702 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22988 n702 p_18_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22987 n714 p_18_2_d2j n715 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22986 n715 p_18_2_d2jbar n716 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22985 n716 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22984 vdd a_30 n714 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22983 vdd p_18_31_t_s n710 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22982 n710 p_18_1_n2j p_18_31_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22981 vdd n715 n711 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22980 n711 n713 p_18_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22979 n713 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22978 vdd n1148 n993 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22977 n992 p_18_1_n2j p_18_30_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22976 vdd p_18_30_t_s n992 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22975 vdd a_28 n994 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22974 n995 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22973 n1150 p_18_2_d2j n995 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22972 n994 p_18_2_d2jbar n1150 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22971 n1148 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22970 n993 n1150 p_18_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22969 vdd c_18_30_a n988 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22968 c_18_30_sum c_18_30_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22967 n990 n1142 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22966 c_18_30_cout n1140 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22965 n988 p_18_30_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22964 n1140 c_18_30_cin n988 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22963 n1140 p_18_30_pi2j n991 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22962 n991 c_18_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22961 c_18_30_s2_s c_18_30_cin n990 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22960 vdd c_18_30_s1_s n1142 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22959 c_18_30_s1_s p_18_30_pi2j n989 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22958 n989 c_18_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22957 c_18_29_sum c_18_29_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22956 n1466 n1462 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22955 c_18_29_cout n1467 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22954 n1456 c_18_29_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22953 vdd p_18_29_pi2j n1456 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22952 n1467 c_18_29_cin n1456 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22951 n1467 c_18_29_a n1465 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22950 n1465 p_18_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22949 c_18_29_s2_s c_18_29_cin n1466 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22948 vdd c_18_29_s1_s n1462 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22947 c_18_29_s1_s c_18_29_a n1463 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22946 n1463 p_18_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22945 n1474 p_18_2_d2j n1475 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22944 n1475 p_18_2_d2jbar n1476 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22943 n1476 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22942 vdd a_28 n1474 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22941 vdd p_18_29_t_s n1470 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22940 n1470 p_18_1_n2j p_18_29_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22939 vdd n1475 n1471 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22938 n1471 n1473 p_18_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22937 n1473 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22936 vdd n1911 n1776 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22935 n1775 p_18_1_n2j p_18_28_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22934 vdd p_18_28_t_s n1775 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22933 vdd a_26 n1777 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22932 n1778 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22931 n1913 p_18_2_d2j n1778 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22930 n1777 p_18_2_d2jbar n1913 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22929 n1911 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22928 n1776 n1913 p_18_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22927 vdd c_18_28_a n1772 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22926 c_18_28_sum c_18_28_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22925 n1773 n1774 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22924 c_18_28_cout n1902 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22923 n1772 p_18_28_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22922 n1902 c_18_28_cin n1772 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22921 n1902 p_18_28_pi2j n1461 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22920 n1461 c_18_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22919 c_18_28_s2_s c_18_28_cin n1773 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22918 vdd c_18_28_s1_s n1774 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22917 c_18_28_s1_s p_18_28_pi2j n1460 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22916 n1460 c_18_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22915 c_18_27_sum c_18_27_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22914 n2135 n2272 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22913 c_18_27_cout n2279 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22912 n2269 c_18_27_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22911 vdd c_18_27_b n2269 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22910 n2279 c_18_27_cin n2269 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22909 n2279 c_18_27_a n2277 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22908 n2277 c_18_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22907 c_18_27_s2_s c_18_27_cin n2135 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22906 vdd c_18_27_s1_s n2272 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22905 c_18_27_s1_s c_18_27_a n2276 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22904 n2276 c_18_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22903 n2137 p_18_2_d2j n2280 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22902 n2280 p_18_2_d2jbar n2139 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22901 n2139 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22900 vdd a_26 n2137 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22899 vdd p_18_27_t_s n2136 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22898 n2136 p_18_1_n2j c_18_27_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22897 vdd n2280 n2286 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22896 n2286 n2283 p_18_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22895 n2283 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22894 vdd n2593 n2284 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22893 n2282 p_18_1_n2j p_18_26_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22892 vdd p_18_26_t_s n2282 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22891 vdd a_24 n2287 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22890 n2288 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22889 n2595 p_18_2_d2j n2288 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22888 n2287 p_18_2_d2jbar n2595 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22887 n2593 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22886 n2284 n2595 p_18_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22885 vdd c_18_26_a n2588 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22884 c_18_26_sum c_18_26_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22883 n2590 n2591 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22882 c_18_26_cout n2736 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22881 n2588 p_18_26_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22880 n2736 c_18_26_cin n2588 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22879 n2736 p_18_26_pi2j n2275 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22878 n2275 c_18_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22877 c_18_26_s2_s c_18_26_cin n2590 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22876 vdd c_18_26_s1_s n2591 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22875 c_18_26_s1_s p_18_26_pi2j n2274 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22874 n2274 c_18_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22873 c_18_25_sum c_18_25_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22872 n2937 n2939 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22871 c_18_25_cout n3107 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22870 n3101 c_18_25_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22869 vdd c_18_25_b n3101 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22868 n3107 c_18_25_cin n3101 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22867 n3107 c_18_25_a n3108 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22866 n3108 c_18_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22865 c_18_25_s2_s c_18_25_cin n2937 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22864 vdd c_18_25_s1_s n2939 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22863 c_18_25_s1_s c_18_25_a n3106 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22862 n3106 c_18_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22861 n2943 p_18_2_d2j n2944 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22860 n2944 p_18_2_d2jbar n2945 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22859 n2945 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22858 vdd a_24 n2943 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22857 vdd p_18_25_t_s n2941 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22856 n2941 p_18_1_n2j c_18_25_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22855 vdd n2944 n2942 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22854 n2942 n3112 p_18_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22853 n3112 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22852 vdd n3361 n3113 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22851 n3110 p_18_1_n2j c_18_24_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22850 vdd p_18_24_t_s n3110 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22849 vdd a_22 n3114 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22848 n3115 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22847 n3362 p_18_2_d2j n3115 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22846 n3114 p_18_2_d2jbar n3362 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22845 n3361 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22844 n3113 n3362 p_18_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22843 vdd c_18_24_a n3100 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22842 c_18_24_sum c_18_24_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22841 n3355 n3356 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22840 c_18_24_cout n3353 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22839 n3100 c_18_24_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22838 n3353 c_18_24_cin n3100 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22837 n3353 c_18_24_b n3104 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22836 n3104 c_18_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22835 c_18_24_s2_s c_18_24_cin n3355 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22834 vdd c_18_24_s1_s n3356 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22833 c_18_24_s1_s c_18_24_b n3103 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22832 n3103 c_18_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22831 c_18_23_sum c_18_23_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22830 n3695 n3699 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22829 c_18_23_cout n3697 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22828 n3949 c_18_23_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22827 vdd c_18_23_b n3949 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22826 n3697 c_18_23_cin n3949 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22825 n3697 c_18_23_a n3694 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22824 n3694 c_18_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22823 c_18_23_s2_s c_18_23_cin n3695 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22822 vdd c_18_23_s1_s n3699 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22821 c_18_23_s1_s c_18_23_a n3692 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22820 n3692 c_18_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22819 n3704 p_18_2_d2j n3705 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22818 n3705 p_18_2_d2jbar n3706 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22817 n3706 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22816 vdd a_22 n3704 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22815 vdd p_18_23_t_s n3700 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22814 n3700 p_18_1_n2j c_18_23_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22813 vdd n3705 n3701 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22812 n3701 n3703 p_18_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22811 n3703 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22810 vdd n4139 n3956 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22809 n3955 p_18_1_n2j p_18_22_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22808 vdd p_18_22_t_s n3955 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22807 vdd a_20 n3957 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22806 n3958 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22805 n4141 p_18_2_d2j n3958 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22804 n3957 p_18_2_d2jbar n4141 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22803 n4139 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22802 n3956 n4141 p_18_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22801 vdd c_18_22_a n3950 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22800 c_18_22_sum c_18_22_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22799 n3952 n4132 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22798 c_18_22_cout n4130 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22797 n3950 p_18_22_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22796 n4130 c_18_22_cin n3950 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22795 n4130 p_18_22_pi2j n3953 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22794 n3953 c_18_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22793 c_18_22_s2_s c_18_22_cin n3952 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22792 vdd c_18_22_s1_s n4132 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22791 c_18_22_s1_s p_18_22_pi2j n3951 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22790 n3951 c_18_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22789 c_18_21_sum c_18_21_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22788 n4454 n4449 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22787 c_18_21_cout n4453 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22786 n4446 c_18_21_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22785 vdd p_18_21_pi2j n4446 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22784 n4453 c_18_21_cin n4446 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22783 n4453 c_18_21_a n4451 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22782 n4451 p_18_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22781 c_18_21_s2_s c_18_21_cin n4454 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22780 vdd c_18_21_s1_s n4449 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22779 c_18_21_s1_s c_18_21_a n4450 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22778 n4450 p_18_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22777 n4461 p_18_2_d2j n4462 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22776 n4462 p_18_2_d2jbar n4463 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22775 n4463 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22774 vdd a_20 n4461 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22773 vdd p_18_21_t_s n4457 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22772 n4457 p_18_1_n2j p_18_21_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22771 vdd n4462 n4458 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22770 n4458 n4460 p_18_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22769 n4460 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22768 vdd n4885 n4736 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22767 n4735 p_18_1_n2j p_18_20_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22766 vdd p_18_20_t_s n4735 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22765 vdd a_18 n4737 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22764 n4738 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22763 n4886 p_18_2_d2j n4738 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22762 n4737 p_18_2_d2jbar n4886 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22761 n4885 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22760 n4736 n4886 p_18_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22759 vdd c_18_20_a n4731 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22758 c_18_20_sum c_18_20_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22757 n4733 n4878 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22756 c_18_20_cout n4876 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22755 n4731 p_18_20_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22754 n4876 c_18_20_cin n4731 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22753 n4876 p_18_20_pi2j n4734 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22752 n4734 c_18_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22751 c_18_20_s2_s c_18_20_cin n4733 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22750 vdd c_18_20_s1_s n4878 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22749 c_18_20_s1_s p_18_20_pi2j n4732 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22748 n4732 c_18_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22747 c_18_19_sum c_18_19_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22746 n5194 n5189 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22745 c_18_19_cout n5193 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22744 n5184 c_18_19_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22743 vdd p_18_19_pi2j n5184 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22742 n5193 c_18_19_cin n5184 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22741 n5193 c_18_19_a n5191 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22740 n5191 p_18_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22739 c_18_19_s2_s c_18_19_cin n5194 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22738 vdd c_18_19_s1_s n5189 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22737 c_18_19_s1_s c_18_19_a n5190 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22736 n5190 p_18_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22735 n5201 p_18_2_d2j n5203 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22734 n5203 p_18_2_d2jbar n5202 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22733 n5202 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22732 vdd a_18 n5201 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22731 vdd p_18_19_t_s n5197 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22730 n5197 p_18_1_n2j p_18_19_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22729 vdd n5203 n5198 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22728 n5198 n5200 p_18_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22727 n5200 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22726 vdd n5637 n5502 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22725 n5501 p_18_1_n2j p_18_18_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22724 vdd p_18_18_t_s n5501 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22723 vdd a_16 n5503 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22722 n5504 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22721 n5640 p_18_2_d2j n5504 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22720 n5503 p_18_2_d2jbar n5640 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22719 n5637 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22718 n5502 n5640 p_18_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22717 vdd c_18_18_a n5498 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22716 c_18_18_sum c_18_18_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22715 n5499 n5500 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22714 c_18_18_cout n5628 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22713 n5498 p_18_18_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22712 n5628 c_18_18_cin n5498 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22711 n5628 p_18_18_pi2j n5188 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22710 n5188 c_18_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22709 c_18_18_s2_s c_18_18_cin n5499 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22708 vdd c_18_18_s1_s n5500 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22707 c_18_18_s1_s p_18_18_pi2j n5187 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22706 n5187 c_18_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22705 c_18_17_sum c_18_17_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22704 n5965 n5958 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22703 c_18_17_cout n5964 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22702 n5955 c_18_17_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22701 vdd p_18_17_pi2j n5955 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22700 n5964 c_18_17_cin n5955 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22699 n5964 c_18_17_a n5966 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22698 n5966 p_18_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22697 c_18_17_s2_s c_18_17_cin n5965 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22696 vdd c_18_17_s1_s n5958 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22695 c_18_17_s1_s c_18_17_a n5963 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22694 n5963 p_18_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22693 n5858 p_18_2_d2j n5968 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22692 n5968 p_18_2_d2jbar n5860 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22691 n5860 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22690 vdd a_16 n5858 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22689 vdd p_18_17_t_s n5970 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22688 n5970 p_18_1_n2j p_18_17_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22687 vdd n5968 n5975 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22686 n5975 n5972 p_18_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22685 n5972 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22684 vdd n6429 n5973 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22683 n5969 p_18_1_n2j p_18_16_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22682 vdd p_18_16_t_s n5969 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22681 vdd a_14 n5976 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22680 n5977 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22679 n6305 p_18_2_d2j n5977 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22678 n5976 p_18_2_d2jbar n6305 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22677 n6429 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22676 n5973 n6305 p_18_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22675 vdd c_18_16_a n6299 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22674 c_18_16_sum c_18_16_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22673 n6301 n6302 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22672 c_18_16_cout n6423 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22671 n6299 p_18_16_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22670 n6423 c_18_16_cin n6299 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22669 n6423 p_18_16_pi2j n5961 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22668 n5961 c_18_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22667 c_18_16_s2_s c_18_16_cin n6301 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22666 vdd c_18_16_s1_s n6302 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22665 c_18_16_s1_s p_18_16_pi2j n5960 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22664 n5960 c_18_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22663 c_18_15_sum c_18_15_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22662 n6638 n6640 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22661 c_18_15_cout n6810 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22660 n6803 c_18_15_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22659 vdd c_18_15_b n6803 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22658 n6810 c_18_15_cin n6803 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22657 n6810 c_18_15_a n6807 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22656 n6807 c_18_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22655 c_18_15_s2_s c_18_15_cin n6638 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22654 vdd c_18_15_s1_s n6640 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22653 c_18_15_s1_s c_18_15_a n6809 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22652 n6809 c_18_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22651 n6644 p_18_2_d2j n6645 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22650 n6645 p_18_2_d2jbar n6646 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22649 n6646 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22648 vdd a_14 n6644 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22647 vdd p_18_15_t_s n6642 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22646 n6642 p_18_1_n2j c_18_15_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22645 vdd n6645 n6643 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22644 n6643 n6814 p_18_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22643 n6814 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22642 vdd n7068 n6815 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22641 n6812 p_18_1_n2j p_18_14_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22640 vdd p_18_14_t_s n6812 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22639 vdd a_12 n6816 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22638 n6817 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22637 n7069 p_18_2_d2j n6817 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22636 n6816 p_18_2_d2jbar n7069 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22635 n7068 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22634 n6815 n7069 p_18_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22633 vdd c_18_14_a n6802 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22632 c_18_14_sum c_18_14_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22631 n7063 n7064 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22630 c_18_14_cout n7061 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22629 n6802 p_18_14_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22628 n7061 c_18_14_cin n6802 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22627 n7061 p_18_14_pi2j n6806 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22626 n6806 c_18_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22625 c_18_14_s2_s c_18_14_cin n7063 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22624 vdd c_18_14_s1_s n7064 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22623 c_18_14_s1_s p_18_14_pi2j n6805 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22622 n6805 c_18_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22621 c_18_13_sum c_18_13_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22620 n7396 n7400 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22619 c_18_13_cout n7397 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22618 n7609 c_18_13_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22617 vdd c_18_13_b n7609 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22616 n7397 c_18_13_cin n7609 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22615 n7397 c_18_13_a n7614 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22614 n7614 c_18_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22613 c_18_13_s2_s c_18_13_cin n7396 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22612 vdd c_18_13_s1_s n7400 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22611 c_18_13_s1_s c_18_13_a n7615 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22610 n7615 c_18_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22609 n7405 p_18_2_d2j n7406 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22608 n7406 p_18_2_d2jbar n7407 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22607 n7407 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22606 vdd a_12 n7405 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22605 vdd p_18_13_t_s n7402 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22604 n7402 p_18_1_n2j c_18_13_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22603 vdd n7406 n7403 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22602 n7403 n7404 p_18_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22601 n7404 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22600 vdd n7832 n7619 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22599 n7617 p_18_1_n2j c_18_12_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22598 vdd p_18_12_t_s n7617 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22597 vdd a_10 n7620 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22596 n7621 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22595 n7834 p_18_2_d2j n7621 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22594 n7620 p_18_2_d2jbar n7834 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22593 n7832 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22592 n7619 n7834 p_18_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22591 vdd c_18_12_a n7610 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22590 c_18_12_sum c_18_12_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22589 n7612 n7826 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22588 c_18_12_cout n7824 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22587 n7610 c_18_12_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22586 n7824 c_18_12_cin n7610 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22585 n7824 c_18_12_b n7613 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22584 n7613 c_18_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22583 c_18_12_s2_s c_18_12_cin n7612 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22582 vdd c_18_12_s1_s n7826 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22581 c_18_12_s1_s c_18_12_b n7611 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22580 n7611 c_18_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22579 c_18_11_sum c_18_11_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22578 n8141 n8137 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22577 c_18_11_cout n8142 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22576 n8134 c_18_11_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22575 vdd p_18_11_pi2j n8134 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22574 n8142 c_18_11_cin n8134 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22573 n8142 c_18_11_a n8140 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22572 n8140 p_18_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22571 c_18_11_s2_s c_18_11_cin n8141 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22570 vdd c_18_11_s1_s n8137 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22569 c_18_11_s1_s c_18_11_a n8138 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22568 n8138 p_18_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22567 n8149 p_18_2_d2j n8150 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22566 n8150 p_18_2_d2jbar n8151 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22565 n8151 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22564 vdd a_10 n8149 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22563 vdd p_18_11_t_s n8145 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22562 n8145 p_18_1_n2j p_18_11_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22561 vdd n8150 n8146 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22560 n8146 n8148 p_18_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22559 n8148 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22558 vdd n8574 n8425 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22557 n8424 p_18_1_n2j p_18_10_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22556 vdd p_18_10_t_s n8424 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22555 vdd a_8 n8426 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22554 n8427 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22553 n8575 p_18_2_d2j n8427 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22552 n8426 p_18_2_d2jbar n8575 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22551 n8574 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22550 n8425 n8575 p_18_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22549 vdd c_18_10_a n8420 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22548 c_18_10_sum c_18_10_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22547 n8422 n8567 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22546 c_18_10_cout n8562 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22545 n8420 p_18_10_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22544 n8562 c_18_10_cin n8420 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22543 n8562 p_18_10_pi2j n8423 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22542 n8423 c_18_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22541 c_18_10_s2_s c_18_10_cin n8422 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22540 vdd c_18_10_s1_s n8567 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22539 c_18_10_s1_s p_18_10_pi2j n8421 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22538 n8421 c_18_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22537 c_18_9_sum c_18_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22536 n8881 n8877 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22535 c_18_9_cout n8882 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22534 n8872 c_18_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22533 vdd p_18_9_pi2j n8872 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22532 n8882 c_18_9_cin n8872 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22531 n8882 c_18_9_a n8880 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22530 n8880 p_18_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22529 c_18_9_s2_s c_18_9_cin n8881 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22528 vdd c_18_9_s1_s n8877 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22527 c_18_9_s1_s c_18_9_a n8878 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22526 n8878 p_18_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22525 n8889 p_18_2_d2j n8891 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22524 n8891 p_18_2_d2jbar n8890 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22523 n8890 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22522 vdd a_8 n8889 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22521 vdd p_18_9_t_s n8885 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22520 n8885 p_18_1_n2j p_18_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22519 vdd n8891 n8886 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22518 n8886 n8888 p_18_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22517 n8888 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22516 vdd n9305 n9188 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22515 n9187 p_18_1_n2j p_18_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22514 vdd p_18_8_t_s n9187 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22513 vdd a_6 n9189 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22512 n9190 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22511 n9308 p_18_2_d2j n9190 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22510 n9189 p_18_2_d2jbar n9308 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22509 n9305 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22508 n9188 n9308 p_18_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22507 vdd c_18_8_a n9185 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22506 c_18_8_sum c_18_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22505 n9186 n9294 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22504 c_18_8_cout n9296 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22503 n9185 p_18_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22502 n9296 c_18_8_cin n9185 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22501 n9296 p_18_8_pi2j n8876 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22500 n8876 c_18_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22499 c_18_8_s2_s c_18_8_cin n9186 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22498 vdd c_18_8_s1_s n9294 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22497 c_18_8_s1_s p_18_8_pi2j n8875 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22496 n8875 c_18_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22495 c_18_7_sum c_18_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22494 n9649 n9646 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22493 c_18_7_cout n9651 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22492 n9640 c_18_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22491 vdd p_18_7_pi2j n9640 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22490 n9651 c_18_7_cin n9640 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22489 n9651 c_18_7_a n9648 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22488 n9648 p_18_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22487 c_18_7_s2_s c_18_7_cin n9649 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22486 vdd c_18_7_s1_s n9646 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22485 c_18_7_s1_s c_18_7_a n9647 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22484 n9647 p_18_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22483 n9536 p_18_2_d2j n9652 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22482 n9652 p_18_2_d2jbar n9538 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22481 n9538 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22480 vdd a_6 n9536 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22479 vdd p_18_7_t_s n9655 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22478 n9655 p_18_1_n2j p_18_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22477 vdd n9652 n9659 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22476 n9659 n9656 p_18_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22475 n9656 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22474 vdd n10091 n9657 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22473 n9653 p_18_1_n2j p_18_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22472 vdd p_18_6_t_s n9653 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22471 vdd a_4 n9660 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22470 n9661 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22469 n10090 p_18_2_d2j n9661 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22468 n9660 p_18_2_d2jbar n10090 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22467 n10091 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22466 n9657 n10090 p_18_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22465 vdd c_18_6_a n9985 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22464 c_18_6_sum c_18_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22463 n9986 n9987 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22462 c_18_6_cout n10084 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22461 n9985 p_18_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22460 n10084 c_18_6_cin n9985 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22459 n10084 p_18_6_pi2j n9644 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22458 n9644 c_18_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22457 c_18_6_s2_s c_18_6_cin n9986 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22456 vdd c_18_6_s1_s n9987 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22455 c_18_6_s1_s p_18_6_pi2j n9643 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22454 n9643 c_18_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22453 c_18_5_sum c_18_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22452 n10313 n10315 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22451 c_18_5_cout n10475 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22450 n10468 c_18_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22449 vdd c_18_5_b n10468 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22448 n10475 c_18_5_cin n10468 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22447 n10475 c_18_5_a n10476 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22446 n10476 c_18_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22445 c_18_5_s2_s c_18_5_cin n10313 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22444 vdd c_18_5_s1_s n10315 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22443 c_18_5_s1_s c_18_5_a n10474 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22442 n10474 c_18_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22441 n10319 p_18_2_d2j n10477 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22440 n10477 p_18_2_d2jbar n10320 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22439 n10320 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22438 vdd a_4 n10319 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22437 vdd p_18_5_t_s n10317 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22436 n10317 p_18_1_n2j c_18_5_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22435 vdd n10477 n10318 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22434 n10318 n10481 p_18_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22433 n10481 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22432 vdd n10742 n10482 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22431 n10479 p_18_1_n2j p_18_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22430 vdd p_18_4_t_s n10479 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22429 vdd a_2 n10483 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22428 n10484 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22427 n10744 p_18_2_d2j n10484 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22426 n10483 p_18_2_d2jbar n10744 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22425 n10742 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22424 n10482 n10744 p_18_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22423 vdd c_18_4_a n10469 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22422 c_18_4_sum c_18_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22421 n10737 n10738 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22420 c_18_4_cout n10735 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22419 n10469 p_18_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22418 n10735 c_18_4_cin n10469 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22417 n10735 p_18_4_pi2j n10472 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22416 n10472 c_18_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22415 c_18_4_s2_s c_18_4_cin n10737 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22414 vdd c_18_4_s1_s n10738 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22413 c_18_4_s1_s p_18_4_pi2j n10471 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22412 n10471 c_18_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22411 c_18_3_sum c_18_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22410 n11061 n11064 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22409 c_18_3_cout n11062 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22408 n11274 c_18_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22407 vdd c_18_3_b n11274 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22406 n11062 c_18_3_cin n11274 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22405 n11062 c_18_3_a n11280 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22404 n11280 c_18_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22403 c_18_3_s2_s c_18_3_cin n11061 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22402 vdd c_18_3_s1_s n11064 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22401 c_18_3_s1_s c_18_3_a n11279 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22400 n11279 c_18_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22399 n11070 p_18_2_d2j n11071 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22398 n11071 p_18_2_d2jbar n11072 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22397 n11072 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22396 vdd a_2 n11070 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22395 vdd p_18_3_t_s n11067 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22394 n11067 p_18_1_n2j c_18_3_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22393 vdd n11071 n11068 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22392 n11068 n11069 p_18_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22391 n11069 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22390 vdd n11495 n11284 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22389 n11282 p_18_1_n2j c_18_2_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22388 vdd p_18_2_t_s n11282 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22387 vdd a_0 n11285 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22386 n11286 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22385 n11496 p_18_2_d2j n11286 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22384 n11285 p_18_2_d2jbar n11496 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22383 n11495 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22382 n11284 n11496 p_18_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22381 vdd c_18_2_a n11275 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22380 c_18_2_sum c_18_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22379 n11277 n11489 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22378 c_18_2_cout n11487 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22377 n11275 c_18_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22376 n11487 c_18_2_cin n11275 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22375 n11487 c_18_2_b n11278 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22374 n11278 c_18_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22373 c_18_2_s2_s c_18_2_cin n11277 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22372 vdd c_18_2_s1_s n11489 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22371 c_18_2_s1_s c_18_2_b n11276 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22370 n11276 c_18_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22369 c_18_1_sum c_18_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22368 n11797 n11792 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22367 c_18_1_cout n11796 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22366 n11788 c_18_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22365 vdd p_18_1_pi2j n11788 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22364 n11796 c_18_1_cin n11788 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22363 n11796 c_18_1_a n11794 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22362 n11794 p_18_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22361 c_18_1_s2_s c_18_1_cin n11797 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22360 vdd c_18_1_s1_s n11792 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22359 c_18_1_s1_s c_18_1_a n11793 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22358 n11793 p_18_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22357 n11806 p_18_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22356 vdd a_0 n11806 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22355 vdd p_18_1_t_s n11801 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22354 n11801 p_18_1_n2j p_18_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22353 vdd n11806 n11803 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22352 n11803 n11805 p_18_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22351 n11805 p_18_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22350 n12089 c_17_1_sum cl4_18_s1_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22349 vdd n12187 n12089 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22348 p_28 cl4_18_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22347 n12176 c_17_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22346 vdd n12187 n12176 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22345 n12175 n12176 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22344 n12172 c_17_1_cout n12088 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22343 n12088 c_17_2_sum n12172 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22342 n12087 c_17_2_sum n12088 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_22341 vdd c_17_1_cout n12087 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_22340 n12088 c_17_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22339 vdd n12187 n12088 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22338 cla_cell0_0_a n12172 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22337 n12086 c_17_2_sum cl4_18_s2_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22336 vdd c_17_1_cout n12086 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22335 n12167 cl4_18_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_22334 n12085 n12175 cl4_18_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22333 vdd n12167 n12085 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22332 p_29 cl4_18_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22331 n68 p_17_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22330 c_17_33_s1_s c_17_31_a n68 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22329 vdd c_17_33_s1_s n65 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22328 c_17_33_s2_s c_17_32_cin n66 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22327 n63 p_17_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22326 n64 c_17_31_a n63 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22325 n64 c_17_32_cin n62 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22324 vdd p_17_33_pi2j n62 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22323 n62 c_17_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22322 c_18_32_cin n64 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22321 n66 n65 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22320 c_18_31_a c_17_33_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22319 n75 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22318 vdd p_17_33_t_s n71 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22317 n71 p_17_1_n2j p_17_33_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22316 vdd n75 n70 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22315 n70 n74 p_17_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22314 n74 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22313 vdd n422 n279 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22312 n278 p_17_1_n2j p_17_32_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22311 vdd p_17_32_t_s n278 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22310 vdd a_30 n280 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22309 n281 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22308 n424 p_17_2_d2j n281 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22307 n280 p_17_2_d2jbar n424 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22306 n422 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22305 n279 n424 p_17_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22304 n277 c_17_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22303 c_17_32_s1_s p_17_32_pi2j n277 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22302 vdd c_17_32_s1_s n418 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22301 c_17_32_s2_s c_17_32_cin n275 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22300 n276 c_17_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22299 n414 p_17_32_pi2j n276 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22298 n414 c_17_32_cin n274 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22297 vdd c_17_31_a n274 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22296 n274 p_17_32_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22295 c_18_31_cin n414 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22294 n275 n418 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22293 c_18_30_a c_17_32_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22292 c_18_29_a c_17_31_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22291 n723 n722 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22290 c_18_30_cin n726 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22289 n717 c_17_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22288 vdd p_17_31_pi2j n717 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22287 n726 c_17_31_cin n717 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22286 n726 c_17_31_a n724 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22285 n724 p_17_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22284 c_17_31_s2_s c_17_31_cin n723 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22283 vdd c_17_31_s1_s n722 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22282 c_17_31_s1_s c_17_31_a n720 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22281 n720 p_17_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22280 n733 p_17_2_d2j n731 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22279 n731 p_17_2_d2jbar n734 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22278 n734 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22277 vdd a_30 n733 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22276 vdd p_17_31_t_s n728 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22275 n728 p_17_1_n2j p_17_31_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22274 vdd n731 n727 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22273 n727 n732 p_17_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22272 n732 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22271 vdd n1163 n1001 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22270 n1000 p_17_1_n2j p_17_30_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22269 vdd p_17_30_t_s n1000 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22268 vdd a_28 n1002 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22267 n1003 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22266 n1165 p_17_2_d2j n1003 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22265 n1002 p_17_2_d2jbar n1165 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22264 n1163 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22263 n1001 n1165 p_17_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22262 n999 c_17_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22261 c_17_30_s1_s p_17_30_pi2j n999 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22260 vdd c_17_30_s1_s n1160 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22259 c_17_30_s2_s c_16_31_cout n998 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22258 n997 c_17_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22257 n1155 p_17_30_pi2j n997 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22256 n1155 c_16_31_cout n996 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22255 vdd c_17_30_a n996 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22254 n996 p_17_30_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22253 c_18_29_cin n1155 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22252 n998 n1160 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22251 c_18_28_a c_17_30_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22250 c_18_27_a c_17_29_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22249 n1485 n1484 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22248 c_18_28_cin n1488 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22247 n1477 c_17_29_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22246 vdd p_17_29_pi2j n1477 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22245 n1488 c_17_29_cin n1477 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22244 n1488 c_17_29_a n1486 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22243 n1486 p_17_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22242 c_17_29_s2_s c_17_29_cin n1485 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22241 vdd c_17_29_s1_s n1484 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22240 c_17_29_s1_s c_17_29_a n1482 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22239 n1482 p_17_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22238 n1494 p_17_2_d2j n1493 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22237 n1493 p_17_2_d2jbar n1496 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22236 n1496 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22235 vdd a_28 n1494 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22234 vdd p_17_29_t_s n1489 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22233 n1489 p_17_1_n2j p_17_29_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22232 vdd n1493 n1490 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22231 n1490 n1495 p_17_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22230 n1495 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22229 vdd n1925 n1782 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22228 n1783 p_17_1_n2j p_17_28_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22227 vdd p_17_28_t_s n1783 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22226 vdd a_26 n1784 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22225 n1785 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22224 n1927 p_17_2_d2j n1785 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22223 n1784 p_17_2_d2jbar n1927 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22222 n1925 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22221 n1782 n1927 p_17_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22220 n1481 c_17_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22219 c_17_28_s1_s p_17_28_pi2j n1481 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22218 vdd c_17_28_s1_s n1781 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22217 c_17_28_s2_s c_16_29_cout n1780 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22216 n1480 c_17_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22215 n1918 p_17_28_pi2j n1480 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22214 n1918 c_16_29_cout n1779 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22213 vdd c_17_28_a n1779 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22212 n1779 p_17_28_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22211 c_18_27_cin n1918 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22210 n1780 n1781 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22209 c_18_26_a c_17_28_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22208 c_18_25_a c_17_27_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22207 n2142 n2291 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22206 c_18_26_cin n2300 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22205 n2290 c_17_27_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22204 vdd c_17_27_b n2290 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22203 n2300 c_17_27_cin n2290 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22202 n2300 c_17_27_a n2297 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22201 n2297 c_17_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22200 c_17_27_s2_s c_17_27_cin n2142 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22199 vdd c_17_27_s1_s n2291 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22198 c_17_27_s1_s c_17_27_a n2299 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22197 n2299 c_17_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22196 n2144 p_17_2_d2j n2301 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22195 n2301 p_17_2_d2jbar n2146 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22194 n2146 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22193 vdd a_26 n2144 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22192 vdd p_17_27_t_s n2143 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22191 n2143 p_17_1_n2j c_17_27_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22190 vdd n2301 n2303 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22189 n2303 n2305 p_17_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22188 n2305 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22187 vdd n2600 n2304 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22186 n2302 p_17_1_n2j p_17_26_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22185 vdd p_17_26_t_s n2302 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22184 vdd a_24 n2307 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22183 n2308 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22182 n2601 p_17_2_d2j n2308 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22181 n2307 p_17_2_d2jbar n2601 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22180 n2600 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22179 n2304 n2601 p_17_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22178 n2296 c_17_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22177 c_17_26_s1_s p_17_26_pi2j n2296 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22176 vdd c_17_26_s1_s n2599 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22175 c_17_26_s2_s c_16_27_cout n2598 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22174 n2295 c_17_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22173 n2749 p_17_26_pi2j n2295 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22172 n2749 c_16_27_cout n2596 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22171 vdd c_17_26_a n2596 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22170 n2596 p_17_26_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22169 c_18_25_cin n2749 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22168 n2598 n2599 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22167 c_18_24_a c_17_26_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22166 c_18_23_a c_17_25_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22165 n2948 n2949 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22164 c_18_24_cin n3123 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22163 n3117 c_17_25_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22162 vdd c_17_25_b n3117 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22161 n3123 c_17_25_cin n3117 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22160 n3123 c_17_25_a n3124 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22159 n3124 c_17_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22158 c_17_25_s2_s c_17_25_cin n2948 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22157 vdd c_17_25_s1_s n2949 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22156 c_17_25_s1_s c_17_25_a n3125 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22155 n3125 c_17_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22154 n2953 p_17_2_d2j n2952 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22153 n2952 p_17_2_d2jbar n2954 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22152 n2954 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22151 vdd a_24 n2953 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22150 vdd p_17_25_t_s n2951 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22149 n2951 p_17_1_n2j c_17_25_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22148 vdd n2952 n2950 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22147 n2950 n3128 p_17_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22146 n3128 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22145 vdd n3371 n3127 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22144 n3126 p_17_1_n2j c_17_24_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22143 vdd p_17_24_t_s n3126 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22142 vdd a_22 n3130 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22141 n3131 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22140 n3372 p_17_2_d2j n3131 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22139 n3130 p_17_2_d2jbar n3372 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22138 n3371 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22137 n3127 n3372 p_17_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22136 n3121 c_17_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22135 c_17_24_s1_s c_17_24_b n3121 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22134 vdd c_17_24_s1_s n3368 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22133 c_17_24_s2_s c_16_25_cout n3366 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22132 n3120 c_17_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22131 n3364 c_17_24_b n3120 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22130 n3364 c_16_25_cout n3116 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22129 vdd c_17_24_a n3116 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22128 n3116 c_17_24_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22127 c_18_23_cin n3364 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22126 n3366 n3368 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22125 c_18_22_a c_17_24_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22124 c_18_21_a c_17_23_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22123 n3711 n3715 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22122 c_18_22_cin n3713 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22121 n3960 c_17_23_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22120 vdd c_17_23_b n3960 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22119 n3713 c_17_23_cin n3960 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22118 n3713 c_17_23_a n3710 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22117 n3710 c_17_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22116 c_17_23_s2_s c_17_23_cin n3711 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22115 vdd c_17_23_s1_s n3715 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22114 c_17_23_s1_s c_17_23_a n3709 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22113 n3709 c_17_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22112 n3721 p_17_2_d2j n3719 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22111 n3719 p_17_2_d2jbar n3722 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22110 n3722 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22109 vdd a_22 n3721 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22108 vdd p_17_23_t_s n3717 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22107 n3717 p_17_1_n2j c_17_23_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22106 vdd n3719 n3716 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22105 n3716 n3720 p_17_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22104 n3720 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22103 vdd n4151 n3966 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22102 n3965 p_17_1_n2j p_17_22_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22101 vdd p_17_22_t_s n3965 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22100 vdd a_20 n3967 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22099 n3968 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22098 n4153 p_17_2_d2j n3968 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22097 n3967 p_17_2_d2jbar n4153 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22096 n4151 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22095 n3966 n4153 p_17_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22094 n3964 c_17_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22093 c_17_22_s1_s p_17_22_pi2j n3964 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22092 vdd c_17_22_s1_s n4147 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22091 c_17_22_s2_s c_16_23_cout n3962 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22090 n3963 c_17_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22089 n4143 p_17_22_pi2j n3963 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22088 n4143 c_16_23_cout n3959 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22087 vdd c_17_22_a n3959 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22086 n3959 p_17_22_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22085 c_18_21_cin n4143 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22084 n3962 n4147 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22083 c_18_20_a c_17_22_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22082 c_18_19_a c_17_21_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22081 n4470 n4469 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22080 c_18_20_cin n4472 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22079 n4464 c_17_21_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22078 vdd p_17_21_pi2j n4464 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22077 n4472 c_17_21_cin n4464 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22076 n4472 c_17_21_a n4471 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22075 n4471 p_17_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22074 c_17_21_s2_s c_17_21_cin n4470 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22073 vdd c_17_21_s1_s n4469 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22072 c_17_21_s1_s c_17_21_a n4467 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22071 n4467 p_17_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22070 n4480 p_17_2_d2j n4478 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22069 n4478 p_17_2_d2jbar n4481 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22068 n4481 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22067 vdd a_20 n4480 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22066 vdd p_17_21_t_s n4475 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22065 n4475 p_17_1_n2j p_17_21_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22064 vdd n4478 n4474 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22063 n4474 n4479 p_17_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22062 n4479 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22061 vdd n4897 n4744 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22060 n4743 p_17_1_n2j p_17_20_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22059 vdd p_17_20_t_s n4743 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22058 vdd a_18 n4745 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22057 n4746 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22056 n4899 p_17_2_d2j n4746 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22055 n4745 p_17_2_d2jbar n4899 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22054 n4897 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22053 n4744 n4899 p_17_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22052 n4742 c_17_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22051 c_17_20_s1_s p_17_20_pi2j n4742 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22050 vdd c_17_20_s1_s n4895 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22049 c_17_20_s2_s c_16_21_cout n4741 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22048 n4740 c_17_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22047 n4890 p_17_20_pi2j n4740 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22046 n4890 c_16_21_cout n4739 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22045 vdd c_17_20_a n4739 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22044 n4739 p_17_20_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22043 c_18_19_cin n4890 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22042 n4741 n4895 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22041 c_18_18_a c_17_20_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22040 c_18_17_a c_17_19_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22039 n5213 n5209 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_22038 c_18_18_cin n5214 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22037 n5204 c_17_19_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22036 vdd p_17_19_pi2j n5204 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22035 n5214 c_17_19_cin n5204 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22034 n5214 c_17_19_a n5212 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22033 n5212 p_17_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22032 c_17_19_s2_s c_17_19_cin n5213 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22031 vdd c_17_19_s1_s n5209 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22030 c_17_19_s1_s c_17_19_a n5210 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22029 n5210 p_17_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22028 n5221 p_17_2_d2j n5220 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22027 n5220 p_17_2_d2jbar n5223 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22026 n5223 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22025 vdd a_18 n5221 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22024 vdd p_17_19_t_s n5216 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22023 n5216 p_17_1_n2j p_17_19_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22022 vdd n5220 n5217 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22021 n5217 n5222 p_17_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22020 n5222 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22019 vdd n5653 n5509 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22018 n5508 p_17_1_n2j p_17_18_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22017 vdd p_17_18_t_s n5508 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22016 vdd a_16 n5510 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22015 n5511 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_22014 n5651 p_17_2_d2j n5511 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22013 n5510 p_17_2_d2jbar n5651 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_22012 n5653 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22011 n5509 n5651 p_17_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_22010 n5207 c_17_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22009 c_17_18_s1_s p_17_18_pi2j n5207 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22008 vdd c_17_18_s1_s n5507 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_22007 c_17_18_s2_s c_16_19_cout n5506 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_22006 n5208 c_17_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22005 n5642 p_17_18_pi2j n5208 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22004 n5642 c_16_19_cout n5505 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22003 vdd c_17_18_a n5505 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22002 n5505 p_17_18_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_22001 c_18_17_cin n5642 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_22000 n5506 n5507 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21999 c_18_16_a c_17_18_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21998 c_18_15_a c_17_17_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21997 n5986 n5979 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21996 c_18_16_cin n5989 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21995 n5978 c_17_17_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21994 vdd p_17_17_pi2j n5978 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21993 n5989 c_17_17_cin n5978 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21992 n5989 c_17_17_a n5987 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21991 n5987 p_17_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21990 c_17_17_s2_s c_17_17_cin n5986 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21989 vdd c_17_17_s1_s n5979 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21988 c_17_17_s1_s c_17_17_a n5985 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21987 n5985 p_17_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21986 n5863 p_17_2_d2j n5990 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21985 n5990 p_17_2_d2jbar n5865 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21984 n5865 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21983 vdd a_16 n5863 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21982 vdd p_17_17_t_s n5994 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21981 n5994 p_17_1_n2j p_17_17_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21980 vdd n5990 n5992 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21979 n5992 n5996 p_17_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21978 n5996 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21977 vdd n6442 n5993 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21976 n5991 p_17_1_n2j p_17_16_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21975 vdd p_17_16_t_s n5991 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21974 vdd a_14 n5998 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21973 n5999 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21972 n6310 p_17_2_d2j n5999 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21971 n5998 p_17_2_d2jbar n6310 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21970 n6442 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21969 n5993 n6310 p_17_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21968 n5983 c_17_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21967 c_17_16_s1_s p_17_16_pi2j n5983 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21966 vdd c_17_16_s1_s n6309 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21965 c_17_16_s2_s c_16_17_cout n6308 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21964 n5982 c_17_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21963 n6436 p_17_16_pi2j n5982 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21962 n6436 c_16_17_cout n6306 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21961 vdd c_17_16_a n6306 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21960 n6306 p_17_16_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21959 c_18_15_cin n6436 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21958 n6308 n6309 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21957 c_18_14_a c_17_16_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21956 c_18_13_a c_17_15_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21955 n6649 n6650 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21954 c_18_14_cin n6826 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21953 n6819 c_17_15_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21952 vdd c_17_15_b n6819 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21951 n6826 c_17_15_cin n6819 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21950 n6826 c_17_15_a n6827 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21949 n6827 c_17_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21948 c_17_15_s2_s c_17_15_cin n6649 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21947 vdd c_17_15_s1_s n6650 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21946 c_17_15_s1_s c_17_15_a n6824 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21945 n6824 c_17_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21944 n6654 p_17_2_d2j n6653 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21943 n6653 p_17_2_d2jbar n6655 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21942 n6655 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21941 vdd a_14 n6654 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21940 vdd p_17_15_t_s n6652 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21939 n6652 p_17_1_n2j c_17_15_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21938 vdd n6653 n6651 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21937 n6651 n6830 p_17_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21936 n6830 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21935 vdd n7077 n6829 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21934 n6828 p_17_1_n2j p_17_14_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21933 vdd p_17_14_t_s n6828 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21932 vdd a_12 n6832 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21931 n6833 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21930 n7078 p_17_2_d2j n6833 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21929 n6832 p_17_2_d2jbar n7078 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21928 n7077 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21927 n6829 n7078 p_17_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21926 n6823 c_17_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21925 c_17_14_s1_s p_17_14_pi2j n6823 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21924 vdd c_17_14_s1_s n7074 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21923 c_17_14_s2_s c_16_15_cout n7072 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21922 n6822 c_17_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21921 n7071 p_17_14_pi2j n6822 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21920 n7071 c_16_15_cout n6818 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21919 vdd c_17_14_a n6818 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21918 n6818 p_17_14_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21917 c_18_13_cin n7071 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21916 n7072 n7074 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21915 c_18_12_a c_17_14_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21914 c_18_11_a c_17_13_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21913 n7410 n7414 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21912 c_18_12_cin n7411 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21911 n7623 c_17_13_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21910 vdd c_17_13_b n7623 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21909 n7411 c_17_13_cin n7623 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21908 n7411 c_17_13_a n7629 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21907 n7629 c_17_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21906 c_17_13_s2_s c_17_13_cin n7410 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21905 vdd c_17_13_s1_s n7414 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21904 c_17_13_s1_s c_17_13_a n7628 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21903 n7628 c_17_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21902 n7419 p_17_2_d2j n7417 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21901 n7417 p_17_2_d2jbar n7420 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21900 n7420 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21899 vdd a_12 n7419 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21898 vdd p_17_13_t_s n7416 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21897 n7416 p_17_1_n2j c_17_13_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21896 vdd n7417 n7415 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21895 n7415 n7418 p_17_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21894 n7418 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21893 vdd n7843 n7631 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21892 n7630 p_17_1_n2j c_17_12_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21891 vdd p_17_12_t_s n7630 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21890 vdd a_10 n7633 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21889 n7634 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21888 n7845 p_17_2_d2j n7634 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21887 n7633 p_17_2_d2jbar n7845 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21886 n7843 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21885 n7631 n7845 p_17_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21884 n7627 c_17_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21883 c_17_12_s1_s c_17_12_b n7627 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21882 vdd c_17_12_s1_s n7840 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21881 c_17_12_s2_s c_16_13_cout n7625 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21880 n7626 c_17_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21879 n7837 c_17_12_b n7626 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21878 n7837 c_16_13_cout n7622 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21877 vdd c_17_12_a n7622 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21876 n7622 c_17_12_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21875 c_18_11_cin n7837 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21874 n7625 n7840 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21873 c_18_10_a c_17_12_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21872 c_18_9_a c_17_11_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21871 n8161 n8155 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21870 c_18_10_cin n8159 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21869 n8152 c_17_11_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21868 vdd p_17_11_pi2j n8152 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21867 n8159 c_17_11_cin n8152 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21866 n8159 c_17_11_a n8157 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21865 n8157 p_17_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21864 c_17_11_s2_s c_17_11_cin n8161 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21863 vdd c_17_11_s1_s n8155 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21862 c_17_11_s1_s c_17_11_a n8156 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21861 n8156 p_17_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21860 n8168 p_17_2_d2j n8166 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21859 n8166 p_17_2_d2jbar n8169 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21858 n8169 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21857 vdd a_10 n8168 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21856 vdd p_17_11_t_s n8163 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21855 n8163 p_17_1_n2j p_17_11_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21854 vdd n8166 n8162 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21853 n8162 n8167 p_17_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21852 n8167 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21851 vdd n8586 n8433 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21850 n8432 p_17_1_n2j p_17_10_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21849 vdd p_17_10_t_s n8432 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21848 vdd a_8 n8434 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21847 n8435 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21846 n8588 p_17_2_d2j n8435 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21845 n8434 p_17_2_d2jbar n8588 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21844 n8586 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21843 n8433 n8588 p_17_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21842 n8431 c_17_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21841 c_17_10_s1_s p_17_10_pi2j n8431 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21840 vdd c_17_10_s1_s n8584 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21839 c_17_10_s2_s c_16_11_cout n8430 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21838 n8429 c_17_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21837 n8579 p_17_10_pi2j n8429 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21836 n8579 c_16_11_cout n8428 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21835 vdd c_17_10_a n8428 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21834 n8428 p_17_10_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21833 c_18_9_cin n8579 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21832 n8430 n8584 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21831 c_18_8_a c_17_10_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21830 c_18_7_a c_17_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21829 n8901 n8897 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21828 c_18_8_cin n8902 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21827 n8892 c_17_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21826 vdd p_17_9_pi2j n8892 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21825 n8902 c_17_9_cin n8892 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21824 n8902 c_17_9_a n8900 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21823 n8900 p_17_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21822 c_17_9_s2_s c_17_9_cin n8901 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21821 vdd c_17_9_s1_s n8897 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21820 c_17_9_s1_s c_17_9_a n8898 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21819 n8898 p_17_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21818 n8909 p_17_2_d2j n8908 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21817 n8908 p_17_2_d2jbar n8911 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21816 n8911 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21815 vdd a_8 n8909 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21814 vdd p_17_9_t_s n8904 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21813 n8904 p_17_1_n2j p_17_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21812 vdd n8908 n8905 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21811 n8905 n8910 p_17_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21810 n8910 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21809 vdd n9322 n9194 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21808 n9193 p_17_1_n2j p_17_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21807 vdd p_17_8_t_s n9193 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21806 vdd a_6 n9195 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21805 n9196 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21804 n9320 p_17_2_d2j n9196 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21803 n9195 p_17_2_d2jbar n9320 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21802 n9322 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21801 n9194 n9320 p_17_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21800 n8895 c_17_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21799 c_17_8_s1_s p_17_8_pi2j n8895 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21798 vdd c_17_8_s1_s n9309 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21797 c_17_8_s2_s c_16_9_cout n9192 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21796 n8896 c_17_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21795 n9311 p_17_8_pi2j n8896 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21794 n9311 c_16_9_cout n9191 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21793 vdd c_17_8_a n9191 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21792 n9191 p_17_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21791 c_18_7_cin n9311 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21790 n9192 n9309 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21789 c_18_6_a c_17_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21788 c_18_5_a c_17_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21787 n9672 n9667 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21786 c_18_6_cin n9670 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21785 n9662 c_17_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21784 vdd p_17_7_pi2j n9662 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21783 n9670 c_17_7_cin n9662 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21782 n9670 c_17_7_a n9673 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21781 n9673 p_17_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21780 c_17_7_s2_s c_17_7_cin n9672 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21779 vdd c_17_7_s1_s n9667 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21778 c_17_7_s1_s c_17_7_a n9668 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21777 n9668 p_17_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21776 n9541 p_17_2_d2j n9674 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21775 n9674 p_17_2_d2jbar n9543 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21774 n9543 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21773 vdd a_6 n9541 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21772 vdd p_17_7_t_s n9677 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21771 n9677 p_17_1_n2j p_17_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21770 vdd n9674 n9678 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21769 n9678 n9680 p_17_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21768 n9680 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21767 vdd n10104 n9675 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21766 n9676 p_17_1_n2j p_17_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21765 vdd p_17_6_t_s n9676 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21764 vdd a_4 n9682 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21763 n9683 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21762 n10105 p_17_2_d2j n9683 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21761 n9682 p_17_2_d2jbar n10105 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21760 n10104 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21759 n9675 n10105 p_17_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21758 n9666 c_17_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21757 c_17_6_s1_s p_17_6_pi2j n9666 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21756 vdd c_17_6_s1_s n9992 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21755 c_17_6_s2_s c_16_7_cout n9991 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21754 n9665 c_17_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21753 n10097 p_17_6_pi2j n9665 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21752 n10097 c_16_7_cout n9990 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21751 vdd c_17_6_a n9990 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21750 n9990 p_17_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21749 c_18_5_cin n10097 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21748 n9991 n9992 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21747 c_18_4_a c_17_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21746 c_18_3_a c_17_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21745 n10323 n10325 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21744 c_18_4_cin n10494 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21743 n10486 c_17_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21742 vdd c_17_5_b n10486 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21741 n10494 c_17_5_cin n10486 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21740 n10494 c_17_5_a n10491 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21739 n10491 c_17_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21738 c_17_5_s2_s c_17_5_cin n10323 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21737 vdd c_17_5_s1_s n10325 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21736 c_17_5_s1_s c_17_5_a n10493 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21735 n10493 c_17_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21734 n10328 p_17_2_d2j n10495 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21733 n10495 p_17_2_d2jbar n10329 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21732 n10329 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21731 vdd a_4 n10328 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21730 vdd p_17_5_t_s n10327 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21729 n10327 p_17_1_n2j c_17_5_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21728 vdd n10495 n10326 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21727 n10326 n10498 p_17_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21726 n10498 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21725 vdd n10751 n10497 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21724 n10496 p_17_1_n2j p_17_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21723 vdd p_17_4_t_s n10496 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21722 vdd a_2 n10500 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21721 n10501 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21720 n10752 p_17_2_d2j n10501 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21719 n10500 p_17_2_d2jbar n10752 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21718 n10751 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21717 n10497 n10752 p_17_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21716 n10490 c_17_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21715 c_17_4_s1_s p_17_4_pi2j n10490 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21714 vdd c_17_4_s1_s n10750 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21713 c_17_4_s2_s c_16_5_cout n10747 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21712 n10489 c_17_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21711 n10745 p_17_4_pi2j n10489 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21710 n10745 c_16_5_cout n10485 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21709 vdd c_17_4_a n10485 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21708 n10485 p_17_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21707 c_18_3_cin n10745 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21706 n10747 n10750 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21705 c_18_2_a c_17_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21704 c_18_1_a c_17_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21703 n11075 n11079 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21702 c_18_2_cin n11076 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21701 n11288 c_17_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21700 vdd c_17_3_b n11288 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21699 n11076 c_17_3_cin n11288 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21698 n11076 c_17_3_a n11294 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21697 n11294 c_17_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21696 c_17_3_s2_s c_17_3_cin n11075 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21695 vdd c_17_3_s1_s n11079 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21694 c_17_3_s1_s c_17_3_a n11293 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21693 n11293 c_17_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21692 n11084 p_17_2_d2j n11082 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21691 n11082 p_17_2_d2jbar n11085 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21690 n11085 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21689 vdd a_2 n11084 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21688 vdd p_17_3_t_s n11081 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21687 n11081 p_17_1_n2j c_17_3_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21686 vdd n11082 n11080 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21685 n11080 n11083 p_17_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21684 n11083 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21683 vdd n11506 n11296 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21682 n11295 p_17_1_n2j c_17_2_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21681 vdd p_17_2_t_s n11295 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21680 vdd a_0 n11298 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21679 n11299 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21678 n11508 p_17_2_d2j n11299 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21677 n11298 p_17_2_d2jbar n11508 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21676 n11506 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21675 n11296 n11508 p_17_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21674 n11292 c_17_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21673 c_17_2_s1_s c_17_2_b n11292 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21672 vdd c_17_2_s1_s n11503 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21671 c_17_2_s2_s c_16_3_cout n11290 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21670 n11291 c_17_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21669 n11500 c_17_2_b n11291 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21668 n11500 c_16_3_cout n11287 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21667 vdd c_17_2_a n11287 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21666 n11287 c_17_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21665 c_18_1_cin n11500 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21664 n11290 n11503 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21663 c_17_2_sum c_17_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21662 c_17_1_sum c_17_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21661 n11814 n11813 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21660 c_17_1_cout n11816 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21659 n11808 c_17_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21658 vdd p_17_1_pi2j n11808 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21657 n11816 c_17_1_cin n11808 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21656 n11816 c_17_1_a n11815 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21655 n11815 p_17_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21654 c_17_1_s2_s c_17_1_cin n11814 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21653 vdd c_17_1_s1_s n11813 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21652 c_17_1_s1_s c_17_1_a n11811 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21651 n11811 p_17_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21650 n11825 p_17_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21649 vdd a_0 n11825 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21648 vdd p_17_1_t_s n11820 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21647 n11820 p_17_1_n2j p_17_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21646 vdd n11825 n11819 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21645 n11819 n11824 p_17_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21644 n11824 p_17_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21643 n12094 c_16_1_sum cl4_17_s1_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21642 vdd n12204 n12094 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21641 p_26 cl4_17_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21640 n12193 c_16_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21639 vdd n12204 n12193 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21638 n12192 n12193 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21637 n12191 c_16_1_cout n12093 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21636 n12093 c_16_2_sum n12191 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21635 n12092 c_16_2_sum n12093 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_21634 vdd c_16_1_cout n12092 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_21633 n12093 c_16_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21632 vdd n12204 n12093 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21631 n12187 n12191 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21630 n12091 c_16_2_sum cl4_17_s2_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21629 vdd c_16_1_cout n12091 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21628 n12185 cl4_17_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_21627 n12090 n12192 cl4_17_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21626 vdd n12185 n12090 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21625 p_27 cl4_17_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21624 n83 p_16_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21623 c_16_33_s1_s c_16_31_a n83 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21622 vdd c_16_33_s1_s n81 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21621 c_16_33_s2_s c_16_32_cin n82 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21620 n79 p_16_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21619 n80 c_16_31_a n79 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21618 n80 c_16_32_cin n77 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21617 vdd p_16_33_pi2j n77 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21616 n77 c_16_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21615 c_17_32_cin n80 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21614 n82 n81 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21613 c_17_31_a c_16_33_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21612 n89 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21611 vdd p_16_33_t_s n78 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21610 n78 p_16_1_n2j p_16_33_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21609 vdd n89 n87 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21608 n87 n88 p_16_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21607 n88 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21606 vdd n435 n287 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21605 n286 p_16_1_n2j p_16_32_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21604 vdd p_16_32_t_s n286 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21603 vdd a_30 n289 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21602 n288 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21601 n437 p_16_2_d2j n288 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21600 n289 p_16_2_d2jbar n437 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21599 n435 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21598 n287 n437 p_16_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21597 n285 c_16_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21596 c_16_32_s1_s p_16_32_pi2j n285 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21595 vdd c_16_32_s1_s n431 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21594 c_16_32_s2_s c_16_32_cin n284 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21593 n283 c_16_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21592 n425 p_16_32_pi2j n283 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21591 n425 c_16_32_cin n282 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21590 vdd c_16_31_a n282 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21589 n282 p_16_32_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21588 c_17_31_cin n425 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21587 n284 n431 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21586 c_17_30_a c_16_32_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21585 c_17_29_a c_16_31_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21584 n744 n740 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21583 c_16_31_cout n745 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21582 n737 c_16_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21581 vdd p_16_31_pi2j n737 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21580 n745 c_16_31_cin n737 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21579 n745 c_16_31_a n743 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21578 n743 p_16_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21577 c_16_31_s2_s c_16_31_cin n744 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21576 vdd c_16_31_s1_s n740 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21575 c_16_31_s1_s c_16_31_a n741 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21574 n741 p_16_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21573 n752 p_16_2_d2j n751 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21572 n751 p_16_2_d2jbar n750 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21571 n750 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21570 vdd a_30 n752 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21569 vdd p_16_31_t_s n739 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21568 n739 p_16_1_n2j p_16_31_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21567 vdd n751 n748 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21566 n748 n749 p_16_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21565 n749 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21564 vdd n1178 n1009 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21563 n1008 p_16_1_n2j p_16_30_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21562 vdd p_16_30_t_s n1008 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21561 vdd a_28 n1011 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21560 n1010 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21559 n1181 p_16_2_d2j n1010 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21558 n1011 p_16_2_d2jbar n1181 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21557 n1178 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21556 n1009 n1181 p_16_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21555 n1007 c_16_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21554 c_16_30_s1_s p_16_30_pi2j n1007 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21553 vdd c_16_30_s1_s n1173 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21552 c_16_30_s2_s c_15_31_cout n1005 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21551 n1006 c_16_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21550 n1167 p_16_30_pi2j n1006 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21549 n1167 c_15_31_cout n1004 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21548 vdd c_16_30_a n1004 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21547 n1004 p_16_30_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21546 c_17_29_cin n1167 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21545 n1005 n1173 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21544 c_17_28_a c_16_30_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21543 c_17_27_a c_16_29_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21542 n1507 n1506 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21541 c_16_29_cout n1509 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21540 n1499 c_16_29_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21539 vdd p_16_29_pi2j n1499 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21538 n1509 c_16_29_cin n1499 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21537 n1509 c_16_29_a n1508 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21536 n1508 p_16_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21535 c_16_29_s2_s c_16_29_cin n1507 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21534 vdd c_16_29_s1_s n1506 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21533 c_16_29_s1_s c_16_29_a n1503 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21532 n1503 p_16_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21531 n1514 p_16_2_d2j n1516 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21530 n1516 p_16_2_d2jbar n1515 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21529 n1515 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21528 vdd a_28 n1514 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21527 vdd p_16_29_t_s n1504 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21526 n1504 p_16_1_n2j p_16_29_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21525 vdd n1516 n1512 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21524 n1512 n1513 p_16_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21523 n1513 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21522 vdd n1939 n1790 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21521 n1788 p_16_1_n2j p_16_28_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21520 vdd p_16_28_t_s n1788 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21519 vdd a_26 n1791 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21518 n1792 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21517 n1942 p_16_2_d2j n1792 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21516 n1791 p_16_2_d2jbar n1942 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21515 n1939 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21514 n1790 n1942 p_16_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21513 n1502 c_16_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21512 c_16_28_s1_s p_16_28_pi2j n1502 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21511 vdd c_16_28_s1_s n1789 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21510 c_16_28_s2_s c_15_29_cout n1787 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21509 n1501 c_16_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21508 n1929 p_16_28_pi2j n1501 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21507 n1929 c_15_29_cout n1786 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21506 vdd c_16_28_a n1786 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21505 n1786 p_16_28_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21504 c_17_27_cin n1929 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21503 n1787 n1789 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21502 c_17_26_a c_16_28_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21501 c_17_25_a c_16_27_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21500 n2150 n2312 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21499 c_16_27_cout n2320 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21498 n2311 c_16_27_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21497 vdd c_16_27_b n2311 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21496 n2320 c_16_27_cin n2311 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21495 n2320 c_16_27_a n2321 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21494 n2321 c_16_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21493 c_16_27_s2_s c_16_27_cin n2150 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21492 vdd c_16_27_s1_s n2312 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21491 c_16_27_s1_s c_16_27_a n2318 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21490 n2318 c_16_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21489 n2152 p_16_2_d2j n2322 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21488 n2322 p_16_2_d2jbar n2151 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21487 n2151 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21486 vdd a_26 n2152 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21485 vdd p_16_27_t_s n2149 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21484 n2149 p_16_1_n2j c_16_27_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21483 vdd n2322 n2325 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21482 n2325 n2323 p_16_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21481 n2323 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21480 vdd n2608 n2326 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21479 n2319 p_16_1_n2j p_16_26_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21478 vdd p_16_26_t_s n2319 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21477 vdd a_24 n2328 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21476 n2327 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21475 n2610 p_16_2_d2j n2327 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21474 n2328 p_16_2_d2jbar n2610 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21473 n2608 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21472 n2326 n2610 p_16_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21471 n2316 c_16_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21470 c_16_26_s1_s p_16_26_pi2j n2316 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21469 vdd c_16_26_s1_s n2607 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21468 c_16_26_s2_s c_15_27_cout n2606 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21467 n2315 c_16_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21466 n2758 p_16_26_pi2j n2315 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21465 n2758 c_15_27_cout n2604 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21464 vdd c_16_26_a n2604 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21463 n2604 p_16_26_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21462 c_17_25_cin n2758 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21461 n2606 n2607 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21460 c_17_24_a c_16_26_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21459 c_17_23_a c_16_25_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21458 n2958 n2959 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21457 c_16_25_cout n3141 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21456 n3133 c_16_25_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21455 vdd c_16_25_b n3133 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21454 n3141 c_16_25_cin n3133 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21453 n3141 c_16_25_a n3142 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21452 n3142 c_16_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21451 c_16_25_s2_s c_16_25_cin n2958 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21450 vdd c_16_25_s1_s n2959 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21449 c_16_25_s1_s c_16_25_a n3139 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21448 n3139 c_16_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21447 n2963 p_16_2_d2j n2962 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21446 n2962 p_16_2_d2jbar n2961 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21445 n2961 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21444 vdd a_24 n2963 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21443 vdd p_16_25_t_s n2957 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21442 n2957 p_16_1_n2j c_16_25_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21441 vdd n2962 n2960 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21440 n2960 n3143 p_16_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21439 n3143 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21438 vdd n3382 n3145 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21437 n3140 p_16_1_n2j c_16_24_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21436 vdd p_16_24_t_s n3140 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21435 vdd a_22 n3147 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21434 n3146 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21433 n3384 p_16_2_d2j n3146 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21432 n3147 p_16_2_d2jbar n3384 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21431 n3382 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21430 n3145 n3384 p_16_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21429 n3137 c_16_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21428 c_16_24_s1_s c_16_24_b n3137 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21427 vdd c_16_24_s1_s n3379 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21426 c_16_24_s2_s c_15_25_cout n3378 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21425 n3136 c_16_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21424 n3375 c_16_24_b n3136 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21423 n3375 c_15_25_cout n3132 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21422 vdd c_16_24_a n3132 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21421 n3132 c_16_24_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21420 c_17_23_cin n3375 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21419 n3378 n3379 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21418 c_17_22_a c_16_24_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21417 c_17_21_a c_16_23_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21416 n3729 n3732 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21415 c_16_23_cout n3731 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21414 n3970 c_16_23_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21413 vdd c_16_23_b n3970 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21412 n3731 c_16_23_cin n3970 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21411 n3731 c_16_23_a n3730 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21410 n3730 c_16_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21409 c_16_23_s2_s c_16_23_cin n3729 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21408 vdd c_16_23_s1_s n3732 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21407 c_16_23_s1_s c_16_23_a n3726 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21406 n3726 c_16_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21405 n3738 p_16_2_d2j n3737 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21404 n3737 p_16_2_d2jbar n3736 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21403 n3736 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21402 vdd a_22 n3738 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21401 vdd p_16_23_t_s n3727 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21400 n3727 p_16_1_n2j c_16_23_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21399 vdd n3737 n3734 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21398 n3734 n3735 p_16_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21397 n3735 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21396 vdd n4166 n3976 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21395 n3975 p_16_1_n2j p_16_22_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21394 vdd p_16_22_t_s n3975 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21393 vdd a_20 n3978 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21392 n3977 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21391 n4168 p_16_2_d2j n3977 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21390 n3978 p_16_2_d2jbar n4168 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21389 n4166 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21388 n3976 n4168 p_16_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21387 n3974 c_16_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21386 c_16_22_s1_s p_16_22_pi2j n3974 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21385 vdd c_16_22_s1_s n4161 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21384 c_16_22_s2_s c_15_23_cout n3973 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21383 n3972 c_16_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21382 n4155 p_16_22_pi2j n3972 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21381 n4155 c_15_23_cout n3969 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21380 vdd c_16_22_a n3969 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21379 n3969 p_16_22_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21378 c_17_21_cin n4155 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21377 n3973 n4161 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21376 c_17_20_a c_16_22_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21375 c_17_19_a c_16_21_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21374 n4490 n4489 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21373 c_16_21_cout n4492 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21372 n4484 c_16_21_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21371 vdd p_16_21_pi2j n4484 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21370 n4492 c_16_21_cin n4484 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21369 n4492 c_16_21_a n4491 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21368 n4491 p_16_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21367 c_16_21_s2_s c_16_21_cin n4490 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21366 vdd c_16_21_s1_s n4489 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21365 c_16_21_s1_s c_16_21_a n4486 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21364 n4486 p_16_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21363 n4499 p_16_2_d2j n4498 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21362 n4498 p_16_2_d2jbar n4497 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21361 n4497 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21360 vdd a_20 n4499 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21359 vdd p_16_21_t_s n4487 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21358 n4487 p_16_1_n2j p_16_21_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21357 vdd n4498 n4495 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21356 n4495 n4496 p_16_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21355 n4496 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21354 vdd n4912 n4752 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21353 n4751 p_16_1_n2j p_16_20_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21352 vdd p_16_20_t_s n4751 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21351 vdd a_18 n4754 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21350 n4753 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21349 n4914 p_16_2_d2j n4753 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21348 n4754 p_16_2_d2jbar n4914 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21347 n4912 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21346 n4752 n4914 p_16_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21345 n4750 c_16_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21344 c_16_20_s1_s p_16_20_pi2j n4750 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21343 vdd c_16_20_s1_s n4909 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21342 c_16_20_s2_s c_15_21_cout n4748 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21341 n4749 c_16_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21340 n4901 p_16_20_pi2j n4749 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21339 n4901 c_15_21_cout n4747 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21338 vdd c_16_20_a n4747 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21337 n4747 p_16_20_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21336 c_17_19_cin n4901 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21335 n4748 n4909 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21334 c_17_18_a c_16_20_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21333 c_17_17_a c_16_19_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21332 n5234 n5232 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21331 c_16_19_cout n5236 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21330 n5226 c_16_19_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21329 vdd p_16_19_pi2j n5226 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21328 n5236 c_16_19_cin n5226 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21327 n5236 c_16_19_a n5235 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21326 n5235 p_16_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21325 c_16_19_s2_s c_16_19_cin n5234 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21324 vdd c_16_19_s1_s n5232 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21323 c_16_19_s1_s c_16_19_a n5233 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21322 n5233 p_16_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21321 n5241 p_16_2_d2j n5243 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21320 n5243 p_16_2_d2jbar n5242 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21319 n5242 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21318 vdd a_18 n5241 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21317 vdd p_16_19_t_s n5230 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21316 n5230 p_16_1_n2j p_16_19_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21315 vdd n5243 n5239 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21314 n5239 n5240 p_16_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21313 n5240 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21312 vdd n5667 n5516 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21311 n5514 p_16_1_n2j p_16_18_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21310 vdd p_16_18_t_s n5514 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21309 vdd a_16 n5518 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21308 n5517 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21307 n5666 p_16_2_d2j n5517 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21306 n5518 p_16_2_d2jbar n5666 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21305 n5667 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21304 n5516 n5666 p_16_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21303 n5229 c_16_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21302 c_16_18_s1_s p_16_18_pi2j n5229 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21301 vdd c_16_18_s1_s n5515 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21300 c_16_18_s2_s c_15_19_cout n5513 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21299 n5228 c_16_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21298 n5656 p_16_18_pi2j n5228 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21297 n5656 c_15_19_cout n5512 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21296 vdd c_16_18_a n5512 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21295 n5512 p_16_18_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21294 c_17_17_cin n5656 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21293 n5513 n5515 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21292 c_17_16_a c_16_18_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21291 c_17_15_a c_16_17_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21290 n6012 n6003 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21289 c_16_17_cout n6013 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21288 n6002 c_16_17_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21287 vdd p_16_17_pi2j n6002 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21286 n6013 c_16_17_cin n6002 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21285 n6013 c_16_17_a n6011 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21284 n6011 p_16_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21283 c_16_17_s2_s c_16_17_cin n6012 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21282 vdd c_16_17_s1_s n6003 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21281 c_16_17_s1_s c_16_17_a n6010 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21280 n6010 p_16_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21279 n5869 p_16_2_d2j n6014 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21278 n6014 p_16_2_d2jbar n5868 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21277 n5868 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21276 vdd a_16 n5869 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21275 vdd p_16_17_t_s n6007 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21274 n6007 p_16_1_n2j p_16_17_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21273 vdd n6014 n6016 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21272 n6016 n6015 p_16_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21271 n6015 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21270 vdd n6454 n6017 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21269 n6008 p_16_1_n2j p_16_16_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21268 vdd p_16_16_t_s n6008 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21267 vdd a_14 n6021 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21266 n6020 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21265 n6318 p_16_2_d2j n6020 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21264 n6021 p_16_2_d2jbar n6318 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21263 n6454 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21262 n6017 n6318 p_16_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21261 n6006 c_16_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21260 c_16_16_s1_s p_16_16_pi2j n6006 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21259 vdd c_16_16_s1_s n6316 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21258 c_16_16_s2_s c_15_17_cout n6315 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21257 n6005 c_16_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21256 n6447 p_16_16_pi2j n6005 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21255 n6447 c_15_17_cout n6313 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21254 vdd c_16_16_a n6313 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21253 n6313 p_16_16_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21252 c_17_15_cin n6447 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21251 n6315 n6316 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21250 c_17_14_a c_16_16_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21249 c_17_13_a c_16_15_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21248 n6659 n6660 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21247 c_16_15_cout n6842 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21246 n6835 c_16_15_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21245 vdd c_16_15_b n6835 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21244 n6842 c_16_15_cin n6835 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21243 n6842 c_16_15_a n6843 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21242 n6843 c_16_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21241 c_16_15_s2_s c_16_15_cin n6659 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21240 vdd c_16_15_s1_s n6660 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21239 c_16_15_s1_s c_16_15_a n6840 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21238 n6840 c_16_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21237 n6664 p_16_2_d2j n6663 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21236 n6663 p_16_2_d2jbar n6662 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21235 n6662 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21234 vdd a_14 n6664 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21233 vdd p_16_15_t_s n6658 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21232 n6658 p_16_1_n2j c_16_15_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21231 vdd n6663 n6661 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21230 n6661 n6845 p_16_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21229 n6845 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21228 vdd n7087 n6847 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21227 n6841 p_16_1_n2j p_16_14_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21226 vdd p_16_14_t_s n6841 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21225 vdd a_12 n6849 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21224 n6848 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21223 n7089 p_16_2_d2j n6848 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21222 n6849 p_16_2_d2jbar n7089 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21221 n7087 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21220 n6847 n7089 p_16_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21219 n6839 c_16_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21218 c_16_14_s1_s p_16_14_pi2j n6839 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21217 vdd c_16_14_s1_s n7084 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21216 c_16_14_s2_s c_15_15_cout n7083 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21215 n6838 c_16_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21214 n7081 p_16_14_pi2j n6838 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21213 n7081 c_15_15_cout n6834 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21212 vdd c_16_14_a n6834 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21211 n6834 p_16_14_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21210 c_17_13_cin n7081 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21209 n7083 n7084 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21208 c_17_12_a c_16_14_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21207 c_17_11_a c_16_13_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21206 n7426 n7428 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21205 c_16_13_cout n7425 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21204 n7636 c_16_13_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21203 vdd c_16_13_b n7636 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21202 n7425 c_16_13_cin n7636 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21201 n7425 c_16_13_a n7641 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21200 n7641 c_16_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21199 c_16_13_s2_s c_16_13_cin n7426 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21198 vdd c_16_13_s1_s n7428 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21197 c_16_13_s1_s c_16_13_a n7642 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21196 n7642 c_16_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21195 n7433 p_16_2_d2j n7432 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21194 n7432 p_16_2_d2jbar n7431 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21193 n7431 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21192 vdd a_12 n7433 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21191 vdd p_16_13_t_s n7424 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21190 n7424 p_16_1_n2j c_16_13_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21189 vdd n7432 n7429 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21188 n7429 n7430 p_16_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21187 n7430 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21186 vdd n7857 n7645 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21185 n7643 p_16_1_n2j c_16_12_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21184 vdd p_16_12_t_s n7643 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21183 vdd a_10 n7647 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21182 n7646 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21181 n7859 p_16_2_d2j n7646 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21180 n7647 p_16_2_d2jbar n7859 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21179 n7857 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21178 n7645 n7859 p_16_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21177 n7640 c_16_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21176 c_16_12_s1_s c_16_12_b n7640 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21175 vdd c_16_12_s1_s n7853 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21174 c_16_12_s2_s c_15_13_cout n7639 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21173 n7638 c_16_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21172 n7847 c_16_12_b n7638 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21171 n7847 c_15_13_cout n7635 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21170 vdd c_16_12_a n7635 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21169 n7635 c_16_12_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21168 c_17_11_cin n7847 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21167 n7639 n7853 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21166 c_17_10_a c_16_12_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21165 c_17_9_a c_16_11_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21164 n8179 n8177 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21163 c_16_11_cout n8178 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21162 n8172 c_16_11_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21161 vdd p_16_11_pi2j n8172 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21160 n8178 c_16_11_cin n8172 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21159 n8178 c_16_11_a n8180 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21158 n8180 p_16_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21157 c_16_11_s2_s c_16_11_cin n8179 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21156 vdd c_16_11_s1_s n8177 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21155 c_16_11_s1_s c_16_11_a n8175 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21154 n8175 p_16_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21153 n8187 p_16_2_d2j n8186 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21152 n8186 p_16_2_d2jbar n8185 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21151 n8185 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21150 vdd a_10 n8187 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21149 vdd p_16_11_t_s n8174 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21148 n8174 p_16_1_n2j p_16_11_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21147 vdd n8186 n8183 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21146 n8183 n8184 p_16_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21145 n8184 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21144 vdd n8601 n8441 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21143 n8440 p_16_1_n2j p_16_10_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21142 vdd p_16_10_t_s n8440 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21141 vdd a_8 n8443 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21140 n8442 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21139 n8603 p_16_2_d2j n8442 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21138 n8443 p_16_2_d2jbar n8603 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21137 n8601 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21136 n8441 n8603 p_16_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21135 n8439 c_16_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21134 c_16_10_s1_s p_16_10_pi2j n8439 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21133 vdd c_16_10_s1_s n8596 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21132 c_16_10_s2_s c_15_11_cout n8437 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21131 n8438 c_16_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21130 n8590 p_16_10_pi2j n8438 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21129 n8590 c_15_11_cout n8436 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21128 vdd c_16_10_a n8436 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21127 n8436 p_16_10_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21126 c_17_9_cin n8590 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21125 n8437 n8596 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21124 c_17_8_a c_16_10_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21123 c_17_7_a c_16_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21122 n8922 n8920 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21121 c_16_9_cout n8924 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21120 n8914 c_16_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21119 vdd p_16_9_pi2j n8914 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21118 n8924 c_16_9_cin n8914 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21117 n8924 c_16_9_a n8923 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21116 n8923 p_16_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21115 c_16_9_s2_s c_16_9_cin n8922 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21114 vdd c_16_9_s1_s n8920 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21113 c_16_9_s1_s c_16_9_a n8921 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21112 n8921 p_16_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21111 n8929 p_16_2_d2j n8931 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21110 n8931 p_16_2_d2jbar n8930 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21109 n8930 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21108 vdd a_8 n8929 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21107 vdd p_16_9_t_s n8918 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21106 n8918 p_16_1_n2j p_16_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21105 vdd n8931 n8927 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21104 n8927 n8928 p_16_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21103 n8928 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21102 vdd n9337 n9200 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21101 n9199 p_16_1_n2j p_16_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21100 vdd p_16_8_t_s n9199 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21099 vdd a_6 n9202 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21098 n9201 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21097 n9336 p_16_2_d2j n9201 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21096 n9202 p_16_2_d2jbar n9336 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21095 n9337 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21094 n9200 n9336 p_16_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21093 n8917 c_16_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21092 c_16_8_s1_s p_16_8_pi2j n8917 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21091 vdd c_16_8_s1_s n9327 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21090 c_16_8_s2_s c_15_9_cout n9198 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21089 n8916 c_16_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21088 n9325 p_16_8_pi2j n8916 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21087 n9325 c_15_9_cout n9197 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21086 vdd c_16_8_a n9197 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21085 n9197 p_16_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21084 c_17_7_cin n9325 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21083 n9198 n9327 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21082 c_17_6_a c_16_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21081 c_17_5_a c_16_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21080 n9695 n9693 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21079 c_16_7_cout n9697 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21078 n9686 c_16_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21077 vdd p_16_7_pi2j n9686 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21076 n9697 c_16_7_cin n9686 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21075 n9697 c_16_7_a n9696 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21074 n9696 p_16_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21073 c_16_7_s2_s c_16_7_cin n9695 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21072 vdd c_16_7_s1_s n9693 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21071 c_16_7_s1_s c_16_7_a n9694 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21070 n9694 p_16_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21069 n9547 p_16_2_d2j n9698 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21068 n9698 p_16_2_d2jbar n9546 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21067 n9546 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21066 vdd a_6 n9547 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21065 vdd p_16_7_t_s n9691 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21064 n9691 p_16_1_n2j p_16_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21063 vdd n9698 n9700 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21062 n9700 n9699 p_16_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21061 n9699 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21060 vdd n10117 n9701 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21059 n9690 p_16_1_n2j p_16_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21058 vdd p_16_6_t_s n9690 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21057 vdd a_4 n9705 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21056 n9704 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21055 n10118 p_16_2_d2j n9704 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21054 n9705 p_16_2_d2jbar n10118 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21053 n10117 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21052 n9701 n10118 p_16_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21051 n9689 c_16_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21050 c_16_6_s1_s p_16_6_pi2j n9689 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21049 vdd c_16_6_s1_s n9997 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21048 c_16_6_s2_s c_15_7_cout n9996 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21047 n9688 c_16_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21046 n10110 p_16_6_pi2j n9688 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21045 n10110 c_15_7_cout n9995 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21044 vdd c_16_6_a n9995 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21043 n9995 p_16_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21042 c_17_5_cin n10110 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21041 n9996 n9997 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21040 c_17_4_a c_16_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21039 c_17_3_a c_16_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21038 n10334 n10335 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_21037 c_16_5_cout n10511 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_21036 n10503 c_16_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21035 vdd c_16_5_b n10503 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21034 n10511 c_16_5_cin n10503 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21033 n10511 c_16_5_a n10512 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21032 n10512 c_16_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21031 c_16_5_s2_s c_16_5_cin n10334 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21030 vdd c_16_5_s1_s n10335 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21029 c_16_5_s1_s c_16_5_a n10509 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21028 n10509 c_16_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21027 n10338 p_16_2_d2j n10513 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21026 n10513 p_16_2_d2jbar n10337 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21025 n10337 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21024 vdd a_4 n10338 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21023 vdd p_16_5_t_s n10333 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21022 n10333 p_16_1_n2j c_16_5_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21021 vdd n10513 n10336 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21020 n10336 n10515 p_16_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21019 n10515 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21018 vdd n10761 n10516 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21017 n10510 p_16_1_n2j p_16_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21016 vdd p_16_4_t_s n10510 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21015 vdd a_2 n10518 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21014 n10517 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_21013 n10763 p_16_2_d2j n10517 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21012 n10518 p_16_2_d2jbar n10763 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21011 n10761 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_21010 n10516 n10763 p_16_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_21009 n10507 c_16_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21008 c_16_4_s1_s p_16_4_pi2j n10507 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21007 vdd c_16_4_s1_s n10759 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_21006 c_16_4_s2_s c_15_5_cout n10757 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_21005 n10506 c_16_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21004 n10755 p_16_4_pi2j n10506 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21003 n10755 c_15_5_cout n10502 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21002 vdd c_16_4_a n10502 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21001 n10502 p_16_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_21000 c_17_3_cin n10755 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20999 n10757 n10759 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20998 c_17_2_a c_16_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20997 c_17_1_a c_16_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20996 n11091 n11093 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20995 c_16_3_cout n11090 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20994 n11301 c_16_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20993 vdd c_16_3_b n11301 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20992 n11090 c_16_3_cin n11301 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20991 n11090 c_16_3_a n11308 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20990 n11308 c_16_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20989 c_16_3_s2_s c_16_3_cin n11091 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20988 vdd c_16_3_s1_s n11093 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20987 c_16_3_s1_s c_16_3_a n11306 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20986 n11306 c_16_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20985 n11098 p_16_2_d2j n11097 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20984 n11097 p_16_2_d2jbar n11096 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20983 n11096 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20982 vdd a_2 n11098 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20981 vdd p_16_3_t_s n11089 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20980 n11089 p_16_1_n2j c_16_3_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20979 vdd n11097 n11094 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20978 n11094 n11095 p_16_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20977 n11095 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20976 vdd n11520 n11310 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20975 n11307 p_16_1_n2j c_16_2_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20974 vdd p_16_2_t_s n11307 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20973 vdd a_0 n11312 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20972 n11311 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20971 n11522 p_16_2_d2j n11311 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20970 n11312 p_16_2_d2jbar n11522 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20969 n11520 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20968 n11310 n11522 p_16_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20967 n11305 c_16_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20966 c_16_2_s1_s c_16_2_b n11305 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20965 vdd c_16_2_s1_s n11516 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20964 c_16_2_s2_s c_15_3_cout n11304 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20963 n11303 c_16_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20962 n11510 c_16_2_b n11303 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20961 n11510 c_15_3_cout n11300 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20960 vdd c_16_2_a n11300 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20959 n11300 c_16_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20958 c_17_1_cin n11510 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20957 n11304 n11516 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20956 c_16_2_sum c_16_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20955 c_16_1_sum c_16_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20954 n11835 n11833 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20953 c_16_1_cout n11837 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20952 n11829 c_16_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20951 vdd p_16_1_pi2j n11829 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20950 n11837 c_16_1_cin n11829 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20949 n11837 c_16_1_a n11836 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20948 n11836 p_16_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20947 c_16_1_s2_s c_16_1_cin n11835 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20946 vdd c_16_1_s1_s n11833 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20945 c_16_1_s1_s c_16_1_a n11834 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20944 n11834 p_16_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20943 n11845 p_16_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20942 vdd a_0 n11845 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20941 vdd p_16_1_t_s n11831 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20940 n11831 p_16_1_n2j p_16_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20939 vdd n11845 n11841 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20938 n11841 n11844 p_16_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20937 n11844 p_16_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20936 n12099 c_15_1_sum cl4_16_s1_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20935 vdd n12221 n12099 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20934 p_24 cl4_16_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20933 n12210 c_15_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20932 vdd n12221 n12210 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20931 n12209 n12210 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20930 n12205 c_15_1_cout n12098 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20929 n12098 c_15_2_sum n12205 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20928 n12097 c_15_2_sum n12098 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_20927 vdd c_15_1_cout n12097 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_20926 n12098 c_15_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20925 vdd n12221 n12098 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20924 n12204 n12205 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20923 n12096 c_15_2_sum cl4_16_s2_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20922 vdd c_15_1_cout n12096 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20921 n12200 cl4_16_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_20920 n12095 n12209 cl4_16_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20919 vdd n12200 n12095 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20918 p_25 cl4_16_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20917 n97 p_15_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20916 c_15_33_s1_s c_15_31_a n97 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20915 vdd c_15_33_s1_s n98 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20914 c_15_33_s2_s c_15_32_cin n92 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20913 n93 p_15_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20912 n91 c_15_31_a n93 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20911 n91 c_15_32_cin n90 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20910 vdd p_15_33_pi2j n90 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20909 n90 c_15_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20908 c_16_32_cin n91 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20907 n92 n98 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20906 c_16_31_a c_15_33_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20905 n103 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20904 vdd p_15_33_t_s n96 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20903 n96 p_15_1_n2j p_15_33_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20902 vdd n103 n102 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20901 n102 n100 p_15_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20900 n100 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20899 vdd n447 n295 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20898 n294 p_15_1_n2j p_15_32_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20897 vdd p_15_32_t_s n294 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20896 vdd a_30 n297 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20895 n296 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20894 n450 p_15_2_d2j n296 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20893 n297 p_15_2_d2jbar n450 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20892 n447 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20891 n295 n450 p_15_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20890 n293 c_15_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20889 c_15_32_s1_s p_15_32_pi2j n293 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20888 vdd c_15_32_s1_s n444 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20887 c_15_32_s2_s c_15_32_cin n292 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20886 n291 c_15_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20885 n439 p_15_32_pi2j n291 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20884 n439 c_15_32_cin n290 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20883 vdd c_15_31_a n290 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20882 n290 p_15_32_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20881 c_16_31_cin n439 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20880 n292 n444 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20879 c_16_30_a c_15_32_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20878 c_16_29_a c_15_31_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20877 n757 n764 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20876 c_15_31_cout n756 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20875 n753 c_15_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20874 vdd p_15_31_pi2j n753 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20873 n756 c_15_31_cin n753 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20872 n756 c_15_31_a n755 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20871 n755 p_15_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20870 c_15_31_s2_s c_15_31_cin n757 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20869 vdd c_15_31_s1_s n764 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20868 c_15_31_s1_s c_15_31_a n761 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20867 n761 p_15_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20866 n770 p_15_2_d2j n769 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20865 n769 p_15_2_d2jbar n768 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20864 n768 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20863 vdd a_30 n770 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20862 vdd p_15_31_t_s n760 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20861 n760 p_15_1_n2j p_15_31_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20860 vdd n769 n766 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20859 n766 n767 p_15_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20858 n767 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20857 vdd n1192 n1017 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20856 n1016 p_15_1_n2j p_15_30_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20855 vdd p_15_30_t_s n1016 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20854 vdd a_28 n1019 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20853 n1018 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20852 n1196 p_15_2_d2j n1018 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20851 n1019 p_15_2_d2jbar n1196 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20850 n1192 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20849 n1017 n1196 p_15_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20848 n1015 c_15_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20847 c_15_30_s1_s p_15_30_pi2j n1015 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20846 vdd c_15_30_s1_s n1188 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20845 c_15_30_s2_s c_14_31_cout n1013 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20844 n1014 c_15_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20843 n1183 p_15_30_pi2j n1014 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20842 n1183 c_14_31_cout n1012 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20841 vdd c_15_30_a n1012 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20840 n1012 p_15_30_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20839 c_16_29_cin n1183 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20838 n1013 n1188 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20837 c_16_28_a c_15_30_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20836 c_16_27_a c_15_29_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20835 n1520 n1527 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20834 c_15_29_cout n1523 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20833 n1517 c_15_29_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20832 vdd p_15_29_pi2j n1517 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20831 n1523 c_15_29_cin n1517 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20830 n1523 c_15_29_a n1521 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20829 n1521 p_15_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20828 c_15_29_s2_s c_15_29_cin n1520 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20827 vdd c_15_29_s1_s n1527 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20826 c_15_29_s1_s c_15_29_a n1528 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20825 n1528 p_15_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20824 n1536 p_15_2_d2j n1534 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20823 n1534 p_15_2_d2jbar n1535 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20822 n1535 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20821 vdd a_28 n1536 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20820 vdd p_15_29_t_s n1526 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20819 n1526 p_15_1_n2j p_15_29_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20818 vdd n1534 n1532 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20817 n1532 n1533 p_15_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20816 n1533 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20815 vdd n1952 n1797 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20814 n1796 p_15_1_n2j p_15_28_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20813 vdd p_15_28_t_s n1796 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20812 vdd a_26 n1798 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20811 n1799 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20810 n1956 p_15_2_d2j n1799 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20809 n1798 p_15_2_d2jbar n1956 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20808 n1952 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20807 n1797 n1956 p_15_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20806 n1525 c_15_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20805 c_15_28_s1_s p_15_28_pi2j n1525 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20804 vdd c_15_28_s1_s n1795 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20803 c_15_28_s2_s c_14_29_cout n1794 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20802 n1519 c_15_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20801 n1945 p_15_28_pi2j n1519 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20800 n1945 c_14_29_cout n1793 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20799 vdd c_15_28_a n1793 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20798 n1793 p_15_28_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20797 c_16_27_cin n1945 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20796 n1794 n1795 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20795 c_16_26_a c_15_28_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20794 c_16_25_a c_15_27_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20793 n2156 n2331 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20792 c_15_27_cout n2335 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20791 n2329 c_15_27_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20790 vdd c_15_27_b n2329 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20789 n2335 c_15_27_cin n2329 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20788 n2335 c_15_27_a n2334 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20787 n2334 c_15_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20786 c_15_27_s2_s c_15_27_cin n2156 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20785 vdd c_15_27_s1_s n2331 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20784 c_15_27_s1_s c_15_27_a n2340 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20783 n2340 c_15_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20782 n2159 p_15_2_d2j n2342 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20781 n2342 p_15_2_d2jbar n2158 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20780 n2158 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20779 vdd a_26 n2159 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20778 vdd p_15_27_t_s n2157 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20777 n2157 p_15_1_n2j c_15_27_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20776 vdd n2342 n2344 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20775 n2344 n2343 p_15_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20774 n2343 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20773 vdd n2616 n2345 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20772 n2341 p_15_1_n2j p_15_26_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20771 vdd p_15_26_t_s n2341 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20770 vdd a_24 n2347 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20769 n2348 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20768 n2618 p_15_2_d2j n2348 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20767 n2347 p_15_2_d2jbar n2618 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20766 n2616 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20765 n2345 n2618 p_15_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20764 n2338 c_15_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20763 c_15_26_s1_s p_15_26_pi2j n2338 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20762 vdd c_15_26_s1_s n2615 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20761 c_15_26_s2_s c_14_27_cout n2613 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20760 n2333 c_15_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20759 n2772 p_15_26_pi2j n2333 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20758 n2772 c_14_27_cout n2612 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20757 vdd c_15_26_a n2612 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20756 n2612 p_15_26_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20755 c_16_25_cin n2772 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20754 n2613 n2615 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20753 c_16_24_a c_15_26_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20752 c_16_23_a c_15_25_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20751 n2964 n2968 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20750 c_15_25_cout n3151 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20749 n3148 c_15_25_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20748 vdd c_15_25_b n3148 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20747 n3151 c_15_25_cin n3148 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20746 n3151 c_15_25_a n3152 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20745 n3152 c_15_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20744 c_15_25_s2_s c_15_25_cin n2964 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20743 vdd c_15_25_s1_s n2968 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20742 c_15_25_s1_s c_15_25_a n3158 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20741 n3158 c_15_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20740 n2972 p_15_2_d2j n2971 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20739 n2971 p_15_2_d2jbar n2970 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20738 n2970 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20737 vdd a_24 n2972 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20736 vdd p_15_25_t_s n2967 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20735 n2967 p_15_1_n2j c_15_25_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20734 vdd n2971 n2969 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20733 n2969 n3159 p_15_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20732 n3159 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20731 vdd n3393 n3161 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20730 n3156 p_15_1_n2j c_15_24_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20729 vdd p_15_24_t_s n3156 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20728 vdd a_22 n3163 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20727 n3162 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20726 n3395 p_15_2_d2j n3162 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20725 n3163 p_15_2_d2jbar n3395 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20724 n3393 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20723 n3161 n3395 p_15_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20722 n3155 c_15_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20721 c_15_24_s1_s c_15_24_b n3155 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20720 vdd c_15_24_s1_s n3390 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20719 c_15_24_s2_s c_14_25_cout n3387 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20718 n3150 c_15_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20717 n3386 c_15_24_b n3150 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20716 n3386 c_14_25_cout n3149 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20715 vdd c_15_24_a n3149 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20714 n3149 c_15_24_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20713 c_16_23_cin n3386 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20712 n3387 n3390 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20711 c_16_22_a c_15_24_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20710 c_16_21_a c_15_23_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20709 n3739 n3747 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20708 c_15_23_cout n3741 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20707 n3979 c_15_23_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20706 vdd c_15_23_b n3979 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20705 n3741 c_15_23_cin n3979 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20704 n3741 c_15_23_a n3740 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20703 n3740 c_15_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20702 c_15_23_s2_s c_15_23_cin n3739 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20701 vdd c_15_23_s1_s n3747 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20700 c_15_23_s1_s c_15_23_a n3748 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20699 n3748 c_15_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20698 n3754 p_15_2_d2j n3753 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20697 n3753 p_15_2_d2jbar n3752 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20696 n3752 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20695 vdd a_22 n3754 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20694 vdd p_15_23_t_s n3745 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20693 n3745 p_15_1_n2j c_15_23_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20692 vdd n3753 n3750 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20691 n3750 n3751 p_15_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20690 n3751 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20689 vdd n4179 n3986 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20688 n3985 p_15_1_n2j p_15_22_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20687 vdd p_15_22_t_s n3985 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20686 vdd a_20 n3988 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20685 n3987 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20684 n4182 p_15_2_d2j n3987 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20683 n3988 p_15_2_d2jbar n4182 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20682 n4179 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20681 n3986 n4182 p_15_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20680 n3984 c_15_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20679 c_15_22_s1_s p_15_22_pi2j n3984 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20678 vdd c_15_22_s1_s n4175 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20677 c_15_22_s2_s c_14_23_cout n3982 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20676 n3981 c_15_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20675 n4170 p_15_22_pi2j n3981 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20674 n4170 c_14_23_cout n3980 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20673 vdd c_15_22_a n3980 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20672 n3980 p_15_22_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20671 c_16_21_cin n4170 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20670 n3982 n4175 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20669 c_16_20_a c_15_22_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20668 c_16_19_a c_15_21_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20667 n4503 n4511 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20666 c_15_21_cout n4504 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20665 n4500 c_15_21_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20664 vdd p_15_21_pi2j n4500 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20663 n4504 c_15_21_cin n4500 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20662 n4504 c_15_21_a n4502 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20661 n4502 p_15_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20660 c_15_21_s2_s c_15_21_cin n4503 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20659 vdd c_15_21_s1_s n4511 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20658 c_15_21_s1_s c_15_21_a n4508 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20657 n4508 p_15_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20656 n4517 p_15_2_d2j n4516 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20655 n4516 p_15_2_d2jbar n4515 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20654 n4515 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20653 vdd a_20 n4517 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20652 vdd p_15_21_t_s n4507 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20651 n4507 p_15_1_n2j p_15_21_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20650 vdd n4516 n4513 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20649 n4513 n4514 p_15_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20648 n4514 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20647 vdd n4925 n4760 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20646 n4759 p_15_1_n2j p_15_20_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20645 vdd p_15_20_t_s n4759 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20644 vdd a_18 n4762 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20643 n4761 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20642 n4928 p_15_2_d2j n4761 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20641 n4762 p_15_2_d2jbar n4928 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20640 n4925 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20639 n4760 n4928 p_15_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20638 n4758 c_15_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20637 c_15_20_s1_s p_15_20_pi2j n4758 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20636 vdd c_15_20_s1_s n4921 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20635 c_15_20_s2_s c_14_21_cout n4756 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20634 n4757 c_15_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20633 n4918 p_15_20_pi2j n4757 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20632 n4918 c_14_21_cout n4755 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20631 vdd c_15_20_a n4755 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20630 n4755 p_15_20_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20629 c_16_19_cin n4918 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20628 n4756 n4921 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20627 c_16_18_a c_15_20_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20626 c_16_17_a c_15_19_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20625 n5248 n5257 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20624 c_15_19_cout n5249 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20623 n5244 c_15_19_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20622 vdd p_15_19_pi2j n5244 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20621 n5249 c_15_19_cin n5244 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20620 n5249 c_15_19_a n5247 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20619 n5247 p_15_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20618 c_15_19_s2_s c_15_19_cin n5248 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20617 vdd c_15_19_s1_s n5257 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20616 c_15_19_s1_s c_15_19_a n5254 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20615 n5254 p_15_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20614 n5263 p_15_2_d2j n5261 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20613 n5261 p_15_2_d2jbar n5262 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20612 n5262 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20611 vdd a_18 n5263 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20610 vdd p_15_19_t_s n5253 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20609 n5253 p_15_1_n2j p_15_19_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20608 vdd n5261 n5259 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20607 n5259 n5260 p_15_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20606 n5260 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20605 vdd n5678 n5523 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20604 n5522 p_15_1_n2j p_15_18_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20603 vdd p_15_18_t_s n5522 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20602 vdd a_16 n5525 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20601 n5524 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20600 n5681 p_15_2_d2j n5524 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20599 n5525 p_15_2_d2jbar n5681 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20598 n5678 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20597 n5523 n5681 p_15_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20596 n5252 c_15_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20595 c_15_18_s1_s p_15_18_pi2j n5252 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20594 vdd c_15_18_s1_s n5521 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20593 c_15_18_s2_s c_14_19_cout n5520 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20592 n5246 c_15_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20591 n5672 p_15_18_pi2j n5246 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20590 n5672 c_14_19_cout n5519 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20589 vdd c_15_18_a n5519 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20588 n5519 p_15_18_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20587 c_16_17_cin n5672 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20586 n5520 n5521 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20585 c_16_16_a c_15_18_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20584 c_16_15_a c_15_17_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20583 n6026 n6023 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20582 c_15_17_cout n6029 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20581 n6022 c_15_17_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20580 vdd p_15_17_pi2j n6022 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20579 n6029 c_15_17_cin n6022 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20578 n6029 c_15_17_a n6027 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20577 n6027 p_15_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20576 c_15_17_s2_s c_15_17_cin n6026 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20575 vdd c_15_17_s1_s n6023 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20574 c_15_17_s1_s c_15_17_a n6035 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20573 n6035 p_15_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20572 n5874 p_15_2_d2j n6037 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20571 n6037 p_15_2_d2jbar n5873 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20570 n5873 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20569 vdd a_16 n5874 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20568 vdd p_15_17_t_s n6033 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20567 n6033 p_15_1_n2j p_15_17_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20566 vdd n6037 n6039 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20565 n6039 n6038 p_15_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20564 n6038 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20563 vdd n6468 n6040 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20562 n6032 p_15_1_n2j c_15_16_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20561 vdd p_15_16_t_s n6032 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20560 vdd a_14 n6043 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20559 n6042 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20558 n6325 p_15_2_d2j n6042 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20557 n6043 p_15_2_d2jbar n6325 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20556 n6468 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20555 n6040 n6325 p_15_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20554 n6031 c_15_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20553 c_15_16_s1_s c_15_16_b n6031 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20552 vdd c_15_16_s1_s n6323 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20551 c_15_16_s2_s c_14_17_cout n6321 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20550 n6025 c_15_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20549 n6462 c_15_16_b n6025 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20548 n6462 c_14_17_cout n6320 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20547 vdd c_15_16_a n6320 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20546 n6320 c_15_16_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20545 c_16_15_cin n6462 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20544 n6321 n6323 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20543 c_16_14_a c_15_16_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20542 c_16_13_a c_15_15_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20541 n6665 n6669 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20540 c_15_15_cout n6854 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20539 n6851 c_15_15_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20538 vdd c_15_15_b n6851 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20537 n6854 c_15_15_cin n6851 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20536 n6854 c_15_15_a n6853 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20535 n6853 c_15_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20534 c_15_15_s2_s c_15_15_cin n6665 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20533 vdd c_15_15_s1_s n6669 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20532 c_15_15_s1_s c_15_15_a n6859 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20531 n6859 c_15_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20530 n6673 p_15_2_d2j n6672 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20529 n6672 p_15_2_d2jbar n6671 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20528 n6671 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20527 vdd a_14 n6673 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20526 vdd p_15_15_t_s n6668 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20525 n6668 p_15_1_n2j c_15_15_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20524 vdd n6672 n6670 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20523 n6670 n6861 p_15_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20522 n6861 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20521 vdd n7097 n6863 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20520 n6860 p_15_1_n2j p_15_14_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20519 vdd p_15_14_t_s n6860 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20518 vdd a_12 n6864 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20517 n6865 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20516 n7099 p_15_2_d2j n6865 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20515 n6864 p_15_2_d2jbar n7099 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20514 n7097 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20513 n6863 n7099 p_15_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20512 n6857 c_15_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20511 c_15_14_s1_s p_15_14_pi2j n6857 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20510 vdd c_15_14_s1_s n7094 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20509 c_15_14_s2_s c_14_15_cout n7092 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20508 n6852 c_15_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20507 n7091 p_15_14_pi2j n6852 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20506 n7091 c_14_15_cout n6850 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20505 vdd c_15_14_a n6850 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20504 n6850 p_15_14_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20503 c_16_13_cin n7091 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20502 n7092 n7094 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20501 c_16_12_a c_15_14_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20500 c_16_11_a c_15_13_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20499 n7435 n7440 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20498 c_15_13_cout n7434 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20497 n7648 c_15_13_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20496 vdd c_15_13_b n7648 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20495 n7434 c_15_13_cin n7648 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20494 n7434 c_15_13_a n7652 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20493 n7652 c_15_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20492 c_15_13_s2_s c_15_13_cin n7435 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20491 vdd c_15_13_s1_s n7440 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20490 c_15_13_s1_s c_15_13_a n7656 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20489 n7656 c_15_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20488 n7446 p_15_2_d2j n7445 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20487 n7445 p_15_2_d2jbar n7444 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20486 n7444 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20485 vdd a_12 n7446 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20484 vdd p_15_13_t_s n7439 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20483 n7439 p_15_1_n2j c_15_13_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20482 vdd n7445 n7442 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20481 n7442 n7443 p_15_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20480 n7443 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20479 vdd n7869 n7658 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20478 n7655 p_15_1_n2j c_15_12_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20477 vdd p_15_12_t_s n7655 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20476 vdd a_10 n7660 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20475 n7659 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20474 n7872 p_15_2_d2j n7659 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20473 n7660 p_15_2_d2jbar n7872 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20472 n7869 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20471 n7658 n7872 p_15_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20470 n7654 c_15_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20469 c_15_12_s1_s c_15_12_b n7654 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20468 vdd c_15_12_s1_s n7866 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20467 c_15_12_s2_s c_14_13_cout n7651 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20466 n7650 c_15_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20465 n7863 c_15_12_b n7650 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20464 n7863 c_14_13_cout n7649 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20463 vdd c_15_12_a n7649 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20462 n7649 c_15_12_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20461 c_16_11_cin n7863 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20460 n7651 n7866 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20459 c_16_10_a c_15_12_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20458 c_16_9_a c_15_11_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20457 n8190 n8196 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20456 c_15_11_cout n8193 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20455 n8188 c_15_11_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20454 vdd p_15_11_pi2j n8188 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20453 n8193 c_15_11_cin n8188 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20452 n8193 c_15_11_a n8191 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20451 n8191 p_15_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20450 c_15_11_s2_s c_15_11_cin n8190 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20449 vdd c_15_11_s1_s n8196 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20448 c_15_11_s1_s c_15_11_a n8197 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20447 n8197 p_15_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20446 n8205 p_15_2_d2j n8204 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20445 n8204 p_15_2_d2jbar n8203 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20444 n8203 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20443 vdd a_10 n8205 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20442 vdd p_15_11_t_s n8195 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20441 n8195 p_15_1_n2j p_15_11_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20440 vdd n8204 n8201 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20439 n8201 n8202 p_15_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20438 n8202 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20437 vdd n8615 n8449 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20436 n8448 p_15_1_n2j p_15_10_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20435 vdd p_15_10_t_s n8448 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20434 vdd a_8 n8451 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20433 n8450 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20432 n8617 p_15_2_d2j n8450 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20431 n8451 p_15_2_d2jbar n8617 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20430 n8615 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20429 n8449 n8617 p_15_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20428 n8447 c_15_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20427 c_15_10_s1_s p_15_10_pi2j n8447 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20426 vdd c_15_10_s1_s n8610 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20425 c_15_10_s2_s c_14_11_cout n8445 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20424 n8446 c_15_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20423 n8605 p_15_10_pi2j n8446 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20422 n8605 c_14_11_cout n8444 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20421 vdd c_15_10_a n8444 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20420 n8444 p_15_10_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20419 c_16_9_cin n8605 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20418 n8445 n8610 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20417 c_16_8_a c_15_10_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20416 c_16_7_a c_15_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20415 n8936 n8945 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20414 c_15_9_cout n8937 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20413 n8932 c_15_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20412 vdd p_15_9_pi2j n8932 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20411 n8937 c_15_9_cin n8932 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20410 n8937 c_15_9_a n8935 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20409 n8935 p_15_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20408 c_15_9_s2_s c_15_9_cin n8936 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20407 vdd c_15_9_s1_s n8945 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20406 c_15_9_s1_s c_15_9_a n8942 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20405 n8942 p_15_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20404 n8951 p_15_2_d2j n8950 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20403 n8950 p_15_2_d2jbar n8949 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20402 n8949 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20401 vdd a_8 n8951 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20400 vdd p_15_9_t_s n8941 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20399 n8941 p_15_1_n2j p_15_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20398 vdd n8950 n8947 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20397 n8947 n8948 p_15_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20396 n8948 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20395 vdd n9349 n9206 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20394 n9205 p_15_1_n2j p_15_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20393 vdd p_15_8_t_s n9205 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20392 vdd a_6 n9208 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20391 n9207 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20390 n9352 p_15_2_d2j n9207 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20389 n9208 p_15_2_d2jbar n9352 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20388 n9349 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20387 n9206 n9352 p_15_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20386 n8940 c_15_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20385 c_15_8_s1_s p_15_8_pi2j n8940 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20384 vdd c_15_8_s1_s n9343 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20383 c_15_8_s2_s c_14_9_cout n9204 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20382 n8934 c_15_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20381 n9341 p_15_8_pi2j n8934 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20380 n9341 c_14_9_cout n9203 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20379 vdd c_15_8_a n9203 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20378 n9203 p_15_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20377 c_16_7_cin n9341 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20376 n9204 n9343 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20375 c_16_6_a c_15_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20374 c_16_5_a c_15_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20373 n9710 n9717 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20372 c_15_7_cout n9711 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20371 n9706 c_15_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20370 vdd p_15_7_pi2j n9706 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20369 n9711 c_15_7_cin n9706 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20368 n9711 c_15_7_a n9709 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20367 n9709 p_15_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20366 c_15_7_s2_s c_15_7_cin n9710 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20365 vdd c_15_7_s1_s n9717 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20364 c_15_7_s1_s c_15_7_a n9718 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20363 n9718 p_15_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20362 n9552 p_15_2_d2j n9721 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20361 n9721 p_15_2_d2jbar n9551 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20360 n9551 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20359 vdd a_6 n9552 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20358 vdd p_15_7_t_s n9716 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20357 n9716 p_15_1_n2j p_15_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20356 vdd n9721 n9723 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20355 n9723 n9722 p_15_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20354 n9722 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20353 vdd n10133 n9724 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20352 n9715 p_15_1_n2j c_15_6_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20351 vdd p_15_6_t_s n9715 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20350 vdd a_4 n9727 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20349 n9726 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20348 n10132 p_15_2_d2j n9726 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20347 n9727 p_15_2_d2jbar n10132 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20346 n10133 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20345 n9724 n10132 p_15_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20344 n9714 c_15_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20343 c_15_6_s1_s c_15_6_b n9714 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20342 vdd c_15_6_s1_s n10002 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20341 c_15_6_s2_s c_14_7_cout n10001 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20340 n9708 c_15_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20339 n10125 c_15_6_b n9708 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20338 n10125 c_14_7_cout n10000 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20337 vdd c_15_6_a n10000 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20336 n10000 c_15_6_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20335 c_16_5_cin n10125 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20334 n10001 n10002 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20333 c_16_4_a c_15_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20332 c_16_3_a c_15_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20331 n10340 n10343 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20330 c_15_5_cout n10523 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20329 n10519 c_15_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20328 vdd c_15_5_b n10519 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20327 n10523 c_15_5_cin n10519 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20326 n10523 c_15_5_a n10522 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20325 n10522 c_15_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20324 c_15_5_s2_s c_15_5_cin n10340 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20323 vdd c_15_5_s1_s n10343 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20322 c_15_5_s1_s c_15_5_a n10529 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20321 n10529 c_15_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20320 n10347 p_15_2_d2j n10530 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20319 n10530 p_15_2_d2jbar n10346 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20318 n10346 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20317 vdd a_4 n10347 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20316 vdd p_15_5_t_s n10344 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20315 n10344 p_15_1_n2j c_15_5_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20314 vdd n10530 n10345 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20313 n10345 n10532 p_15_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20312 n10532 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20311 vdd n10771 n10533 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20310 n10527 p_15_1_n2j p_15_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20309 vdd p_15_4_t_s n10527 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20308 vdd a_2 n10534 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20307 n10535 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20306 n10773 p_15_2_d2j n10535 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20305 n10534 p_15_2_d2jbar n10773 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20304 n10771 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20303 n10533 n10773 p_15_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20302 n10526 c_15_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20301 c_15_4_s1_s p_15_4_pi2j n10526 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20300 vdd c_15_4_s1_s n10768 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20299 c_15_4_s2_s c_14_5_cout n10766 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20298 n10521 c_15_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20297 n10765 p_15_4_pi2j n10521 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20296 n10765 c_14_5_cout n10520 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20295 vdd c_15_4_a n10520 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20294 n10520 p_15_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20293 c_16_3_cin n10765 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20292 n10766 n10768 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20291 c_16_2_a c_15_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20290 c_16_1_a c_15_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20289 n11100 n11105 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20288 c_15_3_cout n11099 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20287 n11313 c_15_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20286 vdd c_15_3_b n11313 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20285 n11099 c_15_3_cin n11313 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20284 n11099 c_15_3_a n11317 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20283 n11317 c_15_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20282 c_15_3_s2_s c_15_3_cin n11100 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20281 vdd c_15_3_s1_s n11105 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20280 c_15_3_s1_s c_15_3_a n11321 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20279 n11321 c_15_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20278 n11111 p_15_2_d2j n11110 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20277 n11110 p_15_2_d2jbar n11109 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20276 n11109 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20275 vdd a_2 n11111 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20274 vdd p_15_3_t_s n11104 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20273 n11104 p_15_1_n2j c_15_3_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20272 vdd n11110 n11107 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20271 n11107 n11108 p_15_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20270 n11108 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20269 vdd n11532 n11323 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20268 n11320 p_15_1_n2j c_15_2_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20267 vdd p_15_2_t_s n11320 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20266 vdd a_0 n11325 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20265 n11324 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20264 n11535 p_15_2_d2j n11324 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20263 n11325 p_15_2_d2jbar n11535 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20262 n11532 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20261 n11323 n11535 p_15_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20260 n11319 c_15_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20259 c_15_2_s1_s c_15_2_b n11319 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20258 vdd c_15_2_s1_s n11529 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20257 c_15_2_s2_s c_14_3_cout n11316 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20256 n11315 c_15_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20255 n11526 c_15_2_b n11315 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20254 n11526 c_14_3_cout n11314 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20253 vdd c_15_2_a n11314 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20252 n11314 c_15_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20251 c_16_1_cin n11526 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20250 n11316 n11529 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20249 c_15_2_sum c_15_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20248 c_15_1_sum c_15_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20247 n11849 n11856 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20246 c_15_1_cout n11850 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20245 n11846 c_15_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20244 vdd p_15_1_pi2j n11846 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20243 n11850 c_15_1_cin n11846 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20242 n11850 c_15_1_a n11848 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20241 n11848 p_15_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20240 c_15_1_s2_s c_15_1_cin n11849 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20239 vdd c_15_1_s1_s n11856 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20238 c_15_1_s1_s c_15_1_a n11857 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20237 n11857 p_15_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20236 n11864 p_15_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20235 vdd a_0 n11864 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20234 vdd p_15_1_t_s n11855 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20233 n11855 p_15_1_n2j p_15_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20232 vdd n11864 n11861 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20231 n11861 n11860 p_15_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20230 n11860 p_15_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20229 n12104 c_14_1_sum cl4_15_s1_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20228 vdd n12236 n12104 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20227 p_22 cl4_15_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20226 n12227 c_14_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20225 vdd n12236 n12227 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20224 n12228 n12227 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20223 n12223 c_14_1_cout n12103 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20222 n12103 c_14_2_sum n12223 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20221 n12102 c_14_2_sum n12103 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_20220 vdd c_14_1_cout n12102 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_20219 n12103 c_14_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20218 vdd n12236 n12103 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20217 n12221 n12223 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20216 n12101 c_14_2_sum cl4_15_s2_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20215 vdd c_14_1_cout n12101 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20214 n12219 cl4_15_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_20213 n12100 n12228 cl4_15_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20212 vdd n12219 n12100 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20211 p_23 cl4_15_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20210 n110 p_14_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20209 c_14_33_s1_s c_14_31_a n110 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20208 vdd c_14_33_s1_s n107 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20207 c_14_33_s2_s c_14_32_cin n108 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20206 n105 p_14_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20205 n106 c_14_31_a n105 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20204 n106 c_14_32_cin n104 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20203 vdd p_14_33_pi2j n104 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20202 n104 c_14_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20201 c_15_32_cin n106 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20200 n108 n107 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20199 c_15_31_a c_14_33_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20198 n117 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20197 vdd p_14_33_t_s n113 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20196 n113 p_14_1_n2j p_14_33_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20195 vdd n117 n114 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20194 n114 n115 p_14_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20193 n115 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20192 vdd n460 n303 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20191 n302 p_14_1_n2j p_14_32_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20190 vdd p_14_32_t_s n302 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20189 vdd a_30 n304 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20188 n305 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20187 n464 p_14_2_d2j n305 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20186 n304 p_14_2_d2jbar n464 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20185 n460 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20184 n303 n464 p_14_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20183 n301 c_14_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20182 c_14_32_s1_s p_14_32_pi2j n301 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20181 vdd c_14_32_s1_s n457 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20180 c_14_32_s2_s c_14_32_cin n300 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20179 n299 c_14_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20178 n452 p_14_32_pi2j n299 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20177 n452 c_14_32_cin n298 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20176 vdd c_14_31_a n298 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20175 n298 p_14_32_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20174 c_15_31_cin n452 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20173 n300 n457 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20172 c_15_30_a c_14_32_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20171 c_15_29_a c_14_31_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20170 n776 n775 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20169 c_14_31_cout n779 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20168 n771 c_14_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20167 vdd p_14_31_pi2j n771 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20166 n779 c_14_31_cin n771 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20165 n779 c_14_31_a n777 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20164 n777 p_14_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20163 c_14_31_s2_s c_14_31_cin n776 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20162 vdd c_14_31_s1_s n775 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20161 c_14_31_s1_s c_14_31_a n773 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20160 n773 p_14_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20159 n786 p_14_2_d2j n788 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20158 n788 p_14_2_d2jbar n787 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20157 n787 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20156 vdd a_30 n786 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20155 vdd p_14_31_t_s n782 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20154 n782 p_14_1_n2j p_14_31_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20153 vdd n788 n783 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20152 n783 n785 p_14_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20151 n785 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20150 vdd n1208 n1025 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20149 n1024 p_14_1_n2j p_14_30_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20148 vdd p_14_30_t_s n1024 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20147 vdd a_28 n1026 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20146 n1027 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20145 n1210 p_14_2_d2j n1027 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20144 n1026 p_14_2_d2jbar n1210 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20143 n1208 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20142 n1025 n1210 p_14_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20141 n1023 c_14_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20140 c_14_30_s1_s p_14_30_pi2j n1023 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20139 vdd c_14_30_s1_s n1204 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20138 c_14_30_s2_s c_12_31_cout n1022 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20137 n1021 c_14_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20136 n1198 p_14_30_pi2j n1021 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20135 n1198 c_12_31_cout n1020 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20134 vdd c_14_30_a n1020 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20133 n1020 p_14_30_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20132 c_15_29_cin n1198 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20131 n1022 n1204 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20130 c_15_28_a c_14_30_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20129 c_15_27_a c_14_29_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20128 n1545 n1541 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20127 c_14_29_cout n1546 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20126 n1537 c_14_29_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20125 vdd p_14_29_pi2j n1537 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20124 n1546 c_14_29_cin n1537 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20123 n1546 c_14_29_a n1544 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20122 n1544 p_14_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20121 c_14_29_s2_s c_14_29_cin n1545 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20120 vdd c_14_29_s1_s n1541 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20119 c_14_29_s1_s c_14_29_a n1542 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20118 n1542 p_14_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20117 n1555 p_14_2_d2j n1554 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20116 n1554 p_14_2_d2jbar n1556 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20115 n1556 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20114 vdd a_28 n1555 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20113 vdd p_14_29_t_s n1550 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20112 n1550 p_14_1_n2j p_14_29_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20111 vdd n1554 n1551 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20110 n1551 n1553 p_14_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20109 n1553 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20108 vdd n1967 n1804 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20107 n1803 p_14_1_n2j p_14_28_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20106 vdd p_14_28_t_s n1803 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20105 vdd a_26 n1806 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20104 n1805 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20103 n1970 p_14_2_d2j n1805 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20102 n1806 p_14_2_d2jbar n1970 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20101 n1967 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20100 n1804 n1970 p_14_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20099 n1540 c_14_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20098 c_14_28_s1_s p_14_28_pi2j n1540 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20097 vdd c_14_28_s1_s n1802 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20096 c_14_28_s2_s c_12_29_cout n1801 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20095 n1539 c_14_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20094 n1958 p_14_28_pi2j n1539 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20093 n1958 c_12_29_cout n1800 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20092 vdd c_14_28_a n1800 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20091 n1800 p_14_28_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20090 c_15_27_cin n1958 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20089 n1801 n1802 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20088 c_15_26_a c_14_28_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20087 c_15_25_a c_14_27_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20086 n2163 n2351 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20085 c_14_27_cout n2358 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20084 n2350 c_14_27_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20083 vdd c_14_27_b n2350 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20082 n2358 c_14_27_cin n2350 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20081 n2358 c_14_27_a n2355 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20080 n2355 c_14_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20079 c_14_27_s2_s c_14_27_cin n2163 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20078 vdd c_14_27_s1_s n2351 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20077 c_14_27_s1_s c_14_27_a n2357 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20076 n2357 c_14_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20075 n2165 p_14_2_d2j n2359 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20074 n2359 p_14_2_d2jbar n2166 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20073 n2166 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20072 vdd a_26 n2165 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20071 vdd p_14_27_t_s n2164 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20070 n2164 p_14_1_n2j c_14_27_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20069 vdd n2359 n2365 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20068 n2365 n2363 p_14_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20067 n2363 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20066 vdd n2624 n2366 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20065 n2362 p_14_1_n2j p_14_26_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20064 vdd p_14_26_t_s n2362 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20063 vdd a_24 n2367 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20062 n2368 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20061 n2627 p_14_2_d2j n2368 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20060 n2367 p_14_2_d2jbar n2627 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20059 n2624 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20058 n2366 n2627 p_14_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20057 n2354 c_14_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20056 c_14_26_s1_s p_14_26_pi2j n2354 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20055 vdd c_14_26_s1_s n2623 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20054 c_14_26_s2_s c_12_27_cout n2621 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20053 n2353 c_14_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20052 n2784 p_14_26_pi2j n2353 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20051 n2784 c_12_27_cout n2620 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20050 vdd c_14_26_a n2620 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20049 n2620 p_14_26_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20048 c_15_25_cin n2784 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20047 n2621 n2623 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20046 c_15_24_a c_14_26_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20045 c_15_23_a c_14_25_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20044 n2973 n2975 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20043 c_14_25_cout n3170 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20042 n3165 c_14_25_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20041 vdd c_14_25_b n3165 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20040 n3170 c_14_25_cin n3165 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20039 n3170 c_14_25_a n3171 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20038 n3171 c_14_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20037 c_14_25_s2_s c_14_25_cin n2973 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20036 vdd c_14_25_s1_s n2975 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20035 c_14_25_s1_s c_14_25_a n3168 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20034 n3168 c_14_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20033 n2979 p_14_2_d2j n2981 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20032 n2981 p_14_2_d2jbar n2980 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20031 n2980 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20030 vdd a_24 n2979 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20029 vdd p_14_25_t_s n2977 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20028 n2977 p_14_1_n2j c_14_25_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20027 vdd n2981 n2978 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20026 n2978 n3176 p_14_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20025 n3176 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20024 vdd n3404 n3177 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20023 n3174 p_14_1_n2j c_14_24_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20022 vdd p_14_24_t_s n3174 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20021 vdd a_22 n3178 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20020 n3179 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_20019 n3407 p_14_2_d2j n3179 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20018 n3178 p_14_2_d2jbar n3407 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_20017 n3404 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20016 n3177 n3407 p_14_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_20015 n3169 c_14_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20014 c_14_24_s1_s c_14_24_b n3169 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20013 vdd c_14_24_s1_s n3401 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_20012 c_14_24_s2_s c_12_25_cout n3398 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_20011 n3166 c_14_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20010 n3397 c_14_24_b n3166 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20009 n3397 c_12_25_cout n3164 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20008 vdd c_14_24_a n3164 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20007 n3164 c_14_24_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20006 c_15_23_cin n3397 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20005 n3398 n3401 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20004 c_15_22_a c_14_24_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20003 c_15_21_a c_14_23_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_20002 n3758 n3762 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_20001 c_14_23_cout n3759 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_20000 n3989 c_14_23_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19999 vdd c_14_23_b n3989 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19998 n3759 c_14_23_cin n3989 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19997 n3759 c_14_23_a n3757 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19996 n3757 c_14_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19995 c_14_23_s2_s c_14_23_cin n3758 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19994 vdd c_14_23_s1_s n3762 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19993 c_14_23_s1_s c_14_23_a n3755 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19992 n3755 c_14_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19991 n3768 p_14_2_d2j n3770 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19990 n3770 p_14_2_d2jbar n3769 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19989 n3769 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19988 vdd a_22 n3768 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19987 vdd p_14_23_t_s n3764 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19986 n3764 p_14_1_n2j c_14_23_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19985 vdd n3770 n3765 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19984 n3765 n3767 p_14_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19983 n3767 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19982 vdd n4194 n3996 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19981 n3995 p_14_1_n2j p_14_22_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19980 vdd p_14_22_t_s n3995 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19979 vdd a_20 n3997 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19978 n3998 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19977 n4197 p_14_2_d2j n3998 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19976 n3997 p_14_2_d2jbar n4197 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19975 n4194 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19974 n3996 n4197 p_14_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19973 n3993 c_14_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19972 c_14_22_s1_s p_14_22_pi2j n3993 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19971 vdd c_14_22_s1_s n4189 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19970 c_14_22_s2_s c_12_23_cout n3992 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19969 n3991 c_14_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19968 n4184 p_14_22_pi2j n3991 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19967 n4184 c_12_23_cout n3990 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19966 vdd c_14_22_a n3990 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19965 n3990 p_14_22_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19964 c_15_21_cin n4184 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19963 n3992 n4189 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19962 c_15_20_a c_14_22_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19961 c_15_19_a c_14_21_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19960 n4525 n4520 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19959 c_14_21_cout n4524 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19958 n4518 c_14_21_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19957 vdd p_14_21_pi2j n4518 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19956 n4524 c_14_21_cin n4518 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19955 n4524 c_14_21_a n4522 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19954 n4522 p_14_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19953 c_14_21_s2_s c_14_21_cin n4525 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19952 vdd c_14_21_s1_s n4520 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19951 c_14_21_s1_s c_14_21_a n4521 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19950 n4521 p_14_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19949 n4533 p_14_2_d2j n4535 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19948 n4535 p_14_2_d2jbar n4534 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19947 n4534 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19946 vdd a_20 n4533 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19945 vdd p_14_21_t_s n4529 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19944 n4529 p_14_1_n2j p_14_21_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19943 vdd n4535 n4530 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19942 n4530 n4532 p_14_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19941 n4532 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19940 vdd n4940 n4768 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19939 n4767 p_14_1_n2j p_14_20_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19938 vdd p_14_20_t_s n4767 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19937 vdd a_18 n4769 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19936 n4770 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19935 n4943 p_14_2_d2j n4770 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19934 n4769 p_14_2_d2jbar n4943 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19933 n4940 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19932 n4768 n4943 p_14_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19931 n4766 c_14_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19930 c_14_20_s1_s p_14_20_pi2j n4766 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19929 vdd c_14_20_s1_s n4936 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19928 c_14_20_s2_s c_12_21_cout n4765 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19927 n4764 c_14_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19926 n4932 p_14_20_pi2j n4764 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19925 n4932 c_12_21_cout n4763 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19924 vdd c_14_20_a n4763 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19923 n4763 p_14_20_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19922 c_15_19_cin n4932 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19921 n4765 n4936 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19920 c_15_18_a c_14_20_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19919 c_15_17_a c_14_19_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19918 n5273 n5268 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19917 c_14_19_cout n5272 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19916 n5264 c_14_19_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19915 vdd p_14_19_pi2j n5264 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19914 n5272 c_14_19_cin n5264 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19913 n5272 c_14_19_a n5270 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19912 n5270 p_14_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19911 c_14_19_s2_s c_14_19_cin n5273 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19910 vdd c_14_19_s1_s n5268 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19909 c_14_19_s1_s c_14_19_a n5269 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19908 n5269 p_14_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19907 n5282 p_14_2_d2j n5281 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19906 n5281 p_14_2_d2jbar n5283 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19905 n5283 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19904 vdd a_18 n5282 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19903 vdd p_14_19_t_s n5277 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19902 n5277 p_14_1_n2j p_14_19_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19901 vdd n5281 n5278 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19900 n5278 n5280 p_14_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19899 n5280 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19898 vdd n5693 n5530 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19897 n5529 p_14_1_n2j p_14_18_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19896 vdd p_14_18_t_s n5529 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19895 vdd a_16 n5531 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19894 n5532 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19893 n5696 p_14_2_d2j n5532 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19892 n5531 p_14_2_d2jbar n5696 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19891 n5693 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19890 n5530 n5696 p_14_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19889 n5266 c_14_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19888 c_14_18_s1_s p_14_18_pi2j n5266 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19887 vdd c_14_18_s1_s n5528 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19886 c_14_18_s2_s c_12_19_cout n5527 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19885 n5267 c_14_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19884 n5686 p_14_18_pi2j n5267 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19883 n5686 c_12_19_cout n5526 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19882 vdd c_14_18_a n5526 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19881 n5526 p_14_18_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19880 c_15_17_cin n5686 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19879 n5527 n5528 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19878 c_15_16_a c_14_18_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19877 c_15_15_a c_14_17_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19876 n6051 n6045 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19875 c_14_17_cout n6053 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19874 n6044 c_14_17_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19873 vdd p_14_17_pi2j n6044 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19872 n6053 c_14_17_cin n6044 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19871 n6053 c_14_17_a n6052 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19870 n6052 p_14_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19869 c_14_17_s2_s c_14_17_cin n6051 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19868 vdd c_14_17_s1_s n6045 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19867 c_14_17_s1_s c_14_17_a n6049 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19866 n6049 p_14_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19865 n5878 p_14_2_d2j n6055 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19864 n6055 p_14_2_d2jbar n5879 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19863 n5879 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19862 vdd a_16 n5878 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19861 vdd p_14_17_t_s n6058 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19860 n6058 p_14_1_n2j p_14_17_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19859 vdd n6055 n6062 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19858 n6062 n6060 p_14_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19857 n6060 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19856 vdd n6481 n6063 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19855 n6057 p_14_1_n2j p_14_16_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19854 vdd p_14_16_t_s n6057 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19853 vdd a_14 n6064 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19852 n6065 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19851 n6333 p_14_2_d2j n6065 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19850 n6064 p_14_2_d2jbar n6333 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19849 n6481 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19848 n6063 n6333 p_14_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19847 n6048 c_14_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19846 c_14_16_s1_s p_14_16_pi2j n6048 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19845 vdd c_14_16_s1_s n6330 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19844 c_14_16_s2_s c_12_17_cout n6328 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19843 n6047 c_14_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19842 n6474 p_14_16_pi2j n6047 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19841 n6474 c_12_17_cout n6327 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19840 vdd c_14_16_a n6327 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19839 n6327 p_14_16_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19838 c_15_15_cin n6474 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19837 n6328 n6330 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19836 c_15_14_a c_14_16_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19835 c_15_13_a c_14_15_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19834 n6674 n6676 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19833 c_14_15_cout n6873 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19832 n6867 c_14_15_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19831 vdd c_14_15_b n6867 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19830 n6873 c_14_15_cin n6867 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19829 n6873 c_14_15_a n6870 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19828 n6870 c_14_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19827 c_14_15_s2_s c_14_15_cin n6674 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19826 vdd c_14_15_s1_s n6676 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19825 c_14_15_s1_s c_14_15_a n6871 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19824 n6871 c_14_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19823 n6680 p_14_2_d2j n6682 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19822 n6682 p_14_2_d2jbar n6681 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19821 n6681 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19820 vdd a_14 n6680 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19819 vdd p_14_15_t_s n6678 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19818 n6678 p_14_1_n2j c_14_15_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19817 vdd n6682 n6679 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19816 n6679 n6878 p_14_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19815 n6878 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19814 vdd n7107 n6879 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19813 n6876 p_14_1_n2j p_14_14_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19812 vdd p_14_14_t_s n6876 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19811 vdd a_12 n6880 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19810 n6881 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19809 n7110 p_14_2_d2j n6881 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19808 n6880 p_14_2_d2jbar n7110 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19807 n7107 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19806 n6879 n7110 p_14_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19805 n6869 c_14_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19804 c_14_14_s1_s p_14_14_pi2j n6869 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19803 vdd c_14_14_s1_s n7104 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19802 c_14_14_s2_s c_12_15_cout n7102 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19801 n6868 c_14_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19800 n7101 p_14_14_pi2j n6868 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19799 n7101 c_12_15_cout n6866 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19798 vdd c_14_14_a n6866 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19797 n6866 p_14_14_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19796 c_15_13_cin n7101 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19795 n7102 n7104 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19794 c_15_12_a c_14_14_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19793 c_15_11_a c_14_13_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19792 n7447 n7452 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19791 c_14_13_cout n7449 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19790 n7661 c_14_13_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19789 vdd c_14_13_b n7661 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19788 n7449 c_14_13_cin n7661 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19787 n7449 c_14_13_a n7665 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19786 n7665 c_14_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19785 c_14_13_s2_s c_14_13_cin n7447 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19784 vdd c_14_13_s1_s n7452 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19783 c_14_13_s1_s c_14_13_a n7666 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19782 n7666 c_14_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19781 n7457 p_14_2_d2j n7459 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19780 n7459 p_14_2_d2jbar n7458 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19779 n7458 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19778 vdd a_12 n7457 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19777 vdd p_14_13_t_s n7454 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19776 n7454 p_14_1_n2j c_14_13_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19775 vdd n7459 n7455 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19774 n7455 n7456 p_14_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19773 n7456 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19772 vdd n7883 n7671 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19771 n7669 p_14_1_n2j c_14_12_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19770 vdd p_14_12_t_s n7669 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19769 vdd a_10 n7672 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19768 n7673 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19767 n7886 p_14_2_d2j n7673 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19766 n7672 p_14_2_d2jbar n7886 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19765 n7883 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19764 n7671 n7886 p_14_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19763 n7667 c_14_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19762 c_14_12_s1_s c_14_12_b n7667 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19761 vdd c_14_12_s1_s n7879 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19760 c_14_12_s2_s c_12_13_cout n7664 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19759 n7663 c_14_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19758 n7876 c_14_12_b n7663 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19757 n7876 c_12_13_cout n7662 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19756 vdd c_14_12_a n7662 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19755 n7662 c_14_12_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19754 c_15_11_cin n7876 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19753 n7664 n7879 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19752 c_15_10_a c_14_12_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19751 c_15_9_a c_14_11_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19750 n8212 n8208 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19749 c_14_11_cout n8213 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19748 n8206 c_14_11_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19747 vdd p_14_11_pi2j n8206 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19746 n8213 c_14_11_cin n8206 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19745 n8213 c_14_11_a n8211 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19744 n8211 p_14_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19743 c_14_11_s2_s c_14_11_cin n8212 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19742 vdd c_14_11_s1_s n8208 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19741 c_14_11_s1_s c_14_11_a n8209 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19740 n8209 p_14_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19739 n8221 p_14_2_d2j n8223 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19738 n8223 p_14_2_d2jbar n8222 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19737 n8222 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19736 vdd a_10 n8221 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19735 vdd p_14_11_t_s n8217 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19734 n8217 p_14_1_n2j p_14_11_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19733 vdd n8223 n8218 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19732 n8218 n8220 p_14_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19731 n8220 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19730 vdd n8629 n8457 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19729 n8456 p_14_1_n2j p_14_10_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19728 vdd p_14_10_t_s n8456 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19727 vdd a_8 n8458 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19726 n8459 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19725 n8632 p_14_2_d2j n8459 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19724 n8458 p_14_2_d2jbar n8632 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19723 n8629 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19722 n8457 n8632 p_14_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19721 n8455 c_14_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19720 c_14_10_s1_s p_14_10_pi2j n8455 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19719 vdd c_14_10_s1_s n8625 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19718 c_14_10_s2_s c_12_11_cout n8454 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19717 n8453 c_14_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19716 n8619 p_14_10_pi2j n8453 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19715 n8619 c_12_11_cout n8452 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19714 vdd c_14_10_a n8452 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19713 n8452 p_14_10_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19712 c_15_9_cin n8619 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19711 n8454 n8625 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19710 c_15_8_a c_14_10_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19709 c_15_7_a c_14_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19708 n8961 n8956 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19707 c_14_9_cout n8960 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19706 n8952 c_14_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19705 vdd p_14_9_pi2j n8952 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19704 n8960 c_14_9_cin n8952 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19703 n8960 c_14_9_a n8958 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19702 n8958 p_14_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19701 c_14_9_s2_s c_14_9_cin n8961 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19700 vdd c_14_9_s1_s n8956 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19699 c_14_9_s1_s c_14_9_a n8957 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19698 n8957 p_14_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19697 n8970 p_14_2_d2j n8969 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19696 n8969 p_14_2_d2jbar n8971 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19695 n8971 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19694 vdd a_8 n8970 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19693 vdd p_14_9_t_s n8965 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19692 n8965 p_14_1_n2j p_14_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19691 vdd n8969 n8966 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19690 n8966 n8968 p_14_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19689 n8968 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19688 vdd n9365 n9212 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19687 n9211 p_14_1_n2j p_14_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19686 vdd p_14_8_t_s n9211 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19685 vdd a_6 n9213 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19684 n9214 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19683 n9368 p_14_2_d2j n9214 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19682 n9213 p_14_2_d2jbar n9368 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19681 n9365 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19680 n9212 n9368 p_14_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19679 n8954 c_14_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19678 c_14_8_s1_s p_14_8_pi2j n8954 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19677 vdd c_14_8_s1_s n9359 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19676 c_14_8_s2_s c_12_9_cout n9210 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19675 n8955 c_14_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19674 n9357 p_14_8_pi2j n8955 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19673 n9357 c_12_9_cout n9209 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19672 vdd c_14_8_a n9209 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19671 n9209 p_14_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19670 c_15_7_cin n9357 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19669 n9210 n9359 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19668 c_15_6_a c_14_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19667 c_15_5_a c_14_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19666 n9736 n9732 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19665 c_14_7_cout n9737 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19664 n9728 c_14_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19663 vdd p_14_7_pi2j n9728 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19662 n9737 c_14_7_cin n9728 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19661 n9737 c_14_7_a n9735 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19660 n9735 p_14_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19659 c_14_7_s2_s c_14_7_cin n9736 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19658 vdd c_14_7_s1_s n9732 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19657 c_14_7_s1_s c_14_7_a n9733 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19656 n9733 p_14_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19655 n9556 p_14_2_d2j n9739 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19654 n9739 p_14_2_d2jbar n9557 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19653 n9557 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19652 vdd a_6 n9556 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19651 vdd p_14_7_t_s n9743 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19650 n9743 p_14_1_n2j p_14_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19649 vdd n9739 n9746 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19648 n9746 n9744 p_14_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19647 n9744 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19646 vdd n10147 n9747 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19645 n9741 p_14_1_n2j p_14_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19644 vdd p_14_6_t_s n9741 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19643 vdd a_4 n9748 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19642 n9749 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19641 n10146 p_14_2_d2j n9749 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19640 n9748 p_14_2_d2jbar n10146 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19639 n10147 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19638 n9747 n10146 p_14_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19637 n9731 c_14_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19636 c_14_6_s1_s p_14_6_pi2j n9731 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19635 vdd c_14_6_s1_s n10007 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19634 c_14_6_s2_s c_12_7_cout n10006 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19633 n9730 c_14_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19632 n10139 p_14_6_pi2j n9730 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19631 n10139 c_12_7_cout n10005 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19630 vdd c_14_6_a n10005 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19629 n10005 p_14_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19628 c_15_5_cin n10139 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19627 n10006 n10007 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19626 c_15_4_a c_14_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19625 c_15_3_a c_14_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19624 n10349 n10351 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19623 c_14_5_cout n10541 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19622 n10537 c_14_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19621 vdd c_14_5_b n10537 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19620 n10541 c_14_5_cin n10537 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19619 n10541 c_14_5_a n10542 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19618 n10542 c_14_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19617 c_14_5_s2_s c_14_5_cin n10349 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19616 vdd c_14_5_s1_s n10351 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19615 c_14_5_s1_s c_14_5_a n10539 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19614 n10539 c_14_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19613 n10355 p_14_2_d2j n10544 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19612 n10544 p_14_2_d2jbar n10356 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19611 n10356 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19610 vdd a_4 n10355 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19609 vdd p_14_5_t_s n10353 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19608 n10353 p_14_1_n2j c_14_5_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19607 vdd n10544 n10354 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19606 n10354 n10549 p_14_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19605 n10549 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19604 vdd n10781 n10550 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19603 n10547 p_14_1_n2j p_14_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19602 vdd p_14_4_t_s n10547 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19601 vdd a_2 n10551 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19600 n10552 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19599 n10784 p_14_2_d2j n10552 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19598 n10551 p_14_2_d2jbar n10784 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19597 n10781 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19596 n10550 n10784 p_14_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19595 n10540 c_14_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19594 c_14_4_s1_s p_14_4_pi2j n10540 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19593 vdd c_14_4_s1_s n10779 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19592 c_14_4_s2_s c_12_5_cout n10776 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19591 n10538 c_14_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19590 n10775 p_14_4_pi2j n10538 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19589 n10775 c_12_5_cout n10536 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19588 vdd c_14_4_a n10536 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19587 n10536 p_14_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19586 c_15_3_cin n10775 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19585 n10776 n10779 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19584 c_15_2_a c_14_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19583 c_15_1_a c_14_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19582 n11112 n11116 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19581 c_14_3_cout n11114 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19580 n11326 c_14_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19579 vdd c_14_3_b n11326 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19578 n11114 c_14_3_cin n11326 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19577 n11114 c_14_3_a n11332 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19576 n11332 c_14_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19575 c_14_3_s2_s c_14_3_cin n11112 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19574 vdd c_14_3_s1_s n11116 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19573 c_14_3_s1_s c_14_3_a n11330 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19572 n11330 c_14_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19571 n11122 p_14_2_d2j n11124 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19570 n11124 p_14_2_d2jbar n11123 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19569 n11123 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19568 vdd a_2 n11122 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19567 vdd p_14_3_t_s n11119 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19566 n11119 p_14_1_n2j c_14_3_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19565 vdd n11124 n11120 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19564 n11120 n11121 p_14_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19563 n11121 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19562 vdd n11546 n11336 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19561 n11334 p_14_1_n2j c_14_2_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19560 vdd p_14_2_t_s n11334 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19559 vdd a_0 n11337 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19558 n11338 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19557 n11549 p_14_2_d2j n11338 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19556 n11337 p_14_2_d2jbar n11549 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19555 n11546 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19554 n11336 n11549 p_14_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19553 n11331 c_14_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19552 c_14_2_s1_s c_14_2_b n11331 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19551 vdd c_14_2_s1_s n11542 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19550 c_14_2_s2_s c_12_3_cout n11329 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19549 n11328 c_14_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19548 n11539 c_14_2_b n11328 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19547 n11539 c_12_3_cout n11327 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19546 vdd c_14_2_a n11327 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19545 n11327 c_14_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19544 c_15_1_cin n11539 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19543 n11329 n11542 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19542 c_14_2_sum c_14_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19541 c_14_1_sum c_14_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19540 n11872 n11867 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19539 c_14_1_cout n11871 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19538 n11865 c_14_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19537 vdd p_14_1_pi2j n11865 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19536 n11871 c_14_1_cin n11865 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19535 n11871 c_14_1_a n11869 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19534 n11869 p_14_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19533 c_14_1_s2_s c_14_1_cin n11872 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19532 vdd c_14_1_s1_s n11867 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19531 c_14_1_s1_s c_14_1_a n11868 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19530 n11868 p_14_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19529 n11883 p_14_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19528 vdd a_0 n11883 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19527 vdd p_14_1_t_s n11877 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19526 n11877 p_14_1_n2j p_14_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19525 vdd n11883 n11879 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19524 n11879 n11880 p_14_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19523 n11880 p_14_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19522 n12109 c_12_1_sum cl4_14_s1_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19521 vdd n12255 n12109 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19520 p_20 cl4_14_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19519 n12244 c_12_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19518 vdd n12255 n12244 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19517 n12243 n12244 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19516 n12239 c_12_1_cout n12108 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19515 n12108 c_12_2_sum n12239 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19514 n12107 c_12_2_sum n12108 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_19513 vdd c_12_1_cout n12107 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_19512 n12108 c_12_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19511 vdd n12255 n12108 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19510 n12236 n12239 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19509 n12106 c_12_2_sum cl4_14_s2_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19508 vdd c_12_1_cout n12106 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19507 n12235 cl4_14_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_19506 n12105 n12243 cl4_14_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19505 vdd n12235 n12105 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19504 p_21 cl4_14_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19503 n125 p_12_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19502 c_12_33_s1_s c_12_31_a n125 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19501 vdd c_12_33_s1_s n123 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19500 c_12_33_s2_s c_12_32_cin n124 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19499 n121 p_12_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19498 n122 c_12_31_a n121 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19497 n122 c_12_32_cin n119 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19496 vdd p_12_33_pi2j n119 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19495 n119 c_12_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19494 c_14_32_cin n122 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19493 n124 n123 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19492 c_14_31_a c_12_33_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19491 n131 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19490 vdd p_12_33_t_s n120 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19489 n120 p_12_1_n2j p_12_33_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19488 vdd n131 n129 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19487 n129 n130 p_12_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19486 n130 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19485 vdd n474 n311 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19484 n310 p_12_1_n2j p_12_32_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19483 vdd p_12_32_t_s n310 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19482 vdd a_30 n313 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19481 n312 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19480 n477 p_12_2_d2j n312 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19479 n313 p_12_2_d2jbar n477 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19478 n474 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19477 n311 n477 p_12_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19476 n309 c_12_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19475 c_12_32_s1_s p_12_32_pi2j n309 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19474 vdd c_12_32_s1_s n470 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19473 c_12_32_s2_s c_12_32_cin n308 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19472 n307 c_12_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19471 n467 p_12_32_pi2j n307 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19470 n467 c_12_32_cin n306 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19469 vdd c_12_31_a n306 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19468 n306 p_12_32_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19467 c_14_31_cin n467 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19466 n308 n470 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19465 c_14_30_a c_12_32_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19464 c_14_29_a c_12_31_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19463 n798 n794 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19462 c_12_31_cout n799 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19461 n791 c_12_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19460 vdd p_12_31_pi2j n791 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19459 n799 c_12_31_cin n791 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19458 n799 c_12_31_a n797 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19457 n797 p_12_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19456 c_12_31_s2_s c_12_31_cin n798 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19455 vdd c_12_31_s1_s n794 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19454 c_12_31_s1_s c_12_31_a n795 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19453 n795 p_12_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19452 n806 p_12_2_d2j n805 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19451 n805 p_12_2_d2jbar n804 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19450 n804 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19449 vdd a_30 n806 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19448 vdd p_12_31_t_s n793 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19447 n793 p_12_1_n2j p_12_31_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19446 vdd n805 n802 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19445 n802 n803 p_12_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19444 n803 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19443 vdd n1223 n1033 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19442 n1032 p_12_1_n2j p_12_30_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19441 vdd p_12_30_t_s n1032 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19440 vdd a_28 n1035 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19439 n1034 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19438 n1226 p_12_2_d2j n1034 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19437 n1035 p_12_2_d2jbar n1226 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19436 n1223 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19435 n1033 n1226 p_12_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19434 n1031 c_12_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19433 c_12_30_s1_s p_12_30_pi2j n1031 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19432 vdd c_12_30_s1_s n1218 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19431 c_12_30_s2_s c_11_31_cout n1029 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19430 n1030 c_12_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19429 n1215 p_12_30_pi2j n1030 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19428 n1215 c_11_31_cout n1028 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19427 vdd c_12_30_a n1028 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19426 n1028 p_12_30_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19425 c_14_29_cin n1215 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19424 n1029 n1218 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19423 c_14_28_a c_12_30_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19422 c_14_27_a c_12_29_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19421 n1567 n1566 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19420 c_12_29_cout n1569 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19419 n1559 c_12_29_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19418 vdd p_12_29_pi2j n1559 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19417 n1569 c_12_29_cin n1559 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19416 n1569 c_12_29_a n1568 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19415 n1568 p_12_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19414 c_12_29_s2_s c_12_29_cin n1567 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19413 vdd c_12_29_s1_s n1566 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19412 c_12_29_s1_s c_12_29_a n1563 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19411 n1563 p_12_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19410 n1574 p_12_2_d2j n1576 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19409 n1576 p_12_2_d2jbar n1575 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19408 n1575 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19407 vdd a_28 n1574 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19406 vdd p_12_29_t_s n1564 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19405 n1564 p_12_1_n2j p_12_29_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19404 vdd n1576 n1571 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19403 n1571 n1573 p_12_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19402 n1573 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19401 vdd n1981 n1811 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19400 n1809 p_12_1_n2j p_12_28_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19399 vdd p_12_28_t_s n1809 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19398 vdd a_26 n1812 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19397 n1813 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19396 n1984 p_12_2_d2j n1813 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19395 n1812 p_12_2_d2jbar n1984 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19394 n1981 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19393 n1811 n1984 p_12_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19392 n1562 c_12_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19391 c_12_28_s1_s p_12_28_pi2j n1562 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19390 vdd c_12_28_s1_s n1810 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19389 c_12_28_s2_s c_11_29_cout n1808 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19388 n1561 c_12_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19387 n1975 p_12_28_pi2j n1561 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19386 n1975 c_11_29_cout n1807 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19385 vdd c_12_28_a n1807 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19384 n1807 p_12_28_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19383 c_14_27_cin n1975 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19382 n1808 n1810 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19381 c_14_26_a c_12_28_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19380 c_14_25_a c_12_27_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19379 n2171 n2372 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19378 c_12_27_cout n2380 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19377 n2371 c_12_27_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19376 vdd c_12_27_b n2371 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19375 n2380 c_12_27_cin n2371 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19374 n2380 c_12_27_a n2381 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19373 n2381 c_12_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19372 c_12_27_s2_s c_12_27_cin n2171 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19371 vdd c_12_27_s1_s n2372 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19370 c_12_27_s1_s c_12_27_a n2378 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19369 n2378 c_12_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19368 n2173 p_12_2_d2j n2382 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19367 n2382 p_12_2_d2jbar n2172 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19366 n2172 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19365 vdd a_26 n2173 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19364 vdd p_12_27_t_s n2170 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19363 n2170 p_12_1_n2j c_12_27_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19362 vdd n2382 n2384 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19361 n2384 n2383 p_12_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19360 n2383 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19359 vdd n2632 n2385 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19358 n2379 p_12_1_n2j p_12_26_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19357 vdd p_12_26_t_s n2379 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19356 vdd a_24 n2388 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19355 n2387 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19354 n2634 p_12_2_d2j n2387 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19353 n2388 p_12_2_d2jbar n2634 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19352 n2632 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19351 n2385 n2634 p_12_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19350 n2376 c_12_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19349 c_12_26_s1_s p_12_26_pi2j n2376 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19348 vdd c_12_26_s1_s n2631 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19347 c_12_26_s2_s c_11_27_cout n2630 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19346 n2375 c_12_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19345 n2799 p_12_26_pi2j n2375 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19344 n2799 c_11_27_cout n2628 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19343 vdd c_12_26_a n2628 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19342 n2628 p_12_26_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19341 c_14_25_cin n2799 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19340 n2630 n2631 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19339 c_14_24_a c_12_26_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19338 c_14_23_a c_12_25_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19337 n2985 n2986 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19336 c_12_25_cout n3189 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19335 n3181 c_12_25_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19334 vdd c_12_25_b n3181 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19333 n3189 c_12_25_cin n3181 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19332 n3189 c_12_25_a n3190 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19331 n3190 c_12_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19330 c_12_25_s2_s c_12_25_cin n2985 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19329 vdd c_12_25_s1_s n2986 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19328 c_12_25_s1_s c_12_25_a n3187 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19327 n3187 c_12_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19326 n2990 p_12_2_d2j n2989 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19325 n2989 p_12_2_d2jbar n2988 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19324 n2988 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19323 vdd a_24 n2990 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19322 vdd p_12_25_t_s n2984 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19321 n2984 p_12_1_n2j c_12_25_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19320 vdd n2989 n2987 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19319 n2987 n3191 p_12_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19318 n3191 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19317 vdd n3415 n3193 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19316 n3188 p_12_1_n2j c_12_24_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19315 vdd p_12_24_t_s n3188 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19314 vdd a_22 n3195 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19313 n3194 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19312 n3417 p_12_2_d2j n3194 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19311 n3195 p_12_2_d2jbar n3417 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19310 n3415 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19309 n3193 n3417 p_12_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19308 n3185 c_12_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19307 c_12_24_s1_s c_12_24_b n3185 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19306 vdd c_12_24_s1_s n3412 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19305 c_12_24_s2_s c_11_25_cout n3411 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19304 n3184 c_12_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19303 n3408 c_12_24_b n3184 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19302 n3408 c_11_25_cout n3180 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19301 vdd c_12_24_a n3180 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19300 n3180 c_12_24_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19299 c_14_23_cin n3408 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19298 n3411 n3412 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19297 c_14_22_a c_12_24_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19296 c_14_21_a c_12_23_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19295 n3777 n3780 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19294 c_12_23_cout n3779 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19293 n4000 c_12_23_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19292 vdd c_12_23_b n4000 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19291 n3779 c_12_23_cin n4000 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19290 n3779 c_12_23_a n3778 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19289 n3778 c_12_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19288 c_12_23_s2_s c_12_23_cin n3777 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19287 vdd c_12_23_s1_s n3780 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19286 c_12_23_s1_s c_12_23_a n3774 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19285 n3774 c_12_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19284 n3786 p_12_2_d2j n3785 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19283 n3785 p_12_2_d2jbar n3784 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19282 n3784 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19281 vdd a_22 n3786 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19280 vdd p_12_23_t_s n3775 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19279 n3775 p_12_1_n2j c_12_23_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19278 vdd n3785 n3782 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19277 n3782 n3783 p_12_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19276 n3783 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19275 vdd n4208 n4006 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19274 n4005 p_12_1_n2j p_12_22_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19273 vdd p_12_22_t_s n4005 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19272 vdd a_20 n4008 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19271 n4007 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19270 n4210 p_12_2_d2j n4007 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19269 n4008 p_12_2_d2jbar n4210 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19268 n4208 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19267 n4006 n4210 p_12_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19266 n4004 c_12_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19265 c_12_22_s1_s p_12_22_pi2j n4004 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19264 vdd c_12_22_s1_s n4203 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19263 c_12_22_s2_s c_11_23_cout n4003 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19262 n4002 c_12_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19261 n4200 p_12_22_pi2j n4002 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19260 n4200 c_11_23_cout n3999 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19259 vdd c_12_22_a n3999 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19258 n3999 p_12_22_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19257 c_14_21_cin n4200 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19256 n4003 n4203 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19255 c_14_20_a c_12_22_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19254 c_14_19_a c_12_21_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19253 n4544 n4543 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19252 c_12_21_cout n4546 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19251 n4538 c_12_21_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19250 vdd p_12_21_pi2j n4538 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19249 n4546 c_12_21_cin n4538 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19248 n4546 c_12_21_a n4545 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19247 n4545 p_12_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19246 c_12_21_s2_s c_12_21_cin n4544 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19245 vdd c_12_21_s1_s n4543 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19244 c_12_21_s1_s c_12_21_a n4540 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19243 n4540 p_12_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19242 n4553 p_12_2_d2j n4552 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19241 n4552 p_12_2_d2jbar n4551 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19240 n4551 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19239 vdd a_20 n4553 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19238 vdd p_12_21_t_s n4541 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19237 n4541 p_12_1_n2j p_12_21_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19236 vdd n4552 n4549 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19235 n4549 n4550 p_12_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19234 n4550 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19233 vdd n4954 n4776 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19232 n4775 p_12_1_n2j p_12_20_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19231 vdd p_12_20_t_s n4775 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19230 vdd a_18 n4778 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19229 n4777 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19228 n4956 p_12_2_d2j n4777 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19227 n4778 p_12_2_d2jbar n4956 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19226 n4954 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19225 n4776 n4956 p_12_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19224 n4774 c_12_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19223 c_12_20_s1_s p_12_20_pi2j n4774 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19222 vdd c_12_20_s1_s n4951 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19221 c_12_20_s2_s c_11_21_cout n4772 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19220 n4773 c_12_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19219 n4946 p_12_20_pi2j n4773 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19218 n4946 c_11_21_cout n4771 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19217 vdd c_12_20_a n4771 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19216 n4771 p_12_20_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19215 c_14_19_cin n4946 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19214 n4772 n4951 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19213 c_14_18_a c_12_20_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19212 c_14_17_a c_12_19_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19211 n5294 n5292 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19210 c_12_19_cout n5296 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19209 n5286 c_12_19_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19208 vdd p_12_19_pi2j n5286 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19207 n5296 c_12_19_cin n5286 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19206 n5296 c_12_19_a n5295 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19205 n5295 p_12_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19204 c_12_19_s2_s c_12_19_cin n5294 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19203 vdd c_12_19_s1_s n5292 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19202 c_12_19_s1_s c_12_19_a n5293 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19201 n5293 p_12_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19200 n5301 p_12_2_d2j n5303 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19199 n5303 p_12_2_d2jbar n5302 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19198 n5302 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19197 vdd a_18 n5301 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19196 vdd p_12_19_t_s n5290 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19195 n5290 p_12_1_n2j p_12_19_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19194 vdd n5303 n5298 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19193 n5298 n5300 p_12_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19192 n5300 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19191 vdd n5709 n5537 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19190 n5535 p_12_1_n2j p_12_18_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19189 vdd p_12_18_t_s n5535 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19188 vdd a_16 n5539 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19187 n5538 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19186 n5708 p_12_2_d2j n5538 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19185 n5539 p_12_2_d2jbar n5708 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19184 n5709 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19183 n5537 n5708 p_12_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19182 n5289 c_12_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19181 c_12_18_s1_s p_12_18_pi2j n5289 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19180 vdd c_12_18_s1_s n5536 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19179 c_12_18_s2_s c_11_19_cout n5534 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19178 n5288 c_12_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19177 n5699 p_12_18_pi2j n5288 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19176 n5699 c_11_19_cout n5533 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19175 vdd c_12_18_a n5533 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19174 n5533 p_12_18_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19173 c_14_17_cin n5699 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19172 n5534 n5536 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19171 c_14_16_a c_12_18_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19170 c_14_15_a c_12_17_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19169 n6078 n6069 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19168 c_12_17_cout n6079 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19167 n6068 c_12_17_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19166 vdd p_12_17_pi2j n6068 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19165 n6079 c_12_17_cin n6068 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19164 n6079 c_12_17_a n6077 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19163 n6077 p_12_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19162 c_12_17_s2_s c_12_17_cin n6078 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19161 vdd c_12_17_s1_s n6069 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19160 c_12_17_s1_s c_12_17_a n6076 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19159 n6076 p_12_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19158 n5884 p_12_2_d2j n6080 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19157 n6080 p_12_2_d2jbar n5883 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19156 n5883 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19155 vdd a_16 n5884 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19154 vdd p_12_17_t_s n6073 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19153 n6073 p_12_1_n2j p_12_17_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19152 vdd n6080 n6082 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19151 n6082 n6081 p_12_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19150 n6081 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19149 vdd n6493 n6083 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19148 n6074 p_12_1_n2j p_12_16_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19147 vdd p_12_16_t_s n6074 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19146 vdd a_14 n6087 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19145 n6086 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19144 n6339 p_12_2_d2j n6086 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19143 n6087 p_12_2_d2jbar n6339 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19142 n6493 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19141 n6083 n6339 p_12_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19140 n6072 c_12_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19139 c_12_16_s1_s p_12_16_pi2j n6072 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19138 vdd c_12_16_s1_s n6337 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19137 c_12_16_s2_s c_11_17_cout n6336 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19136 n6071 c_12_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19135 n6489 p_12_16_pi2j n6071 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19134 n6489 c_11_17_cout n6334 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19133 vdd c_12_16_a n6334 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19132 n6334 p_12_16_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19131 c_14_15_cin n6489 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19130 n6336 n6337 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19129 c_14_14_a c_12_16_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19128 c_14_13_a c_12_15_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19127 n6686 n6687 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19126 c_12_15_cout n6890 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19125 n6883 c_12_15_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19124 vdd c_12_15_b n6883 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19123 n6890 c_12_15_cin n6883 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19122 n6890 c_12_15_a n6891 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19121 n6891 c_12_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19120 c_12_15_s2_s c_12_15_cin n6686 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19119 vdd c_12_15_s1_s n6687 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19118 c_12_15_s1_s c_12_15_a n6888 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19117 n6888 c_12_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19116 n6691 p_12_2_d2j n6690 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19115 n6690 p_12_2_d2jbar n6689 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19114 n6689 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19113 vdd a_14 n6691 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19112 vdd p_12_15_t_s n6685 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19111 n6685 p_12_1_n2j c_12_15_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19110 vdd n6690 n6688 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19109 n6688 n6893 p_12_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19108 n6893 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19107 vdd n7117 n6895 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19106 n6889 p_12_1_n2j p_12_14_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19105 vdd p_12_14_t_s n6889 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19104 vdd a_12 n6897 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19103 n6896 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19102 n7119 p_12_2_d2j n6896 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19101 n6897 p_12_2_d2jbar n7119 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19100 n7117 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19099 n6895 n7119 p_12_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19098 n6887 c_12_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19097 c_12_14_s1_s p_12_14_pi2j n6887 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19096 vdd c_12_14_s1_s n7114 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19095 c_12_14_s2_s c_11_15_cout n7113 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19094 n6886 c_12_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19093 n7111 p_12_14_pi2j n6886 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19092 n7111 c_11_15_cout n6882 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19091 vdd c_12_14_a n6882 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19090 n6882 p_12_14_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19089 c_14_13_cin n7111 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19088 n7113 n7114 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19087 c_14_12_a c_12_14_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19086 c_14_11_a c_12_13_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19085 n7465 n7467 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19084 c_12_13_cout n7464 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19083 n7675 c_12_13_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19082 vdd c_12_13_b n7675 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19081 n7464 c_12_13_cin n7675 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19080 n7464 c_12_13_a n7680 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19079 n7680 c_12_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19078 c_12_13_s2_s c_12_13_cin n7465 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19077 vdd c_12_13_s1_s n7467 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19076 c_12_13_s1_s c_12_13_a n7681 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19075 n7681 c_12_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19074 n7472 p_12_2_d2j n7471 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19073 n7471 p_12_2_d2jbar n7470 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19072 n7470 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19071 vdd a_12 n7472 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19070 vdd p_12_13_t_s n7463 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19069 n7463 p_12_1_n2j c_12_13_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19068 vdd n7471 n7468 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19067 n7468 n7469 p_12_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19066 n7469 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19065 vdd n7896 n7684 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19064 n7682 p_12_1_n2j c_12_12_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19063 vdd p_12_12_t_s n7682 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19062 vdd a_10 n7686 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19061 n7685 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19060 n7898 p_12_2_d2j n7685 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19059 n7686 p_12_2_d2jbar n7898 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19058 n7896 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19057 n7684 n7898 p_12_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19056 n7679 c_12_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19055 c_12_12_s1_s c_12_12_b n7679 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19054 vdd c_12_12_s1_s n7892 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19053 c_12_12_s2_s c_11_13_cout n7678 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19052 n7677 c_12_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19051 n7889 c_12_12_b n7677 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19050 n7889 c_11_13_cout n7674 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19049 vdd c_12_12_a n7674 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19048 n7674 c_12_12_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19047 c_14_11_cin n7889 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19046 n7678 n7892 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19045 c_14_10_a c_12_12_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19044 c_14_9_a c_12_11_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19043 n8233 n8231 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19042 c_12_11_cout n8232 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19041 n8226 c_12_11_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19040 vdd p_12_11_pi2j n8226 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19039 n8232 c_12_11_cin n8226 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19038 n8232 c_12_11_a n8234 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19037 n8234 p_12_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19036 c_12_11_s2_s c_12_11_cin n8233 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19035 vdd c_12_11_s1_s n8231 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19034 c_12_11_s1_s c_12_11_a n8229 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19033 n8229 p_12_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19032 n8241 p_12_2_d2j n8240 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19031 n8240 p_12_2_d2jbar n8239 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19030 n8239 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19029 vdd a_10 n8241 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19028 vdd p_12_11_t_s n8228 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19027 n8228 p_12_1_n2j p_12_11_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19026 vdd n8240 n8237 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19025 n8237 n8238 p_12_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19024 n8238 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19023 vdd n8643 n8465 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19022 n8464 p_12_1_n2j p_12_10_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19021 vdd p_12_10_t_s n8464 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19020 vdd a_8 n8467 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19019 n8466 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_19018 n8645 p_12_2_d2j n8466 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19017 n8467 p_12_2_d2jbar n8645 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_19016 n8643 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19015 n8465 n8645 p_12_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_19014 n8463 c_12_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19013 c_12_10_s1_s p_12_10_pi2j n8463 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19012 vdd c_12_10_s1_s n8638 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_19011 c_12_10_s2_s c_11_11_cout n8461 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_19010 n8462 c_12_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19009 n8635 p_12_10_pi2j n8462 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19008 n8635 c_11_11_cout n8460 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19007 vdd c_12_10_a n8460 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19006 n8460 p_12_10_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19005 c_14_9_cin n8635 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_19004 n8461 n8638 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19003 c_14_8_a c_12_10_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19002 c_14_7_a c_12_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_19001 n8982 n8980 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_19000 c_12_9_cout n8984 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18999 n8974 c_12_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18998 vdd p_12_9_pi2j n8974 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18997 n8984 c_12_9_cin n8974 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18996 n8984 c_12_9_a n8983 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18995 n8983 p_12_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18994 c_12_9_s2_s c_12_9_cin n8982 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18993 vdd c_12_9_s1_s n8980 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18992 c_12_9_s1_s c_12_9_a n8981 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18991 n8981 p_12_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18990 n8989 p_12_2_d2j n8991 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18989 n8991 p_12_2_d2jbar n8990 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18988 n8990 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18987 vdd a_8 n8989 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18986 vdd p_12_9_t_s n8978 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18985 n8978 p_12_1_n2j p_12_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18984 vdd n8991 n8986 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18983 n8986 n8988 p_12_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18982 n8988 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18981 vdd n9382 n9218 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18980 n9217 p_12_1_n2j p_12_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18979 vdd p_12_8_t_s n9217 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18978 vdd a_6 n9220 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18977 n9219 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18976 n9381 p_12_2_d2j n9219 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18975 n9220 p_12_2_d2jbar n9381 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18974 n9382 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18973 n9218 n9381 p_12_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18972 n8977 c_12_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18971 c_12_8_s1_s p_12_8_pi2j n8977 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18970 vdd c_12_8_s1_s n9369 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18969 c_12_8_s2_s c_11_9_cout n9216 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18968 n8976 c_12_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18967 n9372 p_12_8_pi2j n8976 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18966 n9372 c_11_9_cout n9215 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18965 vdd c_12_8_a n9215 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18964 n9215 p_12_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18963 c_14_7_cin n9372 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18962 n9216 n9369 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18961 c_14_6_a c_12_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18960 c_14_5_a c_12_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18959 n9761 n9759 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18958 c_12_7_cout n9763 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18957 n9752 c_12_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18956 vdd p_12_7_pi2j n9752 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18955 n9763 c_12_7_cin n9752 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18954 n9763 c_12_7_a n9762 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18953 n9762 p_12_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18952 c_12_7_s2_s c_12_7_cin n9761 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18951 vdd c_12_7_s1_s n9759 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18950 c_12_7_s1_s c_12_7_a n9760 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18949 n9760 p_12_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18948 n9562 p_12_2_d2j n9765 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18947 n9765 p_12_2_d2jbar n9561 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18946 n9561 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18945 vdd a_6 n9562 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18944 vdd p_12_7_t_s n9757 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18943 n9757 p_12_1_n2j p_12_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18942 vdd n9765 n9766 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18941 n9766 n9764 p_12_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18940 n9764 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18939 vdd n10159 n9767 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18938 n9756 p_12_1_n2j p_12_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18937 vdd p_12_6_t_s n9756 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18936 vdd a_4 n9771 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18935 n9770 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18934 n10160 p_12_2_d2j n9770 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18933 n9771 p_12_2_d2jbar n10160 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18932 n10159 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18931 n9767 n10160 p_12_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18930 n9755 c_12_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18929 c_12_6_s1_s p_12_6_pi2j n9755 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18928 vdd c_12_6_s1_s n10012 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18927 c_12_6_s2_s c_11_7_cout n10011 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18926 n9754 c_12_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18925 n10154 p_12_6_pi2j n9754 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18924 n10154 c_11_7_cout n10010 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18923 vdd c_12_6_a n10010 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18922 n10010 p_12_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18921 c_14_5_cin n10154 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18920 n10011 n10012 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18919 c_14_4_a c_12_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18918 c_14_3_a c_12_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18917 n10361 n10362 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18916 c_12_5_cout n10562 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18915 n10554 c_12_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18914 vdd c_12_5_b n10554 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18913 n10562 c_12_5_cin n10554 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18912 n10562 c_12_5_a n10563 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18911 n10563 c_12_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18910 c_12_5_s2_s c_12_5_cin n10361 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18909 vdd c_12_5_s1_s n10362 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18908 c_12_5_s1_s c_12_5_a n10560 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18907 n10560 c_12_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18906 n10365 p_12_2_d2j n10564 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18905 n10564 p_12_2_d2jbar n10364 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18904 n10364 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18903 vdd a_4 n10365 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18902 vdd p_12_5_t_s n10360 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18901 n10360 p_12_1_n2j c_12_5_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18900 vdd n10564 n10363 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18899 n10363 n10565 p_12_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18898 n10565 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18897 vdd n10791 n10567 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18896 n10561 p_12_1_n2j p_12_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18895 vdd p_12_4_t_s n10561 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18894 vdd a_2 n10569 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18893 n10568 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18892 n10793 p_12_2_d2j n10568 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18891 n10569 p_12_2_d2jbar n10793 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18890 n10791 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18889 n10567 n10793 p_12_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18888 n10558 c_12_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18887 c_12_4_s1_s p_12_4_pi2j n10558 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18886 vdd c_12_4_s1_s n10789 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18885 c_12_4_s2_s c_11_5_cout n10787 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18884 n10557 c_12_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18883 n10785 p_12_4_pi2j n10557 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18882 n10785 c_11_5_cout n10553 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18881 vdd c_12_4_a n10553 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18880 n10553 p_12_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18879 c_14_3_cin n10785 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18878 n10787 n10789 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18877 c_14_2_a c_12_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18876 c_14_1_a c_12_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18875 n11130 n11132 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18874 c_12_3_cout n11129 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18873 n11340 c_12_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18872 vdd c_12_3_b n11340 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18871 n11129 c_12_3_cin n11340 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18870 n11129 c_12_3_a n11347 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18869 n11347 c_12_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18868 c_12_3_s2_s c_12_3_cin n11130 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18867 vdd c_12_3_s1_s n11132 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18866 c_12_3_s1_s c_12_3_a n11345 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18865 n11345 c_12_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18864 n11137 p_12_2_d2j n11136 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18863 n11136 p_12_2_d2jbar n11135 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18862 n11135 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18861 vdd a_2 n11137 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18860 vdd p_12_3_t_s n11128 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18859 n11128 p_12_1_n2j c_12_3_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18858 vdd n11136 n11133 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18857 n11133 n11134 p_12_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18856 n11134 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18855 vdd n11559 n11349 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18854 n11346 p_12_1_n2j c_12_2_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18853 vdd p_12_2_t_s n11346 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18852 vdd a_0 n11351 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18851 n11350 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18850 n11561 p_12_2_d2j n11350 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18849 n11351 p_12_2_d2jbar n11561 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18848 n11559 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18847 n11349 n11561 p_12_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18846 n11344 c_12_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18845 c_12_2_s1_s c_12_2_b n11344 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18844 vdd c_12_2_s1_s n11555 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18843 c_12_2_s2_s c_11_3_cout n11343 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18842 n11342 c_12_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18841 n11552 c_12_2_b n11342 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18840 n11552 c_11_3_cout n11339 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18839 vdd c_12_2_a n11339 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18838 n11339 c_12_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18837 c_14_1_cin n11552 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18836 n11343 n11555 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18835 c_12_2_sum c_12_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18834 c_12_1_sum c_12_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18833 n11892 n11890 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18832 c_12_1_cout n11894 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18831 n11886 c_12_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18830 vdd p_12_1_pi2j n11886 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18829 n11894 c_12_1_cin n11886 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18828 n11894 c_12_1_a n11893 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18827 n11893 p_12_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18826 c_12_1_s2_s c_12_1_cin n11892 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18825 vdd c_12_1_s1_s n11890 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18824 c_12_1_s1_s c_12_1_a n11891 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18823 n11891 p_12_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18822 n11902 p_12_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18821 vdd a_0 n11902 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18820 vdd p_12_1_t_s n11888 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18819 n11888 p_12_1_n2j p_12_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18818 vdd n11902 n11897 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18817 n11897 n11901 p_12_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18816 n11901 p_12_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18815 n12114 c_11_1_sum cl4_12_s1_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18814 vdd n12272 n12114 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18813 p_18 cl4_12_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18812 n12261 c_11_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18811 vdd n12272 n12261 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18810 n12260 n12261 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18809 n12256 c_11_1_cout n12112 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18808 n12112 c_11_2_sum n12256 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18807 n12113 c_11_2_sum n12112 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_18806 vdd c_11_1_cout n12113 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_18805 n12112 c_11_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18804 vdd n12272 n12112 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18803 n12255 n12256 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18802 n12111 c_11_2_sum cl4_12_s2_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18801 vdd c_11_1_cout n12111 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18800 n12252 cl4_12_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_18799 n12110 n12260 cl4_12_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18798 vdd n12252 n12110 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18797 p_19 cl4_12_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18796 n139 p_11_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18795 c_11_33_s1_s c_11_31_a n139 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18794 vdd c_11_33_s1_s n141 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18793 c_11_33_s2_s c_11_32_cin n134 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18792 n135 p_11_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18791 n133 c_11_31_a n135 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18790 n133 c_11_32_cin n132 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18789 vdd p_11_33_pi2j n132 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18788 n132 c_11_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18787 c_12_32_cin n133 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18786 n134 n141 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18785 c_12_31_a c_11_33_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18784 n145 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18783 vdd p_11_33_t_s n137 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18782 n137 p_11_1_n2j p_11_33_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18781 vdd n145 n144 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18780 n144 n142 p_11_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18779 n142 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18778 vdd n486 n319 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18777 n318 p_11_1_n2j p_11_32_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18776 vdd p_11_32_t_s n318 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18775 vdd a_30 n321 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18774 n320 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18773 n489 p_11_2_d2j n320 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18772 n321 p_11_2_d2jbar n489 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18771 n486 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18770 n319 n489 p_11_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18769 n317 c_11_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18768 c_11_32_s1_s p_11_32_pi2j n317 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18767 vdd c_11_32_s1_s n484 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18766 c_11_32_s2_s c_11_32_cin n316 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18765 n315 c_11_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18764 n478 p_11_32_pi2j n315 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18763 n478 c_11_32_cin n314 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18762 vdd c_11_31_a n314 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18761 n314 p_11_32_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18760 c_12_31_cin n478 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18759 n316 n484 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18758 c_12_30_a c_11_32_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18757 c_12_29_a c_11_31_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18756 n811 n815 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18755 c_11_31_cout n810 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18754 n807 c_11_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18753 vdd p_11_31_pi2j n807 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18752 n810 c_11_31_cin n807 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18751 n810 c_11_31_a n809 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18750 n809 p_11_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18749 c_11_31_s2_s c_11_31_cin n811 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18748 vdd c_11_31_s1_s n815 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18747 c_11_31_s1_s c_11_31_a n816 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18746 n816 p_11_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18745 n824 p_11_2_d2j n823 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18744 n823 p_11_2_d2jbar n822 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18743 n822 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18742 vdd a_30 n824 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18741 vdd p_11_31_t_s n814 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18740 n814 p_11_1_n2j p_11_31_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18739 vdd n823 n820 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18738 n820 n821 p_11_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18737 n821 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18736 vdd n1237 n1041 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18735 n1040 p_11_1_n2j p_11_30_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18734 vdd p_11_30_t_s n1040 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18733 vdd a_28 n1043 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18732 n1042 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18731 n1241 p_11_2_d2j n1042 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18730 n1043 p_11_2_d2jbar n1241 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18729 n1237 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18728 n1041 n1241 p_11_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18727 n1039 c_11_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18726 c_11_30_s1_s p_11_30_pi2j n1039 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18725 vdd c_11_30_s1_s n1233 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18724 c_11_30_s2_s c_10_31_cout n1037 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18723 n1038 c_11_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18722 n1228 p_11_30_pi2j n1038 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18721 n1228 c_10_31_cout n1036 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18720 vdd c_11_30_a n1036 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18719 n1036 p_11_30_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18718 c_12_29_cin n1228 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18717 n1037 n1233 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18716 c_12_28_a c_11_30_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18715 c_12_27_a c_11_29_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18714 n1580 n1589 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18713 c_11_29_cout n1583 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18712 n1577 c_11_29_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18711 vdd p_11_29_pi2j n1577 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18710 n1583 c_11_29_cin n1577 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18709 n1583 c_11_29_a n1581 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18708 n1581 p_11_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18707 c_11_29_s2_s c_11_29_cin n1580 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18706 vdd c_11_29_s1_s n1589 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18705 c_11_29_s1_s c_11_29_a n1590 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18704 n1590 p_11_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18703 n1596 p_11_2_d2j n1594 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18702 n1594 p_11_2_d2jbar n1595 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18701 n1595 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18700 vdd a_28 n1596 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18699 vdd p_11_29_t_s n1587 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18698 n1587 p_11_1_n2j p_11_29_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18697 vdd n1594 n1592 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18696 n1592 n1593 p_11_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18695 n1593 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18694 vdd n1994 n1818 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18693 n1816 p_11_1_n2j p_11_28_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18692 vdd p_11_28_t_s n1816 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18691 vdd a_26 n1819 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18690 n1820 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18689 n1998 p_11_2_d2j n1820 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18688 n1819 p_11_2_d2jbar n1998 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18687 n1994 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18686 n1818 n1998 p_11_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18685 n1585 c_11_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18684 c_11_28_s1_s p_11_28_pi2j n1585 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18683 vdd c_11_28_s1_s n1817 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18682 c_11_28_s2_s c_10_29_cout n1815 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18681 n1579 c_11_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18680 n1987 p_11_28_pi2j n1579 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18679 n1987 c_10_29_cout n1814 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18678 vdd c_11_28_a n1814 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18677 n1814 p_11_28_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18676 c_12_27_cin n1987 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18675 n1815 n1817 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18674 c_12_26_a c_11_28_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18673 c_12_25_a c_11_27_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18672 n2177 n2392 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18671 c_11_27_cout n2395 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18670 n2389 c_11_27_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18669 vdd c_11_27_b n2389 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18668 n2395 c_11_27_cin n2389 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18667 n2395 c_11_27_a n2394 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18666 n2394 c_11_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18665 c_11_27_s2_s c_11_27_cin n2177 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18664 vdd c_11_27_s1_s n2392 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18663 c_11_27_s1_s c_11_27_a n2400 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18662 n2400 c_11_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18661 n2180 p_11_2_d2j n2402 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18660 n2402 p_11_2_d2jbar n2179 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18659 n2179 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18658 vdd a_26 n2180 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18657 vdd p_11_27_t_s n2178 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18656 n2178 p_11_1_n2j c_11_27_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18655 vdd n2402 n2404 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18654 n2404 n2403 p_11_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18653 n2403 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18652 vdd n2640 n2405 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18651 n2399 p_11_1_n2j p_11_26_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18650 vdd p_11_26_t_s n2399 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18649 vdd a_24 n2407 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18648 n2408 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18647 n2642 p_11_2_d2j n2408 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18646 n2407 p_11_2_d2jbar n2642 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18645 n2640 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18644 n2405 n2642 p_11_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18643 n2398 c_11_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18642 c_11_26_s1_s p_11_26_pi2j n2398 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18641 vdd c_11_26_s1_s n2639 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18640 c_11_26_s2_s c_10_27_cout n2637 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18639 n2393 c_11_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18638 n2808 p_11_26_pi2j n2393 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18637 n2808 c_10_27_cout n2636 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18636 vdd c_11_26_a n2636 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18635 n2636 p_11_26_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18634 c_12_25_cin n2808 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18633 n2637 n2639 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18632 c_12_24_a c_11_26_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18631 c_12_23_a c_11_25_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18630 n2991 n2995 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18629 c_11_25_cout n3199 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18628 n3196 c_11_25_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18627 vdd c_11_25_b n3196 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18626 n3199 c_11_25_cin n3196 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18625 n3199 c_11_25_a n3200 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18624 n3200 c_11_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18623 c_11_25_s2_s c_11_25_cin n2991 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18622 vdd c_11_25_s1_s n2995 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18621 c_11_25_s1_s c_11_25_a n3205 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18620 n3205 c_11_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18619 n2999 p_11_2_d2j n2998 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18618 n2998 p_11_2_d2jbar n2997 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18617 n2997 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18616 vdd a_24 n2999 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18615 vdd p_11_25_t_s n2994 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18614 n2994 p_11_1_n2j c_11_25_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18613 vdd n2998 n2996 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18612 n2996 n3207 p_11_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18611 n3207 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18610 vdd n3426 n3209 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18609 n3204 p_11_1_n2j c_11_24_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18608 vdd p_11_24_t_s n3204 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18607 vdd a_22 n3211 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18606 n3210 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18605 n3428 p_11_2_d2j n3210 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18604 n3211 p_11_2_d2jbar n3428 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18603 n3426 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18602 n3209 n3428 p_11_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18601 n3203 c_11_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18600 c_11_24_s1_s c_11_24_b n3203 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18599 vdd c_11_24_s1_s n3425 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18598 c_11_24_s2_s c_10_25_cout n3420 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18597 n3198 c_11_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18596 n3419 c_11_24_b n3198 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18595 n3419 c_10_25_cout n3197 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18594 vdd c_11_24_a n3197 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18593 n3197 c_11_24_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18592 c_12_23_cin n3419 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18591 n3420 n3425 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18590 c_12_22_a c_11_24_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18589 c_12_21_a c_11_23_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18588 n3787 n3796 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18587 c_11_23_cout n3789 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18586 n4009 c_11_23_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18585 vdd c_11_23_b n4009 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18584 n3789 c_11_23_cin n4009 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18583 n3789 c_11_23_a n3788 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18582 n3788 c_11_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18581 c_11_23_s2_s c_11_23_cin n3787 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18580 vdd c_11_23_s1_s n3796 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18579 c_11_23_s1_s c_11_23_a n3794 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18578 n3794 c_11_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18577 n3802 p_11_2_d2j n3801 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18576 n3801 p_11_2_d2jbar n3800 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18575 n3800 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18574 vdd a_22 n3802 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18573 vdd p_11_23_t_s n3793 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18572 n3793 p_11_1_n2j c_11_23_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18571 vdd n3801 n3798 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18570 n3798 n3799 p_11_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18569 n3799 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18568 vdd n4221 n4016 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18567 n4015 p_11_1_n2j p_11_22_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18566 vdd p_11_22_t_s n4015 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18565 vdd a_20 n4018 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18564 n4017 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18563 n4224 p_11_2_d2j n4017 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18562 n4018 p_11_2_d2jbar n4224 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18561 n4221 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18560 n4016 n4224 p_11_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18559 n4014 c_11_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18558 c_11_22_s1_s p_11_22_pi2j n4014 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18557 vdd c_11_22_s1_s n4219 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18556 c_11_22_s2_s c_10_23_cout n4012 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18555 n4011 c_11_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18554 n4212 p_11_22_pi2j n4011 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18553 n4212 c_10_23_cout n4010 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18552 vdd c_11_22_a n4010 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18551 n4010 p_11_22_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18550 c_12_21_cin n4212 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18549 n4012 n4219 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18548 c_12_20_a c_11_22_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18547 c_12_19_a c_11_21_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18546 n4557 n4563 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18545 c_11_21_cout n4558 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18544 n4554 c_11_21_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18543 vdd p_11_21_pi2j n4554 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18542 n4558 c_11_21_cin n4554 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18541 n4558 c_11_21_a n4556 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18540 n4556 p_11_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18539 c_11_21_s2_s c_11_21_cin n4557 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18538 vdd c_11_21_s1_s n4563 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18537 c_11_21_s1_s c_11_21_a n4565 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18536 n4565 p_11_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18535 n4571 p_11_2_d2j n4570 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18534 n4570 p_11_2_d2jbar n4569 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18533 n4569 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18532 vdd a_20 n4571 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18531 vdd p_11_21_t_s n4562 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18530 n4562 p_11_1_n2j p_11_21_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18529 vdd n4570 n4567 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18528 n4567 n4568 p_11_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18527 n4568 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18526 vdd n4967 n4784 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18525 n4783 p_11_1_n2j p_11_20_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18524 vdd p_11_20_t_s n4783 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18523 vdd a_18 n4786 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18522 n4785 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18521 n4970 p_11_2_d2j n4785 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18520 n4786 p_11_2_d2jbar n4970 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18519 n4967 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18518 n4784 n4970 p_11_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18517 n4782 c_11_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18516 c_11_20_s1_s p_11_20_pi2j n4782 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18515 vdd c_11_20_s1_s n4963 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18514 c_11_20_s2_s c_10_21_cout n4780 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18513 n4781 c_11_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18512 n4960 p_11_20_pi2j n4781 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18511 n4960 c_10_21_cout n4779 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18510 vdd c_11_20_a n4779 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18509 n4779 p_11_20_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18508 c_12_19_cin n4960 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18507 n4780 n4963 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18506 c_12_18_a c_11_20_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18505 c_12_17_a c_11_19_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18504 n5308 n5315 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18503 c_11_19_cout n5309 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18502 n5304 c_11_19_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18501 vdd p_11_19_pi2j n5304 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18500 n5309 c_11_19_cin n5304 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18499 n5309 c_11_19_a n5307 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18498 n5307 p_11_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18497 c_11_19_s2_s c_11_19_cin n5308 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18496 vdd c_11_19_s1_s n5315 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18495 c_11_19_s1_s c_11_19_a n5316 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18494 n5316 p_11_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18493 n5323 p_11_2_d2j n5321 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18492 n5321 p_11_2_d2jbar n5322 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18491 n5322 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18490 vdd a_18 n5323 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18489 vdd p_11_19_t_s n5313 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18488 n5313 p_11_1_n2j p_11_19_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18487 vdd n5321 n5319 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18486 n5319 n5320 p_11_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18485 n5320 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18484 vdd n5720 n5544 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18483 n5542 p_11_1_n2j p_11_18_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18482 vdd p_11_18_t_s n5542 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18481 vdd a_16 n5546 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18480 n5545 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18479 n5723 p_11_2_d2j n5545 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18478 n5546 p_11_2_d2jbar n5723 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18477 n5720 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18476 n5544 n5723 p_11_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18475 n5312 c_11_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18474 c_11_18_s1_s p_11_18_pi2j n5312 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18473 vdd c_11_18_s1_s n5543 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18472 c_11_18_s2_s c_10_19_cout n5541 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18471 n5306 c_11_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18470 n5714 p_11_18_pi2j n5306 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18469 n5714 c_10_19_cout n5540 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18468 vdd c_11_18_a n5540 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18467 n5540 p_11_18_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18466 c_12_17_cin n5714 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18465 n5541 n5543 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18464 c_12_16_a c_11_18_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18463 c_12_15_a c_11_17_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18462 n6092 n6090 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18461 c_11_17_cout n6095 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18460 n6088 c_11_17_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18459 vdd p_11_17_pi2j n6088 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18458 n6095 c_11_17_cin n6088 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18457 n6095 c_11_17_a n6093 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18456 n6093 p_11_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18455 c_11_17_s2_s c_11_17_cin n6092 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18454 vdd c_11_17_s1_s n6090 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18453 c_11_17_s1_s c_11_17_a n6101 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18452 n6101 p_11_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18451 n5889 p_11_2_d2j n6103 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18450 n6103 p_11_2_d2jbar n5888 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18449 n5888 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18448 vdd a_16 n5889 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18447 vdd p_11_17_t_s n6098 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18446 n6098 p_11_1_n2j p_11_17_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18445 vdd n6103 n6105 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18444 n6105 n6104 p_11_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18443 n6104 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18442 vdd n6507 n6106 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18441 n6099 p_11_1_n2j p_11_16_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18440 vdd p_11_16_t_s n6099 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18439 vdd a_14 n6109 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18438 n6108 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18437 n6346 p_11_2_d2j n6108 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18436 n6109 p_11_2_d2jbar n6346 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18435 n6507 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18434 n6106 n6346 p_11_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18433 n6097 c_11_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18432 c_11_16_s1_s p_11_16_pi2j n6097 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18431 vdd c_11_16_s1_s n6344 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18430 c_11_16_s2_s c_10_17_cout n6342 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18429 n6091 c_11_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18428 n6501 p_11_16_pi2j n6091 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18427 n6501 c_10_17_cout n6341 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18426 vdd c_11_16_a n6341 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18425 n6341 p_11_16_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18424 c_12_15_cin n6501 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18423 n6342 n6344 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18422 c_12_14_a c_11_16_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18421 c_12_13_a c_11_15_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18420 n6692 n6696 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18419 c_11_15_cout n6902 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18418 n6899 c_11_15_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18417 vdd c_11_15_b n6899 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18416 n6902 c_11_15_cin n6899 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18415 n6902 c_11_15_a n6901 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18414 n6901 c_11_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18413 c_11_15_s2_s c_11_15_cin n6692 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18412 vdd c_11_15_s1_s n6696 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18411 c_11_15_s1_s c_11_15_a n6908 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18410 n6908 c_11_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18409 n6700 p_11_2_d2j n6699 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18408 n6699 p_11_2_d2jbar n6698 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18407 n6698 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18406 vdd a_14 n6700 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18405 vdd p_11_15_t_s n6695 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18404 n6695 p_11_1_n2j c_11_15_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18403 vdd n6699 n6697 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18402 n6697 n6909 p_11_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18401 n6909 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18400 vdd n7127 n6911 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18399 n6906 p_11_1_n2j p_11_14_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18398 vdd p_11_14_t_s n6906 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18397 vdd a_12 n6912 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18396 n6913 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18395 n7129 p_11_2_d2j n6913 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18394 n6912 p_11_2_d2jbar n7129 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18393 n7127 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18392 n6911 n7129 p_11_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18391 n6905 c_11_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18390 c_11_14_s1_s p_11_14_pi2j n6905 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18389 vdd c_11_14_s1_s n7126 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18388 c_11_14_s2_s c_10_15_cout n7122 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18387 n6900 c_11_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18386 n7121 p_11_14_pi2j n6900 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18385 n7121 c_10_15_cout n6898 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18384 vdd c_11_14_a n6898 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18383 n6898 p_11_14_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18382 c_12_13_cin n7121 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18381 n7122 n7126 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18380 c_12_12_a c_11_14_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18379 c_12_11_a c_11_13_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18378 n7474 n7480 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18377 c_11_13_cout n7473 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18376 n7687 c_11_13_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18375 vdd c_11_13_b n7687 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18374 n7473 c_11_13_cin n7687 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18373 n7473 c_11_13_a n7691 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18372 n7691 c_11_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18371 c_11_13_s2_s c_11_13_cin n7474 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18370 vdd c_11_13_s1_s n7480 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18369 c_11_13_s1_s c_11_13_a n7694 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18368 n7694 c_11_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18367 n7485 p_11_2_d2j n7484 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18366 n7484 p_11_2_d2jbar n7483 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18365 n7483 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18364 vdd a_12 n7485 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18363 vdd p_11_13_t_s n7478 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18362 n7478 p_11_1_n2j c_11_13_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18361 vdd n7484 n7481 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18360 n7481 n7482 p_11_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18359 n7482 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18358 vdd n7908 n7697 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18357 n7695 p_11_1_n2j c_11_12_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18356 vdd p_11_12_t_s n7695 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18355 vdd a_10 n7699 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18354 n7698 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18353 n7911 p_11_2_d2j n7698 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18352 n7699 p_11_2_d2jbar n7911 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18351 n7908 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18350 n7697 n7911 p_11_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18349 n7693 c_11_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18348 c_11_12_s1_s c_11_12_b n7693 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18347 vdd c_11_12_s1_s n7907 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18346 c_11_12_s2_s c_10_13_cout n7690 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18345 n7689 c_11_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18344 n7902 c_11_12_b n7689 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18343 n7902 c_10_13_cout n7688 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18342 vdd c_11_12_a n7688 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18341 n7688 c_11_12_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18340 c_12_11_cin n7902 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18339 n7690 n7907 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18338 c_12_10_a c_11_12_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18337 c_12_9_a c_11_11_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18336 n8244 n8251 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18335 c_11_11_cout n8247 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18334 n8242 c_11_11_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18333 vdd p_11_11_pi2j n8242 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18332 n8247 c_11_11_cin n8242 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18331 n8247 c_11_11_a n8245 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18330 n8245 p_11_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18329 c_11_11_s2_s c_11_11_cin n8244 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18328 vdd c_11_11_s1_s n8251 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18327 c_11_11_s1_s c_11_11_a n8252 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18326 n8252 p_11_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18325 n8259 p_11_2_d2j n8258 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18324 n8258 p_11_2_d2jbar n8257 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18323 n8257 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18322 vdd a_10 n8259 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18321 vdd p_11_11_t_s n8250 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18320 n8250 p_11_1_n2j p_11_11_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18319 vdd n8258 n8255 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18318 n8255 n8256 p_11_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18317 n8256 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18316 vdd n8657 n8473 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18315 n8472 p_11_1_n2j p_11_10_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18314 vdd p_11_10_t_s n8472 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18313 vdd a_8 n8475 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18312 n8474 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18311 n8659 p_11_2_d2j n8474 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18310 n8475 p_11_2_d2jbar n8659 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18309 n8657 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18308 n8473 n8659 p_11_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18307 n8471 c_11_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18306 c_11_10_s1_s p_11_10_pi2j n8471 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18305 vdd c_11_10_s1_s n8653 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18304 c_11_10_s2_s c_10_11_cout n8469 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18303 n8470 c_11_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18302 n8647 p_11_10_pi2j n8470 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18301 n8647 c_10_11_cout n8468 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18300 vdd c_11_10_a n8468 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18299 n8468 p_11_10_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18298 c_12_9_cin n8647 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18297 n8469 n8653 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18296 c_12_8_a c_11_10_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18295 c_12_7_a c_11_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18294 n8996 n9003 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18293 c_11_9_cout n8997 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18292 n8992 c_11_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18291 vdd p_11_9_pi2j n8992 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18290 n8997 c_11_9_cin n8992 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18289 n8997 c_11_9_a n8995 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18288 n8995 p_11_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18287 c_11_9_s2_s c_11_9_cin n8996 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18286 vdd c_11_9_s1_s n9003 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18285 c_11_9_s1_s c_11_9_a n9004 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18284 n9004 p_11_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18283 n9011 p_11_2_d2j n9010 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18282 n9010 p_11_2_d2jbar n9009 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18281 n9009 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18280 vdd a_8 n9011 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18279 vdd p_11_9_t_s n9001 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18278 n9001 p_11_1_n2j p_11_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18277 vdd n9010 n9007 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18276 n9007 n9008 p_11_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18275 n9008 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18274 vdd n9394 n9224 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18273 n9223 p_11_1_n2j p_11_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18272 vdd p_11_8_t_s n9223 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18271 vdd a_6 n9226 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18270 n9225 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18269 n9397 p_11_2_d2j n9225 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18268 n9226 p_11_2_d2jbar n9397 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18267 n9394 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18266 n9224 n9397 p_11_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18265 n9000 c_11_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18264 c_11_8_s1_s p_11_8_pi2j n9000 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18263 vdd c_11_8_s1_s n9389 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18262 c_11_8_s2_s c_10_9_cout n9222 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18261 n8994 c_11_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18260 n9386 p_11_8_pi2j n8994 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18259 n9386 c_10_9_cout n9221 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18258 vdd c_11_8_a n9221 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18257 n9221 p_11_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18256 c_12_7_cin n9386 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18255 n9222 n9389 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18254 c_12_6_a c_11_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18253 c_12_5_a c_11_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18252 n9776 n9785 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18251 c_11_7_cout n9777 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18250 n9772 c_11_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18249 vdd p_11_7_pi2j n9772 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18248 n9777 c_11_7_cin n9772 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18247 n9777 c_11_7_a n9775 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18246 n9775 p_11_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18245 c_11_7_s2_s c_11_7_cin n9776 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18244 vdd c_11_7_s1_s n9785 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18243 c_11_7_s1_s c_11_7_a n9786 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18242 n9786 p_11_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18241 n9567 p_11_2_d2j n9787 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18240 n9787 p_11_2_d2jbar n9566 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18239 n9566 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18238 vdd a_6 n9567 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18237 vdd p_11_7_t_s n9783 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18236 n9783 p_11_1_n2j p_11_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18235 vdd n9787 n9789 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18234 n9789 n9788 p_11_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18233 n9788 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18232 vdd n10175 n9790 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18231 n9781 p_11_1_n2j c_11_6_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18230 vdd p_11_6_t_s n9781 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18229 vdd a_4 n9793 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18228 n9792 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18227 n10174 p_11_2_d2j n9792 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18226 n9793 p_11_2_d2jbar n10174 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18225 n10175 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18224 n9790 n10174 p_11_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18223 n9780 c_11_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18222 c_11_6_s1_s c_11_6_b n9780 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18221 vdd c_11_6_s1_s n10017 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18220 c_11_6_s2_s c_10_7_cout n10016 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18219 n9774 c_11_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18218 n10167 c_11_6_b n9774 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18217 n10167 c_10_7_cout n10015 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18216 vdd c_11_6_a n10015 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18215 n10015 c_11_6_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18214 c_12_5_cin n10167 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18213 n10016 n10017 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18212 c_12_4_a c_11_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18211 c_12_3_a c_11_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18210 n10367 n10371 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18209 c_11_5_cout n10574 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18208 n10570 c_11_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18207 vdd c_11_5_b n10570 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18206 n10574 c_11_5_cin n10570 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18205 n10574 c_11_5_a n10573 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18204 n10573 c_11_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18203 c_11_5_s2_s c_11_5_cin n10367 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18202 vdd c_11_5_s1_s n10371 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18201 c_11_5_s1_s c_11_5_a n10579 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18200 n10579 c_11_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18199 n10374 p_11_2_d2j n10581 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18198 n10581 p_11_2_d2jbar n10373 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18197 n10373 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18196 vdd a_4 n10374 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18195 vdd p_11_5_t_s n10370 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18194 n10370 p_11_1_n2j c_11_5_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18193 vdd n10581 n10372 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18192 n10372 n10583 p_11_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18191 n10583 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18190 vdd n10801 n10584 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18189 n10578 p_11_1_n2j p_11_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18188 vdd p_11_4_t_s n10578 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18187 vdd a_2 n10585 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18186 n10586 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18185 n10803 p_11_2_d2j n10586 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18184 n10585 p_11_2_d2jbar n10803 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18183 n10801 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18182 n10584 n10803 p_11_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18181 n10577 c_11_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18180 c_11_4_s1_s p_11_4_pi2j n10577 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18179 vdd c_11_4_s1_s n10800 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18178 c_11_4_s2_s c_10_5_cout n10796 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18177 n10572 c_11_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18176 n10795 p_11_4_pi2j n10572 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18175 n10795 c_10_5_cout n10571 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18174 vdd c_11_4_a n10571 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18173 n10571 p_11_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18172 c_12_3_cin n10795 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18171 n10796 n10800 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18170 c_12_2_a c_11_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18169 c_12_1_a c_11_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18168 n11139 n11144 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18167 c_11_3_cout n11138 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18166 n11352 c_11_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18165 vdd c_11_3_b n11352 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18164 n11138 c_11_3_cin n11352 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18163 n11138 c_11_3_a n11356 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18162 n11356 c_11_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18161 c_11_3_s2_s c_11_3_cin n11139 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18160 vdd c_11_3_s1_s n11144 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18159 c_11_3_s1_s c_11_3_a n11360 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18158 n11360 c_11_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18157 n11150 p_11_2_d2j n11149 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18156 n11149 p_11_2_d2jbar n11148 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18155 n11148 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18154 vdd a_2 n11150 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18153 vdd p_11_3_t_s n11143 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18152 n11143 p_11_1_n2j c_11_3_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18151 vdd n11149 n11146 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18150 n11146 n11147 p_11_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18149 n11147 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18148 vdd n11571 n11362 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18147 n11359 p_11_1_n2j c_11_2_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18146 vdd p_11_2_t_s n11359 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18145 vdd a_0 n11364 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18144 n11363 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18143 n11574 p_11_2_d2j n11363 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18142 n11364 p_11_2_d2jbar n11574 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18141 n11571 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18140 n11362 n11574 p_11_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18139 n11358 c_11_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18138 c_11_2_s1_s c_11_2_b n11358 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18137 vdd c_11_2_s1_s n11570 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18136 c_11_2_s2_s c_10_3_cout n11355 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18135 n11354 c_11_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18134 n11565 c_11_2_b n11354 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18133 n11565 c_10_3_cout n11353 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18132 vdd c_11_2_a n11353 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18131 n11353 c_11_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18130 c_12_1_cin n11565 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18129 n11355 n11570 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18128 c_11_2_sum c_11_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18127 c_11_1_sum c_11_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18126 n11906 n11915 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18125 c_11_1_cout n11907 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18124 n11903 c_11_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18123 vdd p_11_1_pi2j n11903 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18122 n11907 c_11_1_cin n11903 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18121 n11907 c_11_1_a n11905 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18120 n11905 p_11_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18119 c_11_1_s2_s c_11_1_cin n11906 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18118 vdd c_11_1_s1_s n11915 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18117 c_11_1_s1_s c_11_1_a n11911 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18116 n11911 p_11_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18115 n11921 p_11_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18114 vdd a_0 n11921 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18113 vdd p_11_1_t_s n11913 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18112 n11913 p_11_1_n2j p_11_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18111 vdd n11921 n11918 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18110 n11918 n11917 p_11_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18109 n11917 p_11_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18108 n12119 c_10_1_sum cl4_11_s1_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18107 vdd n12287 n12119 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18106 p_16 cl4_11_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18105 n12278 c_10_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18104 vdd n12287 n12278 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18103 n12279 n12278 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18102 n12274 c_10_1_cout n12118 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18101 n12118 c_10_2_sum n12274 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18100 n12117 c_10_2_sum n12118 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_18099 vdd c_10_1_cout n12117 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_18098 n12118 c_10_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18097 vdd n12287 n12118 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18096 n12272 n12274 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18095 n12116 c_10_2_sum cl4_11_s2_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18094 vdd c_10_1_cout n12116 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18093 n12270 cl4_11_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_18092 n12115 n12279 cl4_11_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18091 vdd n12270 n12115 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18090 p_17 cl4_11_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18089 n152 p_10_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18088 c_10_33_s1_s c_10_31_a n152 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18087 vdd c_10_33_s1_s n149 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18086 c_10_33_s2_s c_10_32_cin n150 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18085 n147 p_10_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18084 n148 c_10_31_a n147 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18083 n148 c_10_32_cin n146 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18082 vdd p_10_33_pi2j n146 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18081 n146 c_10_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18080 c_11_32_cin n148 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18079 n150 n149 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18078 c_11_31_a c_10_33_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18077 n159 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18076 vdd p_10_33_t_s n155 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18075 n155 p_10_1_n2j p_10_33_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18074 vdd n159 n158 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18073 n158 n156 p_10_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18072 n156 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18071 vdd n499 n327 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18070 n326 p_10_1_n2j p_10_32_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18069 vdd p_10_32_t_s n326 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18068 vdd a_30 n328 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18067 n329 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18066 n503 p_10_2_d2j n329 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18065 n328 p_10_2_d2jbar n503 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18064 n499 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18063 n327 n503 p_10_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18062 n325 c_10_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18061 c_10_32_s1_s p_10_32_pi2j n325 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18060 vdd c_10_32_s1_s n496 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18059 c_10_32_s2_s c_10_32_cin n324 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18058 n323 c_10_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18057 n491 p_10_32_pi2j n323 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18056 n491 c_10_32_cin n322 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18055 vdd c_10_31_a n322 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18054 n322 p_10_32_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18053 c_11_31_cin n491 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18052 n324 n496 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18051 c_11_30_a c_10_32_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18050 c_11_29_a c_10_31_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18049 n830 n829 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18048 c_10_31_cout n833 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18047 n825 c_10_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18046 vdd p_10_31_pi2j n825 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18045 n833 c_10_31_cin n825 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18044 n833 c_10_31_a n831 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18043 n831 p_10_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18042 c_10_31_s2_s c_10_31_cin n830 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18041 vdd c_10_31_s1_s n829 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18040 c_10_31_s1_s c_10_31_a n827 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18039 n827 p_10_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18038 n840 p_10_2_d2j n841 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18037 n841 p_10_2_d2jbar n842 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18036 n842 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18035 vdd a_30 n840 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18034 vdd p_10_31_t_s n836 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18033 n836 p_10_1_n2j p_10_31_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18032 vdd n841 n837 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18031 n837 n839 p_10_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18030 n839 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18029 vdd n1253 n1049 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18028 n1048 p_10_1_n2j p_10_30_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18027 vdd p_10_30_t_s n1048 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18026 vdd a_28 n1050 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18025 n1051 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_18024 n1255 p_10_2_d2j n1051 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18023 n1050 p_10_2_d2jbar n1255 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_18022 n1253 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18021 n1049 n1255 p_10_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_18020 n1047 c_10_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18019 c_10_30_s1_s p_10_30_pi2j n1047 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18018 vdd c_10_30_s1_s n1249 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_18017 c_10_30_s2_s c_9_31_cout n1046 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_18016 n1045 c_10_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18015 n1243 p_10_30_pi2j n1045 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18014 n1243 c_9_31_cout n1044 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18013 vdd c_10_30_a n1044 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18012 n1044 p_10_30_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18011 c_11_29_cin n1243 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18010 n1046 n1249 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18009 c_11_28_a c_10_30_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18008 c_11_27_a c_10_29_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18007 n1605 n1601 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_18006 c_10_29_cout n1606 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_18005 n1597 c_10_29_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18004 vdd p_10_29_pi2j n1597 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18003 n1606 c_10_29_cin n1597 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18002 n1606 c_10_29_a n1604 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18001 n1604 p_10_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_18000 c_10_29_s2_s c_10_29_cin n1605 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17999 vdd c_10_29_s1_s n1601 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17998 c_10_29_s1_s c_10_29_a n1602 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17997 n1602 p_10_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17996 n1614 p_10_2_d2j n1615 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17995 n1615 p_10_2_d2jbar n1616 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17994 n1616 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17993 vdd a_28 n1614 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17992 vdd p_10_29_t_s n1610 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17991 n1610 p_10_1_n2j p_10_29_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17990 vdd n1615 n1612 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17989 n1612 n1613 p_10_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17988 n1613 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17987 vdd n2009 n1825 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17986 n1824 p_10_1_n2j p_10_28_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17985 vdd p_10_28_t_s n1824 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17984 vdd a_26 n1827 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17983 n1826 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17982 n2011 p_10_2_d2j n1826 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17981 n1827 p_10_2_d2jbar n2011 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17980 n2009 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17979 n1825 n2011 p_10_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17978 n1600 c_10_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17977 c_10_28_s1_s p_10_28_pi2j n1600 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17976 vdd c_10_28_s1_s n1823 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17975 c_10_28_s2_s c_9_29_cout n1822 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17974 n1599 c_10_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17973 n2000 p_10_28_pi2j n1599 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17972 n2000 c_9_29_cout n1821 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17971 vdd c_10_28_a n1821 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17970 n1821 p_10_28_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17969 c_11_27_cin n2000 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17968 n1822 n1823 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17967 c_11_26_a c_10_28_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17966 c_11_25_a c_10_27_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17965 n2184 n2410 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17964 c_10_27_cout n2418 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17963 n2409 c_10_27_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17962 vdd c_10_27_b n2409 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17961 n2418 c_10_27_cin n2409 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17960 n2418 c_10_27_a n2415 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17959 n2415 c_10_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17958 c_10_27_s2_s c_10_27_cin n2184 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17957 vdd c_10_27_s1_s n2410 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17956 c_10_27_s1_s c_10_27_a n2417 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17955 n2417 c_10_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17954 n2186 p_10_2_d2j n2419 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17953 n2419 p_10_2_d2jbar n2187 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17952 n2187 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17951 vdd a_26 n2186 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17950 vdd p_10_27_t_s n2185 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17949 n2185 p_10_1_n2j c_10_27_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17948 vdd n2419 n2425 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17947 n2425 n2423 p_10_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17946 n2423 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17945 vdd n2648 n2426 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17944 n2422 p_10_1_n2j p_10_26_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17943 vdd p_10_26_t_s n2422 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17942 vdd a_24 n2428 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17941 n2427 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17940 n2650 p_10_2_d2j n2427 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17939 n2428 p_10_2_d2jbar n2650 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17938 n2648 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17937 n2426 n2650 p_10_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17936 n2414 c_10_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17935 c_10_26_s1_s p_10_26_pi2j n2414 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17934 vdd c_10_26_s1_s n2647 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17933 c_10_26_s2_s c_9_27_cout n2645 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17932 n2413 c_10_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17931 n2820 p_10_26_pi2j n2413 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17930 n2820 c_9_27_cout n2644 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17929 vdd c_10_26_a n2644 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17928 n2644 p_10_26_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17927 c_11_25_cin n2820 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17926 n2645 n2647 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17925 c_11_24_a c_10_26_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17924 c_11_23_a c_10_25_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17923 n3000 n3001 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17922 c_10_25_cout n3218 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17921 n3213 c_10_25_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17920 vdd c_10_25_b n3213 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17919 n3218 c_10_25_cin n3213 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17918 n3218 c_10_25_a n3219 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17917 n3219 c_10_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17916 c_10_25_s2_s c_10_25_cin n3000 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17915 vdd c_10_25_s1_s n3001 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17914 c_10_25_s1_s c_10_25_a n3216 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17913 n3216 c_10_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17912 n3006 p_10_2_d2j n3007 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17911 n3007 p_10_2_d2jbar n3008 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17910 n3008 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17909 vdd a_24 n3006 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17908 vdd p_10_25_t_s n3004 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17907 n3004 p_10_1_n2j c_10_25_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17906 vdd n3007 n3005 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17905 n3005 n3224 p_10_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17904 n3224 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17903 vdd n3437 n3225 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17902 n3222 p_10_1_n2j c_10_24_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17901 vdd p_10_24_t_s n3222 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17900 vdd a_22 n3226 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17899 n3227 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17898 n3439 p_10_2_d2j n3227 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17897 n3226 p_10_2_d2jbar n3439 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17896 n3437 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17895 n3225 n3439 p_10_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17894 n3217 c_10_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17893 c_10_24_s1_s c_10_24_b n3217 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17892 vdd c_10_24_s1_s n3434 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17891 c_10_24_s2_s c_9_25_cout n3431 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17890 n3214 c_10_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17889 n3430 c_10_24_b n3214 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17888 n3430 c_9_25_cout n3212 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17887 vdd c_10_24_a n3212 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17886 n3212 c_10_24_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17885 c_11_23_cin n3430 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17884 n3431 n3434 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17883 c_11_22_a c_10_24_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17882 c_11_21_a c_10_23_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17881 n3806 n3810 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17880 c_10_23_cout n3807 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17879 n4019 c_10_23_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17878 vdd c_10_23_b n4019 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17877 n3807 c_10_23_cin n4019 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17876 n3807 c_10_23_a n3805 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17875 n3805 c_10_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17874 c_10_23_s2_s c_10_23_cin n3806 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17873 vdd c_10_23_s1_s n3810 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17872 c_10_23_s1_s c_10_23_a n3803 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17871 n3803 c_10_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17870 n3816 p_10_2_d2j n3817 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17869 n3817 p_10_2_d2jbar n3818 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17868 n3818 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17867 vdd a_22 n3816 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17866 vdd p_10_23_t_s n3812 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17865 n3812 p_10_1_n2j c_10_23_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17864 vdd n3817 n3813 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17863 n3813 n3815 p_10_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17862 n3815 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17861 vdd n4236 n4026 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17860 n4025 p_10_1_n2j p_10_22_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17859 vdd p_10_22_t_s n4025 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17858 vdd a_20 n4027 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17857 n4028 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17856 n4239 p_10_2_d2j n4028 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17855 n4027 p_10_2_d2jbar n4239 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17854 n4236 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17853 n4026 n4239 p_10_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17852 n4023 c_10_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17851 c_10_22_s1_s p_10_22_pi2j n4023 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17850 vdd c_10_22_s1_s n4231 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17849 c_10_22_s2_s c_9_23_cout n4022 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17848 n4021 c_10_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17847 n4226 p_10_22_pi2j n4021 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17846 n4226 c_9_23_cout n4020 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17845 vdd c_10_22_a n4020 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17844 n4020 p_10_22_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17843 c_11_21_cin n4226 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17842 n4022 n4231 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17841 c_11_20_a c_10_22_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17840 c_11_19_a c_10_21_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17839 n4579 n4574 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17838 c_10_21_cout n4578 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17837 n4572 c_10_21_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17836 vdd p_10_21_pi2j n4572 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17835 n4578 c_10_21_cin n4572 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17834 n4578 c_10_21_a n4576 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17833 n4576 p_10_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17832 c_10_21_s2_s c_10_21_cin n4579 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17831 vdd c_10_21_s1_s n4574 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17830 c_10_21_s1_s c_10_21_a n4575 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17829 n4575 p_10_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17828 n4587 p_10_2_d2j n4588 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17827 n4588 p_10_2_d2jbar n4589 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17826 n4589 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17825 vdd a_20 n4587 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17824 vdd p_10_21_t_s n4583 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17823 n4583 p_10_1_n2j p_10_21_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17822 vdd n4588 n4584 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17821 n4584 n4586 p_10_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17820 n4586 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17819 vdd n4982 n4792 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17818 n4791 p_10_1_n2j p_10_20_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17817 vdd p_10_20_t_s n4791 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17816 vdd a_18 n4793 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17815 n4794 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17814 n4985 p_10_2_d2j n4794 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17813 n4793 p_10_2_d2jbar n4985 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17812 n4982 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17811 n4792 n4985 p_10_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17810 n4790 c_10_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17809 c_10_20_s1_s p_10_20_pi2j n4790 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17808 vdd c_10_20_s1_s n4978 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17807 c_10_20_s2_s c_9_21_cout n4789 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17806 n4788 c_10_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17805 n4974 p_10_20_pi2j n4788 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17804 n4974 c_9_21_cout n4787 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17803 vdd c_10_20_a n4787 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17802 n4787 p_10_20_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17801 c_11_19_cin n4974 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17800 n4789 n4978 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17799 c_11_18_a c_10_20_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17798 c_11_17_a c_10_19_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17797 n5333 n5328 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17796 c_10_19_cout n5332 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17795 n5324 c_10_19_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17794 vdd p_10_19_pi2j n5324 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17793 n5332 c_10_19_cin n5324 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17792 n5332 c_10_19_a n5330 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17791 n5330 p_10_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17790 c_10_19_s2_s c_10_19_cin n5333 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17789 vdd c_10_19_s1_s n5328 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17788 c_10_19_s1_s c_10_19_a n5329 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17787 n5329 p_10_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17786 n5341 p_10_2_d2j n5342 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17785 n5342 p_10_2_d2jbar n5343 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17784 n5343 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17783 vdd a_18 n5341 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17782 vdd p_10_19_t_s n5337 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17781 n5337 p_10_1_n2j p_10_19_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17780 vdd n5342 n5339 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17779 n5339 n5340 p_10_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17778 n5340 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17777 vdd n5735 n5551 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17776 n5550 p_10_1_n2j p_10_18_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17775 vdd p_10_18_t_s n5550 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17774 vdd a_16 n5552 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17773 n5553 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17772 n5737 p_10_2_d2j n5553 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17771 n5552 p_10_2_d2jbar n5737 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17770 n5735 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17769 n5551 n5737 p_10_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17768 n5326 c_10_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17767 c_10_18_s1_s p_10_18_pi2j n5326 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17766 vdd c_10_18_s1_s n5549 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17765 c_10_18_s2_s c_9_19_cout n5548 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17764 n5327 c_10_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17763 n5728 p_10_18_pi2j n5327 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17762 n5728 c_9_19_cout n5547 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17761 vdd c_10_18_a n5547 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17760 n5547 p_10_18_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17759 c_11_17_cin n5728 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17758 n5548 n5549 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17757 c_11_16_a c_10_18_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17756 c_11_15_a c_10_17_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17755 n6117 n6112 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17754 c_10_17_cout n6119 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17753 n6110 c_10_17_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17752 vdd p_10_17_pi2j n6110 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17751 n6119 c_10_17_cin n6110 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17750 n6119 c_10_17_a n6118 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17749 n6118 p_10_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17748 c_10_17_s2_s c_10_17_cin n6117 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17747 vdd c_10_17_s1_s n6112 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17746 c_10_17_s1_s c_10_17_a n6115 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17745 n6115 p_10_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17744 n5893 p_10_2_d2j n6121 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17743 n6121 p_10_2_d2jbar n5894 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17742 n5894 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17741 vdd a_16 n5893 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17740 vdd p_10_17_t_s n6124 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17739 n6124 p_10_1_n2j p_10_17_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17738 vdd n6121 n6128 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17737 n6128 n6126 p_10_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17736 n6126 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17735 vdd n6520 n6129 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17734 n6123 p_10_1_n2j p_10_16_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17733 vdd p_10_16_t_s n6123 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17732 vdd a_14 n6130 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17731 n6131 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17730 n6354 p_10_2_d2j n6131 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17729 n6130 p_10_2_d2jbar n6354 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17728 n6520 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17727 n6129 n6354 p_10_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17726 n6114 c_10_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17725 c_10_16_s1_s p_10_16_pi2j n6114 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17724 vdd c_10_16_s1_s n6351 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17723 c_10_16_s2_s c_9_17_cout n6349 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17722 n6113 c_10_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17721 n6513 p_10_16_pi2j n6113 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17720 n6513 c_9_17_cout n6348 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17719 vdd c_10_16_a n6348 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17718 n6348 p_10_16_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17717 c_11_15_cin n6513 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17716 n6349 n6351 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17715 c_11_14_a c_10_16_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17714 c_11_13_a c_10_15_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17713 n6701 n6702 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17712 c_10_15_cout n6921 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17711 n6915 c_10_15_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17710 vdd c_10_15_b n6915 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17709 n6921 c_10_15_cin n6915 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17708 n6921 c_10_15_a n6918 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17707 n6918 c_10_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17706 c_10_15_s2_s c_10_15_cin n6701 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17705 vdd c_10_15_s1_s n6702 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17704 c_10_15_s1_s c_10_15_a n6919 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17703 n6919 c_10_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17702 n6707 p_10_2_d2j n6708 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17701 n6708 p_10_2_d2jbar n6709 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17700 n6709 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17699 vdd a_14 n6707 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17698 vdd p_10_15_t_s n6705 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17697 n6705 p_10_1_n2j c_10_15_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17696 vdd n6708 n6706 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17695 n6706 n6926 p_10_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17694 n6926 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17693 vdd n7137 n6927 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17692 n6924 p_10_1_n2j p_10_14_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17691 vdd p_10_14_t_s n6924 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17690 vdd a_12 n6928 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17689 n6929 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17688 n7139 p_10_2_d2j n6929 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17687 n6928 p_10_2_d2jbar n7139 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17686 n7137 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17685 n6927 n7139 p_10_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17684 n6917 c_10_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17683 c_10_14_s1_s p_10_14_pi2j n6917 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17682 vdd c_10_14_s1_s n7134 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17681 c_10_14_s2_s c_9_15_cout n7132 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17680 n6916 c_10_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17679 n7131 p_10_14_pi2j n6916 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17678 n7131 c_9_15_cout n6914 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17677 vdd c_10_14_a n6914 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17676 n6914 p_10_14_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17675 c_11_13_cin n7131 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17674 n7132 n7134 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17673 c_11_12_a c_10_14_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17672 c_11_11_a c_10_13_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17671 n7486 n7491 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17670 c_10_13_cout n7487 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17669 n7700 c_10_13_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17668 vdd c_10_13_b n7700 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17667 n7487 c_10_13_cin n7700 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17666 n7487 c_10_13_a n7704 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17665 n7704 c_10_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17664 c_10_13_s2_s c_10_13_cin n7486 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17663 vdd c_10_13_s1_s n7491 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17662 c_10_13_s1_s c_10_13_a n7705 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17661 n7705 c_10_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17660 n7496 p_10_2_d2j n7497 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17659 n7497 p_10_2_d2jbar n7498 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17658 n7498 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17657 vdd a_12 n7496 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17656 vdd p_10_13_t_s n7493 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17655 n7493 p_10_1_n2j c_10_13_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17654 vdd n7497 n7494 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17653 n7494 n7495 p_10_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17652 n7495 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17651 vdd n7922 n7710 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17650 n7708 p_10_1_n2j c_10_12_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17649 vdd p_10_12_t_s n7708 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17648 vdd a_10 n7711 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17647 n7712 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17646 n7925 p_10_2_d2j n7712 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17645 n7711 p_10_2_d2jbar n7925 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17644 n7922 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17643 n7710 n7925 p_10_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17642 n7706 c_10_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17641 c_10_12_s1_s c_10_12_b n7706 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17640 vdd c_10_12_s1_s n7918 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17639 c_10_12_s2_s c_9_13_cout n7703 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17638 n7702 c_10_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17637 n7915 c_10_12_b n7702 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17636 n7915 c_9_13_cout n7701 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17635 vdd c_10_12_a n7701 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17634 n7701 c_10_12_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17633 c_11_11_cin n7915 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17632 n7703 n7918 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17631 c_11_10_a c_10_12_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17630 c_11_9_a c_10_11_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17629 n8266 n8262 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17628 c_10_11_cout n8267 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17627 n8260 c_10_11_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17626 vdd p_10_11_pi2j n8260 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17625 n8267 c_10_11_cin n8260 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17624 n8267 c_10_11_a n8265 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17623 n8265 p_10_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17622 c_10_11_s2_s c_10_11_cin n8266 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17621 vdd c_10_11_s1_s n8262 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17620 c_10_11_s1_s c_10_11_a n8263 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17619 n8263 p_10_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17618 n8275 p_10_2_d2j n8276 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17617 n8276 p_10_2_d2jbar n8277 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17616 n8277 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17615 vdd a_10 n8275 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17614 vdd p_10_11_t_s n8271 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17613 n8271 p_10_1_n2j p_10_11_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17612 vdd n8276 n8272 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17611 n8272 n8274 p_10_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17610 n8274 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17609 vdd n8671 n8481 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17608 n8480 p_10_1_n2j p_10_10_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17607 vdd p_10_10_t_s n8480 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17606 vdd a_8 n8482 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17605 n8483 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17604 n8673 p_10_2_d2j n8483 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17603 n8482 p_10_2_d2jbar n8673 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17602 n8671 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17601 n8481 n8673 p_10_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17600 n8479 c_10_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17599 c_10_10_s1_s p_10_10_pi2j n8479 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17598 vdd c_10_10_s1_s n8667 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17597 c_10_10_s2_s c_9_11_cout n8478 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17596 n8477 c_10_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17595 n8661 p_10_10_pi2j n8477 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17594 n8661 c_9_11_cout n8476 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17593 vdd c_10_10_a n8476 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17592 n8476 p_10_10_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17591 c_11_9_cin n8661 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17590 n8478 n8667 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17589 c_11_8_a c_10_10_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17588 c_11_7_a c_10_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17587 n9021 n9016 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17586 c_10_9_cout n9020 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17585 n9012 c_10_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17584 vdd p_10_9_pi2j n9012 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17583 n9020 c_10_9_cin n9012 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17582 n9020 c_10_9_a n9018 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17581 n9018 p_10_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17580 c_10_9_s2_s c_10_9_cin n9021 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17579 vdd c_10_9_s1_s n9016 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17578 c_10_9_s1_s c_10_9_a n9017 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17577 n9017 p_10_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17576 n9031 p_10_2_d2j n9030 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17575 n9030 p_10_2_d2jbar n9029 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17574 n9029 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17573 vdd a_8 n9031 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17572 vdd p_10_9_t_s n9025 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17571 n9025 p_10_1_n2j p_10_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17570 vdd n9030 n9027 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17569 n9027 n9028 p_10_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17568 n9028 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17567 vdd n9410 n9230 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17566 n9229 p_10_1_n2j p_10_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17565 vdd p_10_8_t_s n9229 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17564 vdd a_6 n9231 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17563 n9232 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17562 n9413 p_10_2_d2j n9232 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17561 n9231 p_10_2_d2jbar n9413 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17560 n9410 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17559 n9230 n9413 p_10_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17558 n9014 c_10_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17557 c_10_8_s1_s p_10_8_pi2j n9014 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17556 vdd c_10_8_s1_s n9405 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17555 c_10_8_s2_s c_9_9_cout n9228 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17554 n9015 c_10_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17553 n9402 p_10_8_pi2j n9015 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17552 n9402 c_9_9_cout n9227 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17551 vdd c_10_8_a n9227 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17550 n9227 p_10_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17549 c_11_7_cin n9402 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17548 n9228 n9405 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17547 c_11_6_a c_10_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17546 c_11_5_a c_10_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17545 n9802 n9798 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17544 c_10_7_cout n9803 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17543 n9794 c_10_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17542 vdd p_10_7_pi2j n9794 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17541 n9803 c_10_7_cin n9794 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17540 n9803 c_10_7_a n9801 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17539 n9801 p_10_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17538 c_10_7_s2_s c_10_7_cin n9802 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17537 vdd c_10_7_s1_s n9798 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17536 c_10_7_s1_s c_10_7_a n9799 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17535 n9799 p_10_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17534 n9571 p_10_2_d2j n9805 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17533 n9805 p_10_2_d2jbar n9572 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17532 n9572 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17531 vdd a_6 n9571 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17530 vdd p_10_7_t_s n9809 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17529 n9809 p_10_1_n2j p_10_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17528 vdd n9805 n9812 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17527 n9812 n9810 p_10_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17526 n9810 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17525 vdd n10189 n9813 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17524 n9807 p_10_1_n2j p_10_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17523 vdd p_10_6_t_s n9807 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17522 vdd a_4 n9814 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17521 n9815 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17520 n10188 p_10_2_d2j n9815 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17519 n9814 p_10_2_d2jbar n10188 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17518 n10189 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17517 n9813 n10188 p_10_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17516 n9797 c_10_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17515 c_10_6_s1_s p_10_6_pi2j n9797 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17514 vdd c_10_6_s1_s n10022 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17513 c_10_6_s2_s c_9_7_cout n10021 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17512 n9796 c_10_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17511 n10181 p_10_6_pi2j n9796 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17510 n10181 c_9_7_cout n10020 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17509 vdd c_10_6_a n10020 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17508 n10020 p_10_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17507 c_11_5_cin n10181 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17506 n10021 n10022 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17505 c_11_4_a c_10_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17504 c_11_3_a c_10_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17503 n10376 n10377 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17502 c_10_5_cout n10592 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17501 n10588 c_10_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17500 vdd c_10_5_b n10588 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17499 n10592 c_10_5_cin n10588 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17498 n10592 c_10_5_a n10593 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17497 n10593 c_10_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17496 c_10_5_s2_s c_10_5_cin n10376 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17495 vdd c_10_5_s1_s n10377 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17494 c_10_5_s1_s c_10_5_a n10590 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17493 n10590 c_10_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17492 n10382 p_10_2_d2j n10595 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17491 n10595 p_10_2_d2jbar n10383 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17490 n10383 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17489 vdd a_4 n10382 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17488 vdd p_10_5_t_s n10380 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17487 n10380 p_10_1_n2j c_10_5_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17486 vdd n10595 n10381 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17485 n10381 n10600 p_10_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17484 n10600 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17483 vdd n10811 n10601 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17482 n10598 p_10_1_n2j p_10_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17481 vdd p_10_4_t_s n10598 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17480 vdd a_2 n10602 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17479 n10603 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17478 n10814 p_10_2_d2j n10603 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17477 n10602 p_10_2_d2jbar n10814 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17476 n10811 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17475 n10601 n10814 p_10_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17474 n10591 c_10_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17473 c_10_4_s1_s p_10_4_pi2j n10591 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17472 vdd c_10_4_s1_s n10809 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17471 c_10_4_s2_s c_9_5_cout n10806 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17470 n10589 c_10_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17469 n10805 p_10_4_pi2j n10589 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17468 n10805 c_9_5_cout n10587 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17467 vdd c_10_4_a n10587 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17466 n10587 p_10_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17465 c_11_3_cin n10805 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17464 n10806 n10809 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17463 c_11_2_a c_10_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17462 c_11_1_a c_10_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17461 n11151 n11155 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17460 c_10_3_cout n11152 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17459 n11365 c_10_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17458 vdd c_10_3_b n11365 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17457 n11152 c_10_3_cin n11365 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17456 n11152 c_10_3_a n11371 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17455 n11371 c_10_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17454 c_10_3_s2_s c_10_3_cin n11151 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17453 vdd c_10_3_s1_s n11155 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17452 c_10_3_s1_s c_10_3_a n11369 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17451 n11369 c_10_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17450 n11161 p_10_2_d2j n11162 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17449 n11162 p_10_2_d2jbar n11163 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17448 n11163 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17447 vdd a_2 n11161 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17446 vdd p_10_3_t_s n11158 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17445 n11158 p_10_1_n2j c_10_3_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17444 vdd n11162 n11159 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17443 n11159 n11160 p_10_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17442 n11160 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17441 vdd n11585 n11375 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17440 n11373 p_10_1_n2j c_10_2_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17439 vdd p_10_2_t_s n11373 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17438 vdd a_0 n11376 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17437 n11377 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17436 n11587 p_10_2_d2j n11377 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17435 n11376 p_10_2_d2jbar n11587 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17434 n11585 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17433 n11375 n11587 p_10_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17432 n11370 c_10_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17431 c_10_2_s1_s c_10_2_b n11370 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17430 vdd c_10_2_s1_s n11581 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17429 c_10_2_s2_s c_9_3_cout n11368 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17428 n11367 c_10_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17427 n11578 c_10_2_b n11367 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17426 n11578 c_9_3_cout n11366 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17425 vdd c_10_2_a n11366 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17424 n11366 c_10_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17423 c_11_1_cin n11578 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17422 n11368 n11581 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17421 c_10_2_sum c_10_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17420 c_10_1_sum c_10_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17419 n11929 n11924 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17418 c_10_1_cout n11928 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17417 n11922 c_10_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17416 vdd p_10_1_pi2j n11922 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17415 n11928 c_10_1_cin n11922 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17414 n11928 c_10_1_a n11926 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17413 n11926 p_10_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17412 c_10_1_s2_s c_10_1_cin n11929 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17411 vdd c_10_1_s1_s n11924 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17410 c_10_1_s1_s c_10_1_a n11925 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17409 n11925 p_10_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17408 n11940 p_10_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17407 vdd a_0 n11940 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17406 vdd p_10_1_t_s n11934 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17405 n11934 p_10_1_n2j p_10_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17404 vdd n11940 n11936 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17403 n11936 n11938 p_10_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17402 n11938 p_10_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17401 n12124 c_9_1_sum cl4_10_s1_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17400 vdd n12305 n12124 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17399 p_14 cl4_10_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17398 n12296 c_9_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17397 vdd n12305 n12296 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17396 n12293 n12296 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17395 n12290 c_9_1_cout n12123 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17394 n12123 c_9_2_sum n12290 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17393 n12122 c_9_2_sum n12123 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_17392 vdd c_9_1_cout n12122 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_17391 n12123 c_9_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17390 vdd n12305 n12123 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17389 n12287 n12290 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17388 n12121 c_9_2_sum cl4_10_s2_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17387 vdd c_9_1_cout n12121 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17386 n12286 cl4_10_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_17385 n12120 n12293 cl4_10_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17384 vdd n12286 n12120 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17383 p_15 cl4_10_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17382 n167 p_9_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17381 c_9_33_s1_s c_9_31_a n167 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17380 vdd c_9_33_s1_s n163 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17379 c_9_33_s2_s c_9_32_cin n165 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17378 n161 p_9_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17377 n162 c_9_31_a n161 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17376 n162 c_9_32_cin n160 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17375 vdd p_9_33_pi2j n160 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17374 n160 c_9_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17373 c_10_32_cin n162 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17372 n165 n163 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17371 c_10_31_a c_9_33_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17370 n173 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17369 vdd p_9_33_t_s n169 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17368 n169 p_9_1_n2j p_9_33_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17367 vdd n173 n168 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17366 n168 n172 p_9_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17365 n172 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17364 vdd n513 n335 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17363 n334 p_9_1_n2j p_9_32_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17362 vdd p_9_32_t_s n334 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17361 vdd a_30 n336 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17360 n337 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17359 n515 p_9_2_d2j n337 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17358 n336 p_9_2_d2jbar n515 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17357 n513 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17356 n335 n515 p_9_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17355 n333 c_9_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17354 c_9_32_s1_s p_9_32_pi2j n333 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17353 vdd c_9_32_s1_s n510 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17352 c_9_32_s2_s c_9_32_cin n331 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17351 n332 c_9_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17350 n505 p_9_32_pi2j n332 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17349 n505 c_9_32_cin n330 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17348 vdd c_9_31_a n330 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17347 n330 p_9_32_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17346 c_10_31_cin n505 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17345 n331 n510 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17344 c_10_30_a c_9_32_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17343 c_10_29_a c_9_31_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17342 n849 n848 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17341 c_9_31_cout n852 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17340 n843 c_9_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17339 vdd p_9_31_pi2j n843 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17338 n852 c_9_31_cin n843 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17337 n852 c_9_31_a n850 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17336 n850 p_9_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17335 c_9_31_s2_s c_9_31_cin n849 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17334 vdd c_9_31_s1_s n848 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17333 c_9_31_s1_s c_9_31_a n846 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17332 n846 p_9_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17331 n859 p_9_2_d2j n857 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17330 n857 p_9_2_d2jbar n860 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17329 n860 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17328 vdd a_30 n859 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17327 vdd p_9_31_t_s n854 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17326 n854 p_9_1_n2j p_9_31_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17325 vdd n857 n853 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17324 n853 n858 p_9_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17323 n858 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17322 vdd n1268 n1057 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17321 n1056 p_9_1_n2j p_9_30_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17320 vdd p_9_30_t_s n1056 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17319 vdd a_28 n1058 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17318 n1059 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17317 n1270 p_9_2_d2j n1059 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17316 n1058 p_9_2_d2jbar n1270 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17315 n1268 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17314 n1057 n1270 p_9_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17313 n1055 c_9_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17312 c_9_30_s1_s p_9_30_pi2j n1055 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17311 vdd c_9_30_s1_s n1263 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17310 c_9_30_s2_s c_8_31_cout n1054 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17309 n1053 c_9_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17308 n1260 p_9_30_pi2j n1053 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17307 n1260 c_8_31_cout n1052 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17306 vdd c_9_30_a n1052 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17305 n1052 p_9_30_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17304 c_10_29_cin n1260 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17303 n1054 n1263 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17302 c_10_28_a c_9_30_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17301 c_10_27_a c_9_29_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17300 n1625 n1624 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17299 c_9_29_cout n1627 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17298 n1617 c_9_29_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17297 vdd p_9_29_pi2j n1617 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17296 n1627 c_9_29_cin n1617 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17295 n1627 c_9_29_a n1626 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17294 n1626 p_9_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17293 c_9_29_s2_s c_9_29_cin n1625 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17292 vdd c_9_29_s1_s n1624 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17291 c_9_29_s1_s c_9_29_a n1622 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17290 n1622 p_9_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17289 n1634 p_9_2_d2j n1633 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17288 n1633 p_9_2_d2jbar n1636 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17287 n1636 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17286 vdd a_28 n1634 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17285 vdd p_9_29_t_s n1629 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17284 n1629 p_9_1_n2j p_9_29_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17283 vdd n1633 n1630 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17282 n1630 n1635 p_9_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17281 n1635 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17280 vdd n2023 n1831 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17279 n1832 p_9_1_n2j p_9_28_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17278 vdd p_9_28_t_s n1832 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17277 vdd a_26 n1833 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17276 n1834 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17275 n2025 p_9_2_d2j n1834 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17274 n1833 p_9_2_d2jbar n2025 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17273 n2023 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17272 n1831 n2025 p_9_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17271 n1621 c_9_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17270 c_9_28_s1_s p_9_28_pi2j n1621 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17269 vdd c_9_28_s1_s n1830 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17268 c_9_28_s2_s c_8_29_cout n1829 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17267 n1620 c_9_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17266 n2015 p_9_28_pi2j n1620 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17265 n2015 c_8_29_cout n1828 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17264 vdd c_9_28_a n1828 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17263 n1828 p_9_28_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17262 c_10_27_cin n2015 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17261 n1829 n1830 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17260 c_10_26_a c_9_28_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17259 c_10_25_a c_9_27_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17258 n2191 n2431 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17257 c_9_27_cout n2438 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17256 n2430 c_9_27_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17255 vdd c_9_27_b n2430 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17254 n2438 c_9_27_cin n2430 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17253 n2438 c_9_27_a n2439 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17252 n2439 c_9_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17251 c_9_27_s2_s c_9_27_cin n2191 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17250 vdd c_9_27_s1_s n2431 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17249 c_9_27_s1_s c_9_27_a n2437 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17248 n2437 c_9_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17247 n2193 p_9_2_d2j n2441 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17246 n2441 p_9_2_d2jbar n2195 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17245 n2195 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17244 vdd a_26 n2193 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17243 vdd p_9_27_t_s n2192 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17242 n2192 p_9_1_n2j c_9_27_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17241 vdd n2441 n2444 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17240 n2444 n2445 p_9_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17239 n2445 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17238 vdd n2656 n2442 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17237 n2443 p_9_1_n2j p_9_26_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17236 vdd p_9_26_t_s n2443 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17235 vdd a_24 n2447 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17234 n2448 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17233 n2657 p_9_2_d2j n2448 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17232 n2447 p_9_2_d2jbar n2657 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17231 n2656 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17230 n2442 n2657 p_9_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17229 n2436 c_9_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17228 c_9_26_s1_s p_9_26_pi2j n2436 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17227 vdd c_9_26_s1_s n2655 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17226 c_9_26_s2_s c_8_27_cout n2654 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17225 n2435 c_9_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17224 n2832 p_9_26_pi2j n2435 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17223 n2832 c_8_27_cout n2652 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17222 vdd c_9_26_a n2652 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17221 n2652 p_9_26_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17220 c_10_25_cin n2832 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17219 n2654 n2655 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17218 c_10_24_a c_9_26_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17217 c_10_23_a c_9_25_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17216 n3011 n3012 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17215 c_9_25_cout n3236 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17214 n3229 c_9_25_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17213 vdd c_9_25_b n3229 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17212 n3236 c_9_25_cin n3229 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17211 n3236 c_9_25_a n3237 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17210 n3237 c_9_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17209 c_9_25_s2_s c_9_25_cin n3011 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17208 vdd c_9_25_s1_s n3012 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17207 c_9_25_s1_s c_9_25_a n3235 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17206 n3235 c_9_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17205 n3016 p_9_2_d2j n3015 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17204 n3015 p_9_2_d2jbar n3017 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17203 n3017 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17202 vdd a_24 n3016 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17201 vdd p_9_25_t_s n3014 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17200 n3014 p_9_1_n2j c_9_25_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17199 vdd n3015 n3013 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17198 n3013 n3240 p_9_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17197 n3240 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17196 vdd n3448 n3239 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17195 n3238 p_9_1_n2j c_9_24_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17194 vdd p_9_24_t_s n3238 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17193 vdd a_22 n3242 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17192 n3243 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17191 n3449 p_9_2_d2j n3243 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17190 n3242 p_9_2_d2jbar n3449 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17189 n3448 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17188 n3239 n3449 p_9_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17187 n3233 c_9_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17186 c_9_24_s1_s c_9_24_b n3233 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17185 vdd c_9_24_s1_s n3447 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17184 c_9_24_s2_s c_8_25_cout n3443 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17183 n3232 c_9_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17182 n3441 c_9_24_b n3232 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17181 n3441 c_8_25_cout n3228 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17180 vdd c_9_24_a n3228 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17179 n3228 c_9_24_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17178 c_10_23_cin n3441 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17177 n3443 n3447 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17176 c_10_22_a c_9_24_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17175 c_10_21_a c_9_23_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17174 n3824 n3827 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17173 c_9_23_cout n3825 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17172 n4030 c_9_23_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17171 vdd c_9_23_b n4030 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17170 n3825 c_9_23_cin n4030 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17169 n3825 c_9_23_a n3823 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17168 n3823 c_9_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17167 c_9_23_s2_s c_9_23_cin n3824 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17166 vdd c_9_23_s1_s n3827 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17165 c_9_23_s1_s c_9_23_a n3821 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17164 n3821 c_9_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17163 n3833 p_9_2_d2j n3831 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17162 n3831 p_9_2_d2jbar n3834 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17161 n3834 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17160 vdd a_22 n3833 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17159 vdd p_9_23_t_s n3829 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17158 n3829 p_9_1_n2j c_9_23_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17157 vdd n3831 n3828 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17156 n3828 n3832 p_9_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17155 n3832 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17154 vdd n4249 n4036 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17153 n4035 p_9_1_n2j p_9_22_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17152 vdd p_9_22_t_s n4035 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17151 vdd a_20 n4037 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17150 n4038 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17149 n4251 p_9_2_d2j n4038 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17148 n4037 p_9_2_d2jbar n4251 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17147 n4249 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17146 n4036 n4251 p_9_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17145 n4034 c_9_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17144 c_9_22_s1_s p_9_22_pi2j n4034 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17143 vdd c_9_22_s1_s n4247 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17142 c_9_22_s2_s c_8_23_cout n4032 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17141 n4033 c_9_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17140 n4241 p_9_22_pi2j n4033 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17139 n4241 c_8_23_cout n4029 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17138 vdd c_9_22_a n4029 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17137 n4029 p_9_22_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17136 c_10_21_cin n4241 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17135 n4032 n4247 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17134 c_10_20_a c_9_22_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17133 c_10_19_a c_9_21_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17132 n4598 n4593 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17131 c_9_21_cout n4596 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17130 n4590 c_9_21_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17129 vdd p_9_21_pi2j n4590 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17128 n4596 c_9_21_cin n4590 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17127 n4596 c_9_21_a n4599 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17126 n4599 p_9_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17125 c_9_21_s2_s c_9_21_cin n4598 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17124 vdd c_9_21_s1_s n4593 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17123 c_9_21_s1_s c_9_21_a n4594 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17122 n4594 p_9_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17121 n4606 p_9_2_d2j n4604 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17120 n4604 p_9_2_d2jbar n4607 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17119 n4607 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17118 vdd a_20 n4606 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17117 vdd p_9_21_t_s n4601 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17116 n4601 p_9_1_n2j p_9_21_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17115 vdd n4604 n4600 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17114 n4600 n4605 p_9_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17113 n4605 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17112 vdd n4995 n4800 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17111 n4799 p_9_1_n2j p_9_20_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17110 vdd p_9_20_t_s n4799 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17109 vdd a_18 n4801 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17108 n4802 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17107 n4997 p_9_2_d2j n4802 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17106 n4801 p_9_2_d2jbar n4997 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17105 n4995 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17104 n4800 n4997 p_9_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17103 n4798 c_9_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17102 c_9_20_s1_s p_9_20_pi2j n4798 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17101 vdd c_9_20_s1_s n4993 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17100 c_9_20_s2_s c_8_21_cout n4797 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17099 n4796 c_9_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17098 n4987 p_9_20_pi2j n4796 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17097 n4987 c_8_21_cout n4795 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17096 vdd c_9_20_a n4795 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17095 n4795 p_9_20_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17094 c_10_19_cin n4987 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17093 n4797 n4993 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17092 c_10_18_a c_9_20_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17091 c_10_17_a c_9_19_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17090 n5352 n5351 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17089 c_9_19_cout n5355 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17088 n5344 c_9_19_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17087 vdd p_9_19_pi2j n5344 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17086 n5355 c_9_19_cin n5344 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17085 n5355 c_9_19_a n5353 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17084 n5353 p_9_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17083 c_9_19_s2_s c_9_19_cin n5352 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17082 vdd c_9_19_s1_s n5351 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17081 c_9_19_s1_s c_9_19_a n5349 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17080 n5349 p_9_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17079 n5361 p_9_2_d2j n5360 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17078 n5360 p_9_2_d2jbar n5363 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17077 n5363 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17076 vdd a_18 n5361 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17075 vdd p_9_19_t_s n5356 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17074 n5356 p_9_1_n2j p_9_19_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17073 vdd n5360 n5357 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17072 n5357 n5362 p_9_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17071 n5362 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17070 vdd n5750 n5558 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17069 n5557 p_9_1_n2j p_9_18_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17068 vdd p_9_18_t_s n5557 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17067 vdd a_16 n5559 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17066 n5560 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17065 n5749 p_9_2_d2j n5560 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17064 n5559 p_9_2_d2jbar n5749 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17063 n5750 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17062 n5558 n5749 p_9_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17061 n5347 c_9_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17060 c_9_18_s1_s p_9_18_pi2j n5347 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17059 vdd c_9_18_s1_s n5556 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17058 c_9_18_s2_s c_8_19_cout n5555 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17057 n5348 c_9_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17056 n5740 p_9_18_pi2j n5348 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17055 n5740 c_8_19_cout n5554 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17054 vdd c_9_18_a n5554 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17053 n5554 p_9_18_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17052 c_10_17_cin n5740 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17051 n5555 n5556 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17050 c_10_16_a c_9_18_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17049 c_10_15_a c_9_17_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17048 n6141 n6133 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17047 c_9_17_cout n6143 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17046 n6132 c_9_17_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17045 vdd p_9_17_pi2j n6132 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17044 n6143 c_9_17_cin n6132 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17043 n6143 c_9_17_a n6142 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17042 n6142 p_9_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17041 c_9_17_s2_s c_9_17_cin n6141 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17040 vdd c_9_17_s1_s n6133 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17039 c_9_17_s1_s c_9_17_a n6138 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17038 n6138 p_9_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17037 n5898 p_9_2_d2j n6144 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17036 n6144 p_9_2_d2jbar n5900 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17035 n5900 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17034 vdd a_16 n5898 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17033 vdd p_9_17_t_s n6147 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17032 n6147 p_9_1_n2j p_9_17_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17031 vdd n6144 n6148 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17030 n6148 n6150 p_9_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17029 n6150 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17028 vdd n6533 n6145 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17027 n6146 p_9_1_n2j p_9_16_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17026 vdd p_9_16_t_s n6146 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17025 vdd a_14 n6152 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17024 n6153 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_17023 n6359 p_9_2_d2j n6153 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17022 n6152 p_9_2_d2jbar n6359 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_17021 n6533 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17020 n6145 n6359 p_9_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_17019 n6137 c_9_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17018 c_9_16_s1_s p_9_16_pi2j n6137 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17017 vdd c_9_16_s1_s n6358 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_17016 c_9_16_s2_s c_8_17_cout n6357 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_17015 n6136 c_9_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17014 n6526 p_9_16_pi2j n6136 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17013 n6526 c_8_17_cout n6355 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17012 vdd c_9_16_a n6355 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17011 n6355 p_9_16_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17010 c_10_15_cin n6526 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17009 n6357 n6358 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17008 c_10_14_a c_9_16_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17007 c_10_13_a c_9_15_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17006 n6712 n6713 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_17005 c_9_15_cout n6939 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_17004 n6931 c_9_15_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17003 vdd c_9_15_b n6931 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17002 n6939 c_9_15_cin n6931 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17001 n6939 c_9_15_a n6936 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_17000 n6936 c_9_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16999 c_9_15_s2_s c_9_15_cin n6712 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16998 vdd c_9_15_s1_s n6713 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16997 c_9_15_s1_s c_9_15_a n6937 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16996 n6937 c_9_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16995 n6717 p_9_2_d2j n6716 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16994 n6716 p_9_2_d2jbar n6718 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16993 n6718 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16992 vdd a_14 n6717 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16991 vdd p_9_15_t_s n6715 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16990 n6715 p_9_1_n2j c_9_15_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16989 vdd n6716 n6714 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16988 n6714 n6942 p_9_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16987 n6942 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16986 vdd n7147 n6941 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16985 n6940 p_9_1_n2j p_9_14_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16984 vdd p_9_14_t_s n6940 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16983 vdd a_12 n6944 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16982 n6945 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16981 n7148 p_9_2_d2j n6945 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16980 n6944 p_9_2_d2jbar n7148 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16979 n7147 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16978 n6941 n7148 p_9_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16977 n6935 c_9_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16976 c_9_14_s1_s p_9_14_pi2j n6935 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16975 vdd c_9_14_s1_s n7146 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16974 c_9_14_s2_s c_8_15_cout n7142 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16973 n6934 c_9_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16972 n7141 p_9_14_pi2j n6934 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16971 n7141 c_8_15_cout n6930 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16970 vdd c_9_14_a n6930 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16969 n6930 p_9_14_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16968 c_10_13_cin n7141 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16967 n7142 n7146 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16966 c_10_12_a c_9_14_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16965 c_10_11_a c_9_13_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16964 n7501 n7505 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16963 c_9_13_cout n7503 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16962 n7714 c_9_13_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16961 vdd c_9_13_b n7714 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16960 n7503 c_9_13_cin n7714 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16959 n7503 c_9_13_a n7719 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16958 n7719 c_9_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16957 c_9_13_s2_s c_9_13_cin n7501 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16956 vdd c_9_13_s1_s n7505 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16955 c_9_13_s1_s c_9_13_a n7720 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16954 n7720 c_9_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16953 n7510 p_9_2_d2j n7508 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16952 n7508 p_9_2_d2jbar n7511 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16951 n7511 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16950 vdd a_12 n7510 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16949 vdd p_9_13_t_s n7507 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16948 n7507 p_9_1_n2j c_9_13_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16947 vdd n7508 n7506 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16946 n7506 n7509 p_9_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16945 n7509 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16944 vdd n7934 n7722 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16943 n7721 p_9_1_n2j c_9_12_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16942 vdd p_9_12_t_s n7721 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16941 vdd a_10 n7724 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16940 n7725 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16939 n7936 p_9_2_d2j n7725 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16938 n7724 p_9_2_d2jbar n7936 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16937 n7934 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16936 n7722 n7936 p_9_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16935 n7718 c_9_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16934 c_9_12_s1_s c_9_12_b n7718 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16933 vdd c_9_12_s1_s n7933 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16932 c_9_12_s2_s c_8_13_cout n7716 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16931 n7717 c_9_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16930 n7928 c_9_12_b n7717 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16929 n7928 c_8_13_cout n7713 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16928 vdd c_9_12_a n7713 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16927 n7713 c_9_12_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16926 c_10_11_cin n7928 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16925 n7716 n7933 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16924 c_10_10_a c_9_12_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16923 c_10_9_a c_9_11_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16922 n8285 n8281 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16921 c_9_11_cout n8286 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16920 n8278 c_9_11_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16919 vdd p_9_11_pi2j n8278 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16918 n8286 c_9_11_cin n8278 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16917 n8286 c_9_11_a n8284 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16916 n8284 p_9_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16915 c_9_11_s2_s c_9_11_cin n8285 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16914 vdd c_9_11_s1_s n8281 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16913 c_9_11_s1_s c_9_11_a n8282 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16912 n8282 p_9_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16911 n8294 p_9_2_d2j n8292 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16910 n8292 p_9_2_d2jbar n8295 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16909 n8295 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16908 vdd a_10 n8294 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16907 vdd p_9_11_t_s n8289 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16906 n8289 p_9_1_n2j p_9_11_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16905 vdd n8292 n8288 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16904 n8288 n8293 p_9_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16903 n8293 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16902 vdd n8684 n8489 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16901 n8488 p_9_1_n2j p_9_10_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16900 vdd p_9_10_t_s n8488 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16899 vdd a_8 n8490 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16898 n8491 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16897 n8686 p_9_2_d2j n8491 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16896 n8490 p_9_2_d2jbar n8686 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16895 n8684 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16894 n8489 n8686 p_9_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16893 n8487 c_9_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16892 c_9_10_s1_s p_9_10_pi2j n8487 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16891 vdd c_9_10_s1_s n8680 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16890 c_9_10_s2_s c_8_11_cout n8486 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16889 n8485 c_9_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16888 n8676 p_9_10_pi2j n8485 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16887 n8676 c_8_11_cout n8484 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16886 vdd c_9_10_a n8484 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16885 n8484 p_9_10_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16884 c_10_9_cin n8676 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16883 n8486 n8680 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16882 c_10_8_a c_9_10_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16881 c_10_7_a c_9_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16880 n9040 n9039 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16879 c_9_9_cout n9043 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16878 n9032 c_9_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16877 vdd p_9_9_pi2j n9032 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16876 n9043 c_9_9_cin n9032 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16875 n9043 c_9_9_a n9041 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16874 n9041 p_9_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16873 c_9_9_s2_s c_9_9_cin n9040 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16872 vdd c_9_9_s1_s n9039 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16871 c_9_9_s1_s c_9_9_a n9037 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16870 n9037 p_9_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16869 n9049 p_9_2_d2j n9048 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16868 n9048 p_9_2_d2jbar n9051 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16867 n9051 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16866 vdd a_8 n9049 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16865 vdd p_9_9_t_s n9044 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16864 n9044 p_9_1_n2j p_9_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16863 vdd n9048 n9045 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16862 n9045 n9050 p_9_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16861 n9050 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16860 vdd n9426 n9236 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16859 n9235 p_9_1_n2j p_9_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16858 vdd p_9_8_t_s n9235 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16857 vdd a_6 n9237 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16856 n9238 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16855 n9425 p_9_2_d2j n9238 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16854 n9237 p_9_2_d2jbar n9425 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16853 n9426 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16852 n9236 n9425 p_9_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16851 n9035 c_9_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16850 c_9_8_s1_s p_9_8_pi2j n9035 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16849 vdd c_9_8_s1_s n9414 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16848 c_9_8_s2_s c_8_9_cout n9234 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16847 n9036 c_9_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16846 n9416 p_9_8_pi2j n9036 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16845 n9416 c_8_9_cout n9233 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16844 vdd c_9_8_a n9233 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16843 n9233 p_9_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16842 c_10_7_cin n9416 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16841 n9234 n9414 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16840 c_10_6_a c_9_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16839 c_10_5_a c_9_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16838 n9825 n9821 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16837 c_9_7_cout n9826 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16836 n9816 c_9_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16835 vdd p_9_7_pi2j n9816 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16834 n9826 c_9_7_cin n9816 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16833 n9826 c_9_7_a n9824 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16832 n9824 p_9_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16831 c_9_7_s2_s c_9_7_cin n9825 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16830 vdd c_9_7_s1_s n9821 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16829 c_9_7_s1_s c_9_7_a n9822 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16828 n9822 p_9_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16827 n9576 p_9_2_d2j n9828 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16826 n9828 p_9_2_d2jbar n9578 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16825 n9578 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16824 vdd a_6 n9576 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16823 vdd p_9_7_t_s n9831 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16822 n9831 p_9_1_n2j p_9_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16821 vdd n9828 n9832 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16820 n9832 n9834 p_9_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16819 n9834 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16818 vdd n10202 n9829 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16817 n9830 p_9_1_n2j p_9_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16816 vdd p_9_6_t_s n9830 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16815 vdd a_4 n9836 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16814 n9837 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16813 n10203 p_9_2_d2j n9837 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16812 n9836 p_9_2_d2jbar n10203 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16811 n10202 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16810 n9829 n10203 p_9_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16809 n9820 c_9_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16808 c_9_6_s1_s p_9_6_pi2j n9820 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16807 vdd c_9_6_s1_s n10027 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16806 c_9_6_s2_s c_8_7_cout n10026 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16805 n9819 c_9_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16804 n10195 p_9_6_pi2j n9819 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16803 n10195 c_8_7_cout n10025 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16802 vdd c_9_6_a n10025 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16801 n10025 p_9_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16800 c_10_5_cin n10195 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16799 n10026 n10027 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16798 c_10_4_a c_9_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16797 c_10_3_a c_9_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16796 n10386 n10388 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16795 c_9_5_cout n10611 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16794 n10605 c_9_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16793 vdd c_9_5_b n10605 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16792 n10611 c_9_5_cin n10605 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16791 n10611 c_9_5_a n10612 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16790 n10612 c_9_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16789 c_9_5_s2_s c_9_5_cin n10386 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16788 vdd c_9_5_s1_s n10388 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16787 c_9_5_s1_s c_9_5_a n10610 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16786 n10610 c_9_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16785 n10391 p_9_2_d2j n10614 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16784 n10614 p_9_2_d2jbar n10392 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16783 n10392 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16782 vdd a_4 n10391 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16781 vdd p_9_5_t_s n10390 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16780 n10390 p_9_1_n2j c_9_5_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16779 vdd n10614 n10389 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16778 n10389 n10617 p_9_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16777 n10617 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16776 vdd n10821 n10616 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16775 n10615 p_9_1_n2j p_9_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16774 vdd p_9_4_t_s n10615 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16773 vdd a_2 n10619 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16772 n10620 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16771 n10822 p_9_2_d2j n10620 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16770 n10619 p_9_2_d2jbar n10822 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16769 n10821 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16768 n10616 n10822 p_9_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16767 n10609 c_9_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16766 c_9_4_s1_s p_9_4_pi2j n10609 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16765 vdd c_9_4_s1_s n10820 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16764 c_9_4_s2_s c_8_5_cout n10817 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16763 n10608 c_9_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16762 n10815 p_9_4_pi2j n10608 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16761 n10815 c_8_5_cout n10604 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16760 vdd c_9_4_a n10604 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16759 n10604 p_9_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16758 c_10_3_cin n10815 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16757 n10817 n10820 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16756 c_10_2_a c_9_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16755 c_10_1_a c_9_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16754 n11166 n11170 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16753 c_9_3_cout n11168 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16752 n11379 c_9_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16751 vdd c_9_3_b n11379 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16750 n11168 c_9_3_cin n11379 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16749 n11168 c_9_3_a n11385 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16748 n11385 c_9_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16747 c_9_3_s2_s c_9_3_cin n11166 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16746 vdd c_9_3_s1_s n11170 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16745 c_9_3_s1_s c_9_3_a n11384 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16744 n11384 c_9_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16743 n11175 p_9_2_d2j n11173 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16742 n11173 p_9_2_d2jbar n11176 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16741 n11176 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16740 vdd a_2 n11175 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16739 vdd p_9_3_t_s n11172 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16738 n11172 p_9_1_n2j c_9_3_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16737 vdd n11173 n11171 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16736 n11171 n11174 p_9_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16735 n11174 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16734 vdd n11597 n11387 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16733 n11386 p_9_1_n2j c_9_2_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16732 vdd p_9_2_t_s n11386 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16731 vdd a_0 n11389 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16730 n11390 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16729 n11599 p_9_2_d2j n11390 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16728 n11389 p_9_2_d2jbar n11599 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16727 n11597 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16726 n11387 n11599 p_9_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16725 n11383 c_9_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16724 c_9_2_s1_s c_9_2_b n11383 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16723 vdd c_9_2_s1_s n11596 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16722 c_9_2_s2_s c_8_3_cout n11381 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16721 n11382 c_9_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16720 n11590 c_9_2_b n11382 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16719 n11590 c_8_3_cout n11378 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16718 vdd c_9_2_a n11378 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16717 n11378 c_9_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16716 c_10_1_cin n11590 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16715 n11381 n11596 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16714 c_9_2_sum c_9_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16713 c_9_1_sum c_9_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16712 n11949 n11944 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16711 c_9_1_cout n11947 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16710 n11941 c_9_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16709 vdd p_9_1_pi2j n11941 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16708 n11947 c_9_1_cin n11941 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16707 n11947 c_9_1_a n11950 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16706 n11950 p_9_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16705 c_9_1_s2_s c_9_1_cin n11949 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16704 vdd c_9_1_s1_s n11944 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16703 c_9_1_s1_s c_9_1_a n11945 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16702 n11945 p_9_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16701 n11958 p_9_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16700 vdd a_0 n11958 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16699 vdd p_9_1_t_s n11953 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16698 n11953 p_9_1_n2j p_9_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16697 vdd n11958 n11952 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16696 n11952 n11957 p_9_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16695 n11957 p_9_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16694 n12129 c_8_1_sum cl4_9_s1_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16693 vdd n12323 n12129 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16692 p_12 cl4_9_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16691 n12312 c_8_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16690 vdd n12323 n12312 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16689 n12311 n12312 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16688 n12309 c_8_1_cout n12128 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16687 n12128 c_8_2_sum n12309 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16686 n12127 c_8_2_sum n12128 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_16685 vdd c_8_1_cout n12127 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_16684 n12128 c_8_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16683 vdd n12323 n12128 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16682 n12305 n12309 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16681 n12126 c_8_2_sum cl4_9_s2_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16680 vdd c_8_1_cout n12126 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16679 n12304 cl4_9_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_16678 n12125 n12311 cl4_9_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16677 vdd n12304 n12125 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16676 p_13 cl4_9_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16675 n180 p_8_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16674 c_8_33_s1_s c_8_31_a n180 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16673 vdd c_8_33_s1_s n181 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16672 c_8_33_s2_s c_8_32_cin n179 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16671 n177 p_8_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16670 n178 c_8_31_a n177 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16669 n178 c_8_32_cin n174 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16668 vdd p_8_33_pi2j n174 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16667 n174 c_8_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16666 c_9_32_cin n178 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16665 n179 n181 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16664 c_9_31_a c_8_33_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16663 n187 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16662 vdd p_8_33_t_s n176 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16661 n176 p_8_1_n2j p_8_33_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16660 vdd n187 n185 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16659 n185 n186 p_8_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16658 n186 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16657 vdd n526 n343 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16656 n341 p_8_1_n2j p_8_32_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16655 vdd p_8_32_t_s n341 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16654 vdd a_30 n344 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16653 n345 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16652 n529 p_8_2_d2j n345 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16651 n344 p_8_2_d2jbar n529 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16650 n526 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16649 n343 n529 p_8_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16648 n342 c_8_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16647 c_8_32_s1_s p_8_32_pi2j n342 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16646 vdd c_8_32_s1_s n522 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16645 c_8_32_s2_s c_8_32_cin n340 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16644 n339 c_8_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16643 n517 p_8_32_pi2j n339 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16642 n517 c_8_32_cin n338 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16641 vdd c_8_31_a n338 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16640 n338 p_8_32_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16639 c_9_31_cin n517 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16638 n340 n522 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16637 c_9_30_a c_8_32_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16636 c_9_29_a c_8_31_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16635 n869 n868 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16634 c_8_31_cout n871 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16633 n862 c_8_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16632 vdd p_8_31_pi2j n862 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16631 n871 c_8_31_cin n862 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16630 n871 c_8_31_a n870 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16629 n870 p_8_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16628 c_8_31_s2_s c_8_31_cin n869 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16627 vdd c_8_31_s1_s n868 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16626 c_8_31_s1_s c_8_31_a n865 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16625 n865 p_8_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16624 n877 p_8_2_d2j n875 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16623 n875 p_8_2_d2jbar n876 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16622 n876 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16621 vdd a_30 n877 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16620 vdd p_8_31_t_s n866 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16619 n866 p_8_1_n2j p_8_31_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16618 vdd n875 n874 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16617 n874 n878 p_8_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16616 n878 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16615 vdd n1283 n1065 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16614 n1064 p_8_1_n2j p_8_30_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16613 vdd p_8_30_t_s n1064 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16612 vdd a_28 n1066 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16611 n1067 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16610 n1286 p_8_2_d2j n1067 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16609 n1066 p_8_2_d2jbar n1286 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16608 n1283 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16607 n1065 n1286 p_8_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16606 n1063 c_8_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16605 c_8_30_s1_s p_8_30_pi2j n1063 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16604 vdd c_8_30_s1_s n1280 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16603 c_8_30_s2_s c_6_31_cout n1061 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16602 n1062 c_8_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16601 n1275 p_8_30_pi2j n1062 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16600 n1275 c_6_31_cout n1060 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16599 vdd c_8_30_a n1060 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16598 n1060 p_8_30_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16597 c_9_29_cin n1275 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16596 n1061 n1280 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16595 c_9_28_a c_8_30_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16594 c_9_27_a c_8_29_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16593 n1648 n1644 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16592 c_8_29_cout n1649 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16591 n1638 c_8_29_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16590 vdd p_8_29_pi2j n1638 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16589 n1649 c_8_29_cin n1638 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16588 n1649 c_8_29_a n1647 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16587 n1647 p_8_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16586 c_8_29_s2_s c_8_29_cin n1648 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16585 vdd c_8_29_s1_s n1644 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16584 c_8_29_s1_s c_8_29_a n1645 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16583 n1645 p_8_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16582 n1655 p_8_2_d2j n1654 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16581 n1654 p_8_2_d2jbar n1653 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16580 n1653 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16579 vdd a_28 n1655 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16578 vdd p_8_29_t_s n1643 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16577 n1643 p_8_1_n2j p_8_29_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16576 vdd n1654 n1651 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16575 n1651 n1656 p_8_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16574 n1656 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16573 vdd n2040 n1839 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16572 n1837 p_8_1_n2j p_8_28_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16571 vdd p_8_28_t_s n1837 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16570 vdd a_26 n1841 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16569 n1840 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16568 n2039 p_8_2_d2j n1840 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16567 n1841 p_8_2_d2jbar n2039 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16566 n2040 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16565 n1839 n2039 p_8_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16564 n1642 c_8_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16563 c_8_28_s1_s p_8_28_pi2j n1642 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16562 vdd c_8_28_s1_s n1838 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16561 c_8_28_s2_s c_6_29_cout n1836 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16560 n1641 c_8_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16559 n2031 p_8_28_pi2j n1641 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16558 n2031 c_6_29_cout n1835 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16557 vdd c_8_28_a n1835 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16556 n1835 p_8_28_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16555 c_9_27_cin n2031 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16554 n1836 n1838 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16553 c_9_26_a c_8_28_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16552 c_9_25_a c_8_27_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16551 n2199 n2451 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16550 c_8_27_cout n2461 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16549 n2450 c_8_27_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16548 vdd c_8_27_b n2450 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16547 n2461 c_8_27_cin n2450 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16546 n2461 c_8_27_a n2460 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16545 n2460 c_8_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16544 c_8_27_s2_s c_8_27_cin n2199 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16543 vdd c_8_27_s1_s n2451 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16542 c_8_27_s1_s c_8_27_a n2459 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16541 n2459 c_8_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16540 n2201 p_8_2_d2j n2462 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16539 n2462 p_8_2_d2jbar n2200 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16538 n2200 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16537 vdd a_26 n2201 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16536 vdd p_8_27_t_s n2198 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16535 n2198 p_8_1_n2j c_8_27_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16534 vdd n2462 n2463 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16533 n2463 n2466 p_8_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16532 n2466 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16531 vdd n2664 n2464 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16530 n2456 p_8_1_n2j p_8_26_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16529 vdd p_8_26_t_s n2456 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16528 vdd a_24 n2467 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16527 n2468 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16526 n2667 p_8_2_d2j n2468 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16525 n2467 p_8_2_d2jbar n2667 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16524 n2664 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16523 n2464 n2667 p_8_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16522 n2457 c_8_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16521 c_8_26_s1_s p_8_26_pi2j n2457 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16520 vdd c_8_26_s1_s n2663 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16519 c_8_26_s2_s c_6_27_cout n2662 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16518 n2455 c_8_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16517 n2845 p_8_26_pi2j n2455 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16516 n2845 c_6_27_cout n2660 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16515 vdd c_8_26_a n2660 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16514 n2660 p_8_26_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16513 c_9_25_cin n2845 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16512 n2662 n2663 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16511 c_9_24_a c_8_26_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16510 c_9_23_a c_8_25_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16509 n3021 n3022 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16508 c_8_25_cout n3254 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16507 n3245 c_8_25_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16506 vdd c_8_25_b n3245 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16505 n3254 c_8_25_cin n3245 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16504 n3254 c_8_25_a n3253 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16503 n3253 c_8_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16502 c_8_25_s2_s c_8_25_cin n3021 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16501 vdd c_8_25_s1_s n3022 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16500 c_8_25_s1_s c_8_25_a n3252 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16499 n3252 c_8_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16498 n3026 p_8_2_d2j n3024 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16497 n3024 p_8_2_d2jbar n3025 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16496 n3025 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16495 vdd a_24 n3026 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16494 vdd p_8_25_t_s n3020 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16493 n3020 p_8_1_n2j c_8_25_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16492 vdd n3024 n3023 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16491 n3023 n3257 p_8_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16490 n3257 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16489 vdd n3459 n3256 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16488 n3249 p_8_1_n2j c_8_24_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16487 vdd p_8_24_t_s n3249 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16486 vdd a_22 n3258 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16485 n3259 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16484 n3462 p_8_2_d2j n3259 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16483 n3258 p_8_2_d2jbar n3462 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16482 n3459 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16481 n3256 n3462 p_8_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16480 n3250 c_8_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16479 c_8_24_s1_s c_8_24_b n3250 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16478 vdd c_8_24_s1_s n3456 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16477 c_8_24_s2_s c_6_25_cout n3455 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16476 n3248 c_8_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16475 n3452 c_8_24_b n3248 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16474 n3452 c_6_25_cout n3244 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16473 vdd c_8_24_a n3244 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16472 n3244 c_8_24_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16471 c_9_23_cin n3452 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16470 n3455 n3456 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16469 c_9_22_a c_8_24_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16468 c_9_21_a c_8_23_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16467 n3841 n3844 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16466 c_8_23_cout n3843 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16465 n4040 c_8_23_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16464 vdd c_8_23_b n4040 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16463 n3843 c_8_23_cin n4040 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16462 n3843 c_8_23_a n3840 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16461 n3840 c_8_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16460 c_8_23_s2_s c_8_23_cin n3841 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16459 vdd c_8_23_s1_s n3844 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16458 c_8_23_s1_s c_8_23_a n3839 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16457 n3839 c_8_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16456 n3849 p_8_2_d2j n3847 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16455 n3847 p_8_2_d2jbar n3848 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16454 n3848 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16453 vdd a_22 n3849 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16452 vdd p_8_23_t_s n3838 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16451 n3838 p_8_1_n2j c_8_23_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16450 vdd n3847 n3846 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16449 n3846 n3850 p_8_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16448 n3850 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16447 vdd n4264 n4046 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16446 n4044 p_8_1_n2j p_8_22_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16445 vdd p_8_22_t_s n4044 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16444 vdd a_20 n4047 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16443 n4048 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16442 n4267 p_8_2_d2j n4048 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16441 n4047 p_8_2_d2jbar n4267 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16440 n4264 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16439 n4046 n4267 p_8_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16438 n4045 c_8_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16437 c_8_22_s1_s p_8_22_pi2j n4045 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16436 vdd c_8_22_s1_s n4259 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16435 c_8_22_s2_s c_6_23_cout n4043 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16434 n4042 c_8_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16433 n4254 p_8_22_pi2j n4042 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16432 n4254 c_6_23_cout n4039 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16431 vdd c_8_22_a n4039 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16430 n4039 p_8_22_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16429 c_9_21_cin n4254 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16428 n4043 n4259 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16427 c_9_20_a c_8_22_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16426 c_9_19_a c_8_21_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16425 n4618 n4613 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16424 c_8_21_cout n4617 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16423 n4608 c_8_21_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16422 vdd p_8_21_pi2j n4608 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16421 n4617 c_8_21_cin n4608 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16420 n4617 c_8_21_a n4615 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16419 n4615 p_8_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16418 c_8_21_s2_s c_8_21_cin n4618 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16417 vdd c_8_21_s1_s n4613 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16416 c_8_21_s1_s c_8_21_a n4614 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16415 n4614 p_8_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16414 n4624 p_8_2_d2j n4622 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16413 n4622 p_8_2_d2jbar n4623 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16412 n4623 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16411 vdd a_20 n4624 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16410 vdd p_8_21_t_s n4612 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16409 n4612 p_8_1_n2j p_8_21_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16408 vdd n4622 n4621 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16407 n4621 n4625 p_8_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16406 n4625 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16405 vdd n5010 n4808 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16404 n4807 p_8_1_n2j p_8_20_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16403 vdd p_8_20_t_s n4807 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16402 vdd a_18 n4809 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16401 n4810 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16400 n5013 p_8_2_d2j n4810 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16399 n4809 p_8_2_d2jbar n5013 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16398 n5010 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16397 n4808 n5013 p_8_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16396 n4806 c_8_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16395 c_8_20_s1_s p_8_20_pi2j n4806 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16394 vdd c_8_20_s1_s n5006 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16393 c_8_20_s2_s c_6_21_cout n4804 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16392 n4805 c_8_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16391 n5002 p_8_20_pi2j n4805 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16390 n5002 c_6_21_cout n4803 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16389 vdd c_8_20_a n4803 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16388 n4803 p_8_20_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16387 c_9_19_cin n5002 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16386 n4804 n5006 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16385 c_9_18_a c_8_20_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16384 c_9_17_a c_8_19_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16383 n5375 n5371 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16382 c_8_19_cout n5376 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16381 n5364 c_8_19_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16380 vdd p_8_19_pi2j n5364 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16379 n5376 c_8_19_cin n5364 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16378 n5376 c_8_19_a n5374 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16377 n5374 p_8_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16376 c_8_19_s2_s c_8_19_cin n5375 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16375 vdd c_8_19_s1_s n5371 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16374 c_8_19_s1_s c_8_19_a n5372 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16373 n5372 p_8_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16372 n5382 p_8_2_d2j n5381 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16371 n5381 p_8_2_d2jbar n5380 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16370 n5380 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16369 vdd a_18 n5382 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16368 vdd p_8_19_t_s n5370 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16367 n5370 p_8_1_n2j p_8_19_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16366 vdd n5381 n5378 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16365 n5378 n5383 p_8_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16364 n5383 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16363 vdd n5764 n5565 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16362 n5563 p_8_1_n2j p_8_18_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16361 vdd p_8_18_t_s n5563 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16360 vdd a_16 n5566 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16359 n5567 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16358 n5766 p_8_2_d2j n5567 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16357 n5566 p_8_2_d2jbar n5766 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16356 n5764 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16355 n5565 n5766 p_8_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16354 n5369 c_8_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16353 c_8_18_s1_s p_8_18_pi2j n5369 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16352 vdd c_8_18_s1_s n5564 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16351 c_8_18_s2_s c_6_19_cout n5562 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16350 n5368 c_8_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16349 n5757 p_8_18_pi2j n5368 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16348 n5757 c_6_19_cout n5561 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16347 vdd c_8_18_a n5561 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16346 n5561 p_8_18_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16345 c_9_17_cin n5757 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16344 n5562 n5564 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16343 c_9_16_a c_8_18_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16342 c_9_15_a c_8_17_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16341 n6165 n6156 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16340 c_8_17_cout n6167 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16339 n6155 c_8_17_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16338 vdd p_8_17_pi2j n6155 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16337 n6167 c_8_17_cin n6155 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16336 n6167 c_8_17_a n6166 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16335 n6166 p_8_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16334 c_8_17_s2_s c_8_17_cin n6165 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16333 vdd c_8_17_s1_s n6156 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16332 c_8_17_s1_s c_8_17_a n6163 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16331 n6163 p_8_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16330 n5904 p_8_2_d2j n6168 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16329 n6168 p_8_2_d2jbar n5903 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16328 n5903 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16327 vdd a_16 n5904 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16326 vdd p_8_17_t_s n6161 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16325 n6161 p_8_1_n2j p_8_17_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16324 vdd n6168 n6169 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16323 n6169 n6173 p_8_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16322 n6173 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16321 vdd n6546 n6170 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16320 n6162 p_8_1_n2j p_8_16_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16319 vdd p_8_16_t_s n6162 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16318 vdd a_14 n6174 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16317 n6175 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16316 n6368 p_8_2_d2j n6175 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16315 n6174 p_8_2_d2jbar n6368 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16314 n6546 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16313 n6170 n6368 p_8_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16312 n6160 c_8_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16311 c_8_16_s1_s p_8_16_pi2j n6160 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16310 vdd c_8_16_s1_s n6365 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16309 c_8_16_s2_s c_6_17_cout n6364 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16308 n6159 c_8_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16307 n6540 p_8_16_pi2j n6159 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16306 n6540 c_6_17_cout n6362 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16305 vdd c_8_16_a n6362 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16304 n6362 p_8_16_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16303 c_9_15_cin n6540 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16302 n6364 n6365 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16301 c_9_14_a c_8_16_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16300 c_9_13_a c_8_15_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16299 n6722 n6723 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16298 c_8_15_cout n6955 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16297 n6947 c_8_15_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16296 vdd c_8_15_b n6947 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16295 n6955 c_8_15_cin n6947 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16294 n6955 c_8_15_a n6956 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16293 n6956 c_8_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16292 c_8_15_s2_s c_8_15_cin n6722 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16291 vdd c_8_15_s1_s n6723 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16290 c_8_15_s1_s c_8_15_a n6953 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16289 n6953 c_8_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16288 n6727 p_8_2_d2j n6725 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16287 n6725 p_8_2_d2jbar n6726 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16286 n6726 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16285 vdd a_14 n6727 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16284 vdd p_8_15_t_s n6721 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16283 n6721 p_8_1_n2j c_8_15_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16282 vdd n6725 n6724 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16281 n6724 n6959 p_8_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16280 n6959 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16279 vdd n7157 n6958 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16278 n6954 p_8_1_n2j p_8_14_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16277 vdd p_8_14_t_s n6954 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16276 vdd a_12 n6960 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16275 n6961 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16274 n7160 p_8_2_d2j n6961 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16273 n6960 p_8_2_d2jbar n7160 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16272 n7157 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16271 n6958 n7160 p_8_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16270 n6951 c_8_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16269 c_8_14_s1_s p_8_14_pi2j n6951 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16268 vdd c_8_14_s1_s n7154 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16267 c_8_14_s2_s c_6_15_cout n7153 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16266 n6950 c_8_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16265 n7151 p_8_14_pi2j n6950 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16264 n7151 c_6_15_cout n6946 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16263 vdd c_8_14_a n6946 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16262 n6946 p_8_14_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16261 c_9_13_cin n7151 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16260 n7153 n7154 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16259 c_9_12_a c_8_14_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16258 c_9_11_a c_8_13_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16257 n7516 n7519 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16256 c_8_13_cout n7517 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16255 n7727 c_8_13_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16254 vdd c_8_13_b n7727 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16253 n7517 c_8_13_cin n7727 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16252 n7517 c_8_13_a n7733 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16251 n7733 c_8_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16250 c_8_13_s2_s c_8_13_cin n7516 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16249 vdd c_8_13_s1_s n7519 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16248 c_8_13_s1_s c_8_13_a n7734 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16247 n7734 c_8_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16246 n7523 p_8_2_d2j n7521 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16245 n7521 p_8_2_d2jbar n7522 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16244 n7522 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16243 vdd a_12 n7523 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16242 vdd p_8_13_t_s n7515 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16241 n7515 p_8_1_n2j c_8_13_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16240 vdd n7521 n7520 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16239 n7520 n7524 p_8_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16238 n7524 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16237 vdd n7948 n7736 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16236 n7731 p_8_1_n2j c_8_12_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16235 vdd p_8_12_t_s n7731 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16234 vdd a_10 n7737 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16233 n7738 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16232 n7951 p_8_2_d2j n7738 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16231 n7737 p_8_2_d2jbar n7951 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16230 n7948 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16229 n7736 n7951 p_8_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16228 n7732 c_8_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16227 c_8_12_s1_s c_8_12_b n7732 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16226 vdd c_8_12_s1_s n7944 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16225 c_8_12_s2_s c_6_13_cout n7730 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16224 n7729 c_8_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16223 n7941 c_8_12_b n7729 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16222 n7941 c_6_13_cout n7726 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16221 vdd c_8_12_a n7726 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16220 n7726 c_8_12_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16219 c_9_11_cin n7941 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16218 n7730 n7944 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16217 c_9_10_a c_8_12_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16216 c_9_9_a c_8_11_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16215 n8305 n8301 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16214 c_8_11_cout n8306 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16213 n8297 c_8_11_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16212 vdd p_8_11_pi2j n8297 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16211 n8306 c_8_11_cin n8297 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16210 n8306 c_8_11_a n8304 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16209 n8304 p_8_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16208 c_8_11_s2_s c_8_11_cin n8305 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16207 vdd c_8_11_s1_s n8301 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16206 c_8_11_s1_s c_8_11_a n8302 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16205 n8302 p_8_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16204 n8312 p_8_2_d2j n8310 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16203 n8310 p_8_2_d2jbar n8311 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16202 n8311 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16201 vdd a_10 n8312 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16200 vdd p_8_11_t_s n8300 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16199 n8300 p_8_1_n2j p_8_11_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16198 vdd n8310 n8309 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16197 n8309 n8313 p_8_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16196 n8313 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16195 vdd n8699 n8497 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16194 n8496 p_8_1_n2j p_8_10_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16193 vdd p_8_10_t_s n8496 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16192 vdd a_8 n8498 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16191 n8499 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16190 n8702 p_8_2_d2j n8499 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16189 n8498 p_8_2_d2jbar n8702 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16188 n8699 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16187 n8497 n8702 p_8_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16186 n8495 c_8_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16185 c_8_10_s1_s p_8_10_pi2j n8495 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16184 vdd c_8_10_s1_s n8696 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16183 c_8_10_s2_s c_6_11_cout n8493 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16182 n8494 c_8_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16181 n8691 p_8_10_pi2j n8494 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16180 n8691 c_6_11_cout n8492 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16179 vdd c_8_10_a n8492 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16178 n8492 p_8_10_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16177 c_9_9_cin n8691 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16176 n8493 n8696 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16175 c_9_8_a c_8_10_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16174 c_9_7_a c_8_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16173 n9063 n9059 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16172 c_8_9_cout n9064 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16171 n9053 c_8_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16170 vdd p_8_9_pi2j n9053 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16169 n9064 c_8_9_cin n9053 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16168 n9064 c_8_9_a n9062 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16167 n9062 p_8_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16166 c_8_9_s2_s c_8_9_cin n9063 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16165 vdd c_8_9_s1_s n9059 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16164 c_8_9_s1_s c_8_9_a n9060 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16163 n9060 p_8_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16162 n9070 p_8_2_d2j n9069 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16161 n9069 p_8_2_d2jbar n9068 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16160 n9068 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16159 vdd a_8 n9070 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16158 vdd p_8_9_t_s n9058 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16157 n9058 p_8_1_n2j p_8_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16156 vdd n9069 n9066 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16155 n9066 n9071 p_8_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16154 n9071 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16153 vdd n9441 n9242 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16152 n9241 p_8_1_n2j p_8_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16151 vdd p_8_8_t_s n9241 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16150 vdd a_6 n9243 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16149 n9244 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16148 n9443 p_8_2_d2j n9244 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16147 n9243 p_8_2_d2jbar n9443 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16146 n9441 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16145 n9242 n9443 p_8_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16144 n9057 c_8_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16143 c_8_8_s1_s p_8_8_pi2j n9057 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16142 vdd c_8_8_s1_s n9429 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16141 c_8_8_s2_s c_6_9_cout n9240 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16140 n9056 c_8_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16139 n9432 p_8_8_pi2j n9056 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16138 n9432 c_6_9_cout n9239 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16137 vdd c_8_8_a n9239 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16136 n9239 p_8_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16135 c_9_7_cin n9432 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16134 n9240 n9429 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16133 c_9_6_a c_8_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16132 c_9_5_a c_8_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16131 n9849 n9846 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16130 c_8_7_cout n9851 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16129 n9839 c_8_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16128 vdd p_8_7_pi2j n9839 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16127 n9851 c_8_7_cin n9839 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16126 n9851 c_8_7_a n9848 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16125 n9848 p_8_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16124 c_8_7_s2_s c_8_7_cin n9849 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16123 vdd c_8_7_s1_s n9846 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16122 c_8_7_s1_s c_8_7_a n9847 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16121 n9847 p_8_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16120 n9582 p_8_2_d2j n9852 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16119 n9852 p_8_2_d2jbar n9581 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16118 n9581 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16117 vdd a_6 n9582 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16116 vdd p_8_7_t_s n9844 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16115 n9844 p_8_1_n2j p_8_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16114 vdd n9852 n9853 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16113 n9853 n9857 p_8_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16112 n9857 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16111 vdd n10217 n9854 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16110 n9845 p_8_1_n2j p_8_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16109 vdd p_8_6_t_s n9845 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16108 vdd a_4 n9858 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16107 n9859 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16106 n10215 p_8_2_d2j n9859 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16105 n9858 p_8_2_d2jbar n10215 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16104 n10217 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16103 n9854 n10215 p_8_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16102 n9843 c_8_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16101 c_8_6_s1_s p_8_6_pi2j n9843 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16100 vdd c_8_6_s1_s n10032 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16099 c_8_6_s2_s c_6_7_cout n10031 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16098 n9842 c_8_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16097 n10210 p_8_6_pi2j n9842 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16096 n10210 c_6_7_cout n10030 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16095 vdd c_8_6_a n10030 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16094 n10030 p_8_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16093 c_9_5_cin n10210 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16092 n10031 n10032 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16091 c_9_4_a c_8_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16090 c_9_3_a c_8_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16089 n10397 n10398 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16088 c_8_5_cout n10631 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16087 n10622 c_8_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16086 vdd c_8_5_b n10622 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16085 n10631 c_8_5_cin n10622 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16084 n10631 c_8_5_a n10630 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16083 n10630 c_8_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16082 c_8_5_s2_s c_8_5_cin n10397 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16081 vdd c_8_5_s1_s n10398 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16080 c_8_5_s1_s c_8_5_a n10629 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16079 n10629 c_8_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16078 n10401 p_8_2_d2j n10632 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16077 n10632 p_8_2_d2jbar n10400 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16076 n10400 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16075 vdd a_4 n10401 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16074 vdd p_8_5_t_s n10396 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16073 n10396 p_8_1_n2j c_8_5_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16072 vdd n10632 n10399 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16071 n10399 n10635 p_8_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16070 n10635 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16069 vdd n10831 n10634 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16068 n10626 p_8_1_n2j p_8_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16067 vdd p_8_4_t_s n10626 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16066 vdd a_2 n10636 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16065 n10637 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16064 n10834 p_8_2_d2j n10637 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16063 n10636 p_8_2_d2jbar n10834 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16062 n10831 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16061 n10634 n10834 p_8_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16060 n10627 c_8_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16059 c_8_4_s1_s p_8_4_pi2j n10627 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16058 vdd c_8_4_s1_s n10830 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16057 c_8_4_s2_s c_6_5_cout n10827 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16056 n10625 c_8_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16055 n10825 p_8_4_pi2j n10625 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16054 n10825 c_6_5_cout n10621 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16053 vdd c_8_4_a n10621 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16052 n10621 p_8_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16051 c_9_3_cin n10825 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16050 n10827 n10830 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16049 c_9_2_a c_8_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16048 c_9_1_a c_8_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16047 n11181 n11184 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16046 c_8_3_cout n11182 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16045 n11392 c_8_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16044 vdd c_8_3_b n11392 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16043 n11182 c_8_3_cin n11392 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16042 n11182 c_8_3_a n11398 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16041 n11398 c_8_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16040 c_8_3_s2_s c_8_3_cin n11181 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16039 vdd c_8_3_s1_s n11184 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16038 c_8_3_s1_s c_8_3_a n11399 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16037 n11399 c_8_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16036 n11188 p_8_2_d2j n11186 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16035 n11186 p_8_2_d2jbar n11187 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16034 n11187 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16033 vdd a_2 n11188 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16032 vdd p_8_3_t_s n11180 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16031 n11180 p_8_1_n2j c_8_3_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16030 vdd n11186 n11185 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16029 n11185 n11189 p_8_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16028 n11189 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16027 vdd n11611 n11401 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16026 n11396 p_8_1_n2j c_8_2_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16025 vdd p_8_2_t_s n11396 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16024 vdd a_0 n11402 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16023 n11403 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_16022 n11614 p_8_2_d2j n11403 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16021 n11402 p_8_2_d2jbar n11614 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_16020 n11611 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16019 n11401 n11614 p_8_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_16018 n11397 c_8_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16017 c_8_2_s1_s c_8_2_b n11397 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16016 vdd c_8_2_s1_s n11607 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_16015 c_8_2_s2_s c_6_3_cout n11395 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_16014 n11394 c_8_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16013 n11604 c_8_2_b n11394 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16012 n11604 c_6_3_cout n11391 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16011 vdd c_8_2_a n11391 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16010 n11391 c_8_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16009 c_9_1_cin n11604 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16008 n11395 n11607 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16007 c_8_2_sum c_8_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16006 c_8_1_sum c_8_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16005 n11969 n11967 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_16004 c_8_1_cout n11968 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_16003 n11961 c_8_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16002 vdd p_8_1_pi2j n11961 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16001 n11968 c_8_1_cin n11961 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_16000 n11968 c_8_1_a n11970 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15999 n11970 p_8_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15998 c_8_1_s2_s c_8_1_cin n11969 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15997 vdd c_8_1_s1_s n11967 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15996 c_8_1_s1_s c_8_1_a n11964 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15995 n11964 p_8_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15994 n11978 p_8_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15993 vdd a_0 n11978 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15992 vdd p_8_1_t_s n11965 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15991 n11965 p_8_1_n2j p_8_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15990 vdd n11978 n11973 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15989 n11973 n11977 p_8_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15988 n11977 p_8_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15987 n12134 c_6_1_sum cl4_8_s1_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15986 vdd n12339 n12134 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15985 p_10 cl4_8_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15984 n12329 c_6_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15983 vdd n12339 n12329 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15982 n12328 n12329 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15981 n12324 c_6_1_cout n12132 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15980 n12132 c_6_2_sum n12324 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15979 n12133 c_6_2_sum n12132 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_15978 vdd c_6_1_cout n12133 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_15977 n12132 c_6_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15976 vdd n12339 n12132 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15975 n12323 n12324 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15974 n12131 c_6_2_sum cl4_8_s2_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15973 vdd c_6_1_cout n12131 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15972 n12320 cl4_8_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_15971 n12130 n12328 cl4_8_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15970 vdd n12320 n12130 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15969 p_11 cl4_8_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15968 n194 p_6_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15967 c_6_33_s1_s c_6_31_a n194 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15966 vdd c_6_33_s1_s n191 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15965 c_6_33_s2_s c_6_32_cin n192 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15964 n189 p_6_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15963 n190 c_6_31_a n189 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15962 n190 c_6_32_cin n188 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15961 vdd p_6_33_pi2j n188 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15960 n188 c_6_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15959 c_8_32_cin n190 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15958 n192 n191 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15957 c_8_31_a c_6_33_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15956 n201 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15955 vdd p_6_33_t_s n197 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15954 n197 p_6_1_n2j p_6_33_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15953 vdd n201 n200 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15952 n200 n198 p_6_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15951 n198 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15950 vdd n538 n351 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15949 n350 p_6_1_n2j p_6_32_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15948 vdd p_6_32_t_s n350 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15947 vdd a_30 n352 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15946 n353 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15945 n541 p_6_2_d2j n353 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15944 n352 p_6_2_d2jbar n541 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15943 n538 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15942 n351 n541 p_6_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15941 n349 c_6_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15940 c_6_32_s1_s p_6_32_pi2j n349 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15939 vdd c_6_32_s1_s n535 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15938 c_6_32_s2_s c_6_32_cin n348 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15937 n347 c_6_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15936 n530 p_6_32_pi2j n347 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15935 n530 c_6_32_cin n346 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15934 vdd c_6_31_a n346 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15933 n346 p_6_32_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15932 c_8_31_cin n530 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15931 n348 n535 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15930 c_8_30_a c_6_32_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15929 c_8_29_a c_6_31_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15928 n884 n883 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15927 c_6_31_cout n887 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15926 n879 c_6_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15925 vdd p_6_31_pi2j n879 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15924 n887 c_6_31_cin n879 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15923 n887 c_6_31_a n885 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15922 n885 p_6_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15921 c_6_31_s2_s c_6_31_cin n884 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15920 vdd c_6_31_s1_s n883 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15919 c_6_31_s1_s c_6_31_a n881 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15918 n881 p_6_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15917 n894 p_6_2_d2j n895 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15916 n895 p_6_2_d2jbar n896 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15915 n896 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15914 vdd a_30 n894 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15913 vdd p_6_31_t_s n890 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15912 n890 p_6_1_n2j p_6_31_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15911 vdd n895 n891 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15910 n891 n893 p_6_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15909 n893 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15908 vdd n1298 n1073 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15907 n1072 p_6_1_n2j p_6_30_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15906 vdd p_6_30_t_s n1072 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15905 vdd a_28 n1074 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15904 n1075 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15903 n1301 p_6_2_d2j n1075 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15902 n1074 p_6_2_d2jbar n1301 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15901 n1298 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15900 n1073 n1301 p_6_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15899 n1071 c_6_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15898 c_6_30_s1_s p_6_30_pi2j n1071 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15897 vdd c_6_30_s1_s n1293 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15896 c_6_30_s2_s c_5_31_cout n1070 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15895 n1069 c_6_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15894 n1288 p_6_30_pi2j n1069 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15893 n1288 c_5_31_cout n1068 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15892 vdd c_6_30_a n1068 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15891 n1068 p_6_30_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15890 c_8_29_cin n1288 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15889 n1070 n1293 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15888 c_8_28_a c_6_30_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15887 c_8_27_a c_6_29_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15886 n1665 n1661 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15885 c_6_29_cout n1666 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15884 n1657 c_6_29_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15883 vdd p_6_29_pi2j n1657 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15882 n1666 c_6_29_cin n1657 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15881 n1666 c_6_29_a n1664 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15880 n1664 p_6_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15879 c_6_29_s2_s c_6_29_cin n1665 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15878 vdd c_6_29_s1_s n1661 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15877 c_6_29_s1_s c_6_29_a n1662 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15876 n1662 p_6_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15875 n1674 p_6_2_d2j n1675 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15874 n1675 p_6_2_d2jbar n1676 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15873 n1676 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15872 vdd a_28 n1674 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15871 vdd p_6_29_t_s n1669 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15870 n1669 p_6_1_n2j p_6_29_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15869 vdd n1675 n1672 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15868 n1672 n1673 p_6_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15867 n1673 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15866 vdd n2051 n1846 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15865 n1845 p_6_1_n2j p_6_28_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15864 vdd p_6_28_t_s n1845 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15863 vdd a_26 n1848 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15862 n1847 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15861 n2054 p_6_2_d2j n1847 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15860 n1848 p_6_2_d2jbar n2054 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15859 n2051 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15858 n1846 n2054 p_6_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15857 n1660 c_6_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15856 c_6_28_s1_s p_6_28_pi2j n1660 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15855 vdd c_6_28_s1_s n1844 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15854 c_6_28_s2_s c_5_29_cout n1843 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15853 n1659 c_6_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15852 n2044 p_6_28_pi2j n1659 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15851 n2044 c_5_29_cout n1842 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15850 vdd c_6_28_a n1842 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15849 n1842 p_6_28_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15848 c_8_27_cin n2044 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15847 n1843 n1844 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15846 c_8_26_a c_6_28_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15845 c_8_25_a c_6_27_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15844 n2205 n2470 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15843 c_6_27_cout n2478 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15842 n2469 c_6_27_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15841 vdd c_6_27_b n2469 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15840 n2478 c_6_27_cin n2469 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15839 n2478 c_6_27_a n2475 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15838 n2475 c_6_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15837 c_6_27_s2_s c_6_27_cin n2205 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15836 vdd c_6_27_s1_s n2470 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15835 c_6_27_s1_s c_6_27_a n2477 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15834 n2477 c_6_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15833 n2207 p_6_2_d2j n2479 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15832 n2479 p_6_2_d2jbar n2208 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15831 n2208 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15830 vdd a_26 n2207 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15829 vdd p_6_27_t_s n2206 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15828 n2206 p_6_1_n2j c_6_27_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15827 vdd n2479 n2485 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15826 n2485 n2483 p_6_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15825 n2483 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15824 vdd n2672 n2486 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15823 n2482 p_6_1_n2j p_6_26_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15822 vdd p_6_26_t_s n2482 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15821 vdd a_24 n2488 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15820 n2487 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15819 n2675 p_6_2_d2j n2487 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15818 n2488 p_6_2_d2jbar n2675 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15817 n2672 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15816 n2486 n2675 p_6_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15815 n2474 c_6_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15814 c_6_26_s1_s p_6_26_pi2j n2474 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15813 vdd c_6_26_s1_s n2671 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15812 c_6_26_s2_s c_5_27_cout n2669 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15811 n2473 c_6_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15810 n2857 p_6_26_pi2j n2473 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15809 n2857 c_5_27_cout n2668 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15808 vdd c_6_26_a n2668 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15807 n2668 p_6_26_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15806 c_8_25_cin n2857 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15805 n2669 n2671 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15804 c_8_24_a c_6_26_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15803 c_8_23_a c_6_25_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15802 n3027 n3028 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15801 c_6_25_cout n3266 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15800 n3260 c_6_25_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15799 vdd c_6_25_b n3260 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15798 n3266 c_6_25_cin n3260 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15797 n3266 c_6_25_a n3267 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15796 n3267 c_6_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15795 c_6_25_s2_s c_6_25_cin n3027 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15794 vdd c_6_25_s1_s n3028 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15793 c_6_25_s1_s c_6_25_a n3264 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15792 n3264 c_6_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15791 n3033 p_6_2_d2j n3034 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15790 n3034 p_6_2_d2jbar n3035 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15789 n3035 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15788 vdd a_24 n3033 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15787 vdd p_6_25_t_s n3031 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15786 n3031 p_6_1_n2j c_6_25_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15785 vdd n3034 n3032 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15784 n3032 n3272 p_6_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15783 n3272 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15782 vdd n3470 n3273 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15781 n3270 p_6_1_n2j c_6_24_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15780 vdd p_6_24_t_s n3270 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15779 vdd a_22 n3274 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15778 n3275 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15777 n3471 p_6_2_d2j n3275 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15776 n3274 p_6_2_d2jbar n3471 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15775 n3470 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15774 n3273 n3471 p_6_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15773 n3265 c_6_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15772 c_6_24_s1_s c_6_24_b n3265 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15771 vdd c_6_24_s1_s n3467 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15770 c_6_24_s2_s c_5_25_cout n3464 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15769 n3262 c_6_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15768 n3463 c_6_24_b n3262 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15767 n3463 c_5_25_cout n3261 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15766 vdd c_6_24_a n3261 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15765 n3261 c_6_24_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15764 c_8_23_cin n3463 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15763 n3464 n3467 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15762 c_8_22_a c_6_24_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15761 c_8_21_a c_6_23_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15760 n3854 n3858 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15759 c_6_23_cout n3855 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15758 n4049 c_6_23_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15757 vdd c_6_23_b n4049 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15756 n3855 c_6_23_cin n4049 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15755 n3855 c_6_23_a n3853 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15754 n3853 c_6_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15753 c_6_23_s2_s c_6_23_cin n3854 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15752 vdd c_6_23_s1_s n3858 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15751 c_6_23_s1_s c_6_23_a n3851 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15750 n3851 c_6_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15749 n3864 p_6_2_d2j n3865 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15748 n3865 p_6_2_d2jbar n3866 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15747 n3866 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15746 vdd a_22 n3864 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15745 vdd p_6_23_t_s n3860 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15744 n3860 p_6_1_n2j c_6_23_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15743 vdd n3865 n3861 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15742 n3861 n3863 p_6_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15741 n3863 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15740 vdd n4278 n4056 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15739 n4055 p_6_1_n2j p_6_22_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15738 vdd p_6_22_t_s n4055 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15737 vdd a_20 n4057 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15736 n4058 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15735 n4280 p_6_2_d2j n4058 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15734 n4057 p_6_2_d2jbar n4280 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15733 n4278 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15732 n4056 n4280 p_6_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15731 n4053 c_6_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15730 c_6_22_s1_s p_6_22_pi2j n4053 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15729 vdd c_6_22_s1_s n4273 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15728 c_6_22_s2_s c_5_23_cout n4052 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15727 n4051 c_6_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15726 n4268 p_6_22_pi2j n4051 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15725 n4268 c_5_23_cout n4050 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15724 vdd c_6_22_a n4050 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15723 n4050 p_6_22_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15722 c_8_21_cin n4268 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15721 n4052 n4273 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15720 c_8_20_a c_6_22_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15719 c_8_19_a c_6_21_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15718 n4633 n4628 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15717 c_6_21_cout n4632 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15716 n4626 c_6_21_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15715 vdd p_6_21_pi2j n4626 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15714 n4632 c_6_21_cin n4626 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15713 n4632 c_6_21_a n4630 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15712 n4630 p_6_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15711 c_6_21_s2_s c_6_21_cin n4633 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15710 vdd c_6_21_s1_s n4628 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15709 c_6_21_s1_s c_6_21_a n4629 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15708 n4629 p_6_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15707 n4641 p_6_2_d2j n4642 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15706 n4642 p_6_2_d2jbar n4643 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15705 n4643 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15704 vdd a_20 n4641 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15703 vdd p_6_21_t_s n4637 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15702 n4637 p_6_1_n2j p_6_21_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15701 vdd n4642 n4638 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15700 n4638 n4640 p_6_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15699 n4640 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15698 vdd n5024 n4816 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15697 n4815 p_6_1_n2j p_6_20_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15696 vdd p_6_20_t_s n4815 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15695 vdd a_18 n4817 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15694 n4818 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15693 n5027 p_6_2_d2j n4818 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15692 n4817 p_6_2_d2jbar n5027 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15691 n5024 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15690 n4816 n5027 p_6_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15689 n4814 c_6_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15688 c_6_20_s1_s p_6_20_pi2j n4814 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15687 vdd c_6_20_s1_s n5019 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15686 c_6_20_s2_s c_5_21_cout n4813 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15685 n4812 c_6_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15684 n5016 p_6_20_pi2j n4812 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15683 n5016 c_5_21_cout n4811 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15682 vdd c_6_20_a n4811 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15681 n4811 p_6_20_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15680 c_8_19_cin n5016 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15679 n4813 n5019 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15678 c_8_18_a c_6_20_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15677 c_8_17_a c_6_19_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15676 n5393 n5388 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15675 c_6_19_cout n5392 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15674 n5384 c_6_19_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15673 vdd p_6_19_pi2j n5384 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15672 n5392 c_6_19_cin n5384 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15671 n5392 c_6_19_a n5390 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15670 n5390 p_6_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15669 c_6_19_s2_s c_6_19_cin n5393 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15668 vdd c_6_19_s1_s n5388 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15667 c_6_19_s1_s c_6_19_a n5389 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15666 n5389 p_6_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15665 n5401 p_6_2_d2j n5402 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15664 n5402 p_6_2_d2jbar n5403 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15663 n5403 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15662 vdd a_18 n5401 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15661 vdd p_6_19_t_s n5396 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15660 n5396 p_6_1_n2j p_6_19_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15659 vdd n5402 n5399 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15658 n5399 n5400 p_6_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15657 n5400 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15656 vdd n5777 n5572 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15655 n5571 p_6_1_n2j p_6_18_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15654 vdd p_6_18_t_s n5571 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15653 vdd a_16 n5573 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15652 n5574 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15651 n5780 p_6_2_d2j n5574 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15650 n5573 p_6_2_d2jbar n5780 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15649 n5777 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15648 n5572 n5780 p_6_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15647 n5386 c_6_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15646 c_6_18_s1_s p_6_18_pi2j n5386 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15645 vdd c_6_18_s1_s n5570 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15644 c_6_18_s2_s c_5_19_cout n5569 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15643 n5387 c_6_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15642 n5769 p_6_18_pi2j n5387 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15641 n5769 c_5_19_cout n5568 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15640 vdd c_6_18_a n5568 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15639 n5568 p_6_18_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15638 c_8_17_cin n5769 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15637 n5569 n5570 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15636 c_8_16_a c_6_18_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15635 c_8_15_a c_6_17_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15634 n6183 n6178 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15633 c_6_17_cout n6185 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15632 n6176 c_6_17_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15631 vdd p_6_17_pi2j n6176 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15630 n6185 c_6_17_cin n6176 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15629 n6185 c_6_17_a n6184 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15628 n6184 p_6_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15627 c_6_17_s2_s c_6_17_cin n6183 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15626 vdd c_6_17_s1_s n6178 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15625 c_6_17_s1_s c_6_17_a n6181 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15624 n6181 p_6_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15623 n5908 p_6_2_d2j n6187 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15622 n6187 p_6_2_d2jbar n5909 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15621 n5909 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15620 vdd a_16 n5908 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15619 vdd p_6_17_t_s n6190 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15618 n6190 p_6_1_n2j p_6_17_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15617 vdd n6187 n6194 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15616 n6194 n6192 p_6_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15615 n6192 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15614 vdd n6559 n6195 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15613 n6189 p_6_1_n2j p_6_16_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15612 vdd p_6_16_t_s n6189 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15611 vdd a_14 n6196 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15610 n6197 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15609 n6374 p_6_2_d2j n6197 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15608 n6196 p_6_2_d2jbar n6374 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15607 n6559 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15606 n6195 n6374 p_6_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15605 n6180 c_6_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15604 c_6_16_s1_s p_6_16_pi2j n6180 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15603 vdd c_6_16_s1_s n6372 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15602 c_6_16_s2_s c_5_17_cout n6370 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15601 n6179 c_6_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15600 n6552 p_6_16_pi2j n6179 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15599 n6552 c_5_17_cout n6369 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15598 vdd c_6_16_a n6369 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15597 n6369 p_6_16_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15596 c_8_15_cin n6552 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15595 n6370 n6372 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15594 c_8_14_a c_6_16_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15593 c_8_13_a c_6_15_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15592 n6728 n6729 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15591 c_6_15_cout n6969 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15590 n6963 c_6_15_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15589 vdd c_6_15_b n6963 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15588 n6969 c_6_15_cin n6963 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15587 n6969 c_6_15_a n6966 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15586 n6966 c_6_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15585 c_6_15_s2_s c_6_15_cin n6728 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15584 vdd c_6_15_s1_s n6729 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15583 c_6_15_s1_s c_6_15_a n6967 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15582 n6967 c_6_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15581 n6734 p_6_2_d2j n6735 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15580 n6735 p_6_2_d2jbar n6736 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15579 n6736 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15578 vdd a_14 n6734 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15577 vdd p_6_15_t_s n6732 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15576 n6732 p_6_1_n2j c_6_15_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15575 vdd n6735 n6733 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15574 n6733 n6974 p_6_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15573 n6974 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15572 vdd n7167 n6975 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15571 n6972 p_6_1_n2j p_6_14_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15570 vdd p_6_14_t_s n6972 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15569 vdd a_12 n6976 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15568 n6977 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15567 n7168 p_6_2_d2j n6977 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15566 n6976 p_6_2_d2jbar n7168 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15565 n7167 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15564 n6975 n7168 p_6_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15563 n6965 c_6_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15562 c_6_14_s1_s p_6_14_pi2j n6965 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15561 vdd c_6_14_s1_s n7164 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15560 c_6_14_s2_s c_5_15_cout n7162 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15559 n6964 c_6_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15558 n7161 p_6_14_pi2j n6964 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15557 n7161 c_5_15_cout n6962 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15556 vdd c_6_14_a n6962 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15555 n6962 p_6_14_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15554 c_8_13_cin n7161 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15553 n7162 n7164 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15552 c_8_12_a c_6_14_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15551 c_8_11_a c_6_13_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15550 n7525 n7529 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15549 c_6_13_cout n7526 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15548 n7739 c_6_13_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15547 vdd c_6_13_b n7739 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15546 n7526 c_6_13_cin n7739 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15545 n7526 c_6_13_a n7743 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15544 n7743 c_6_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15543 c_6_13_s2_s c_6_13_cin n7525 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15542 vdd c_6_13_s1_s n7529 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15541 c_6_13_s1_s c_6_13_a n7744 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15540 n7744 c_6_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15539 n7535 p_6_2_d2j n7536 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15538 n7536 p_6_2_d2jbar n7537 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15537 n7537 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15536 vdd a_12 n7535 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15535 vdd p_6_13_t_s n7531 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15534 n7531 p_6_1_n2j c_6_13_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15533 vdd n7536 n7533 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15532 n7533 n7534 p_6_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15531 n7534 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15530 vdd n7961 n7749 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15529 n7747 p_6_1_n2j c_6_12_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15528 vdd p_6_12_t_s n7747 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15527 vdd a_10 n7750 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15526 n7751 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15525 n7964 p_6_2_d2j n7751 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15524 n7750 p_6_2_d2jbar n7964 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15523 n7961 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15522 n7749 n7964 p_6_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15521 n7745 c_6_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15520 c_6_12_s1_s c_6_12_b n7745 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15519 vdd c_6_12_s1_s n7957 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15518 c_6_12_s2_s c_5_13_cout n7742 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15517 n7741 c_6_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15516 n7954 c_6_12_b n7741 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15515 n7954 c_5_13_cout n7740 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15514 vdd c_6_12_a n7740 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15513 n7740 c_6_12_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15512 c_8_11_cin n7954 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15511 n7742 n7957 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15510 c_8_10_a c_6_12_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15509 c_8_9_a c_6_11_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15508 n8320 n8316 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15507 c_6_11_cout n8321 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15506 n8314 c_6_11_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15505 vdd p_6_11_pi2j n8314 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15504 n8321 c_6_11_cin n8314 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15503 n8321 c_6_11_a n8319 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15502 n8319 p_6_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15501 c_6_11_s2_s c_6_11_cin n8320 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15500 vdd c_6_11_s1_s n8316 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15499 c_6_11_s1_s c_6_11_a n8317 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15498 n8317 p_6_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15497 n8329 p_6_2_d2j n8330 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15496 n8330 p_6_2_d2jbar n8331 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15495 n8331 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15494 vdd a_10 n8329 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15493 vdd p_6_11_t_s n8325 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15492 n8325 p_6_1_n2j p_6_11_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15491 vdd n8330 n8326 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15490 n8326 n8328 p_6_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15489 n8328 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15488 vdd n8713 n8505 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15487 n8504 p_6_1_n2j p_6_10_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15486 vdd p_6_10_t_s n8504 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15485 vdd a_8 n8506 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15484 n8507 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15483 n8716 p_6_2_d2j n8507 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15482 n8506 p_6_2_d2jbar n8716 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15481 n8713 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15480 n8505 n8716 p_6_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15479 n8503 c_6_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15478 c_6_10_s1_s p_6_10_pi2j n8503 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15477 vdd c_6_10_s1_s n8708 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15476 c_6_10_s2_s c_5_11_cout n8502 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15475 n8501 c_6_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15474 n8703 p_6_10_pi2j n8501 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15473 n8703 c_5_11_cout n8500 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15472 vdd c_6_10_a n8500 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15471 n8500 p_6_10_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15470 c_8_9_cin n8703 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15469 n8502 n8708 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15468 c_8_8_a c_6_10_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15467 c_8_7_a c_6_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15466 n9081 n9076 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15465 c_6_9_cout n9080 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15464 n9072 c_6_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15463 vdd p_6_9_pi2j n9072 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15462 n9080 c_6_9_cin n9072 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15461 n9080 c_6_9_a n9078 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15460 n9078 p_6_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15459 c_6_9_s2_s c_6_9_cin n9081 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15458 vdd c_6_9_s1_s n9076 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15457 c_6_9_s1_s c_6_9_a n9077 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15456 n9077 p_6_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15455 n9091 p_6_2_d2j n9090 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15454 n9090 p_6_2_d2jbar n9089 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15453 n9089 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15452 vdd a_8 n9091 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15451 vdd p_6_9_t_s n9084 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15450 n9084 p_6_1_n2j p_6_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15449 vdd n9090 n9087 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15448 n9087 n9088 p_6_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15447 n9088 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15446 vdd n9455 n9248 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15445 n9247 p_6_1_n2j p_6_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15444 vdd p_6_8_t_s n9247 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15443 vdd a_6 n9249 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15442 n9250 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15441 n9457 p_6_2_d2j n9250 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15440 n9249 p_6_2_d2jbar n9457 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15439 n9455 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15438 n9248 n9457 p_6_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15437 n9074 c_6_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15436 c_6_8_s1_s p_6_8_pi2j n9074 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15435 vdd c_6_8_s1_s n9450 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15434 c_6_8_s2_s c_5_9_cout n9246 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15433 n9075 c_6_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15432 n9445 p_6_8_pi2j n9075 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15431 n9445 c_5_9_cout n9245 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15430 vdd c_6_8_a n9245 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15429 n9245 p_6_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15428 c_8_7_cin n9445 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15427 n9246 n9450 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15426 c_8_6_a c_6_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15425 c_8_5_a c_6_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15424 n9868 n9864 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15423 c_6_7_cout n9869 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15422 n9860 c_6_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15421 vdd p_6_7_pi2j n9860 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15420 n9869 c_6_7_cin n9860 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15419 n9869 c_6_7_a n9867 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15418 n9867 p_6_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15417 c_6_7_s2_s c_6_7_cin n9868 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15416 vdd c_6_7_s1_s n9864 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15415 c_6_7_s1_s c_6_7_a n9865 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15414 n9865 p_6_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15413 n9586 p_6_2_d2j n9871 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15412 n9871 p_6_2_d2jbar n9587 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15411 n9587 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15410 vdd a_6 n9586 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15409 vdd p_6_7_t_s n9874 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15408 n9874 p_6_1_n2j p_6_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15407 vdd n9871 n9878 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15406 n9878 n9876 p_6_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15405 n9876 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15404 vdd n10231 n9879 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15403 n9873 p_6_1_n2j p_6_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15402 vdd p_6_6_t_s n9873 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15401 vdd a_4 n9880 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15400 n9881 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15399 n10230 p_6_2_d2j n9881 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15398 n9880 p_6_2_d2jbar n10230 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15397 n10231 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15396 n9879 n10230 p_6_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15395 n9863 c_6_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15394 c_6_6_s1_s p_6_6_pi2j n9863 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15393 vdd c_6_6_s1_s n10037 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15392 c_6_6_s2_s c_5_7_cout n10036 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15391 n9862 c_6_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15390 n10223 p_6_6_pi2j n9862 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15389 n10223 c_5_7_cout n10035 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15388 vdd c_6_6_a n10035 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15387 n10035 p_6_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15386 c_8_5_cin n10223 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15385 n10036 n10037 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15384 c_8_4_a c_6_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15383 c_8_3_a c_6_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15382 n10403 n10404 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15381 c_6_5_cout n10643 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15380 n10639 c_6_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15379 vdd c_6_5_b n10639 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15378 n10643 c_6_5_cin n10639 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15377 n10643 c_6_5_a n10644 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15376 n10644 c_6_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15375 c_6_5_s2_s c_6_5_cin n10403 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15374 vdd c_6_5_s1_s n10404 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15373 c_6_5_s1_s c_6_5_a n10641 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15372 n10641 c_6_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15371 n10409 p_6_2_d2j n10646 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15370 n10646 p_6_2_d2jbar n10410 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15369 n10410 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15368 vdd a_4 n10409 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15367 vdd p_6_5_t_s n10407 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15366 n10407 p_6_1_n2j c_6_5_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15365 vdd n10646 n10408 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15364 n10408 n10651 p_6_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15363 n10651 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15362 vdd n10841 n10652 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15361 n10649 p_6_1_n2j p_6_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15360 vdd p_6_4_t_s n10649 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15359 vdd a_2 n10653 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15358 n10654 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15357 n10844 p_6_2_d2j n10654 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15356 n10653 p_6_2_d2jbar n10844 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15355 n10841 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15354 n10652 n10844 p_6_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15353 n10642 c_6_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15352 c_6_4_s1_s p_6_4_pi2j n10642 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15351 vdd c_6_4_s1_s n10838 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15350 c_6_4_s2_s c_5_5_cout n10836 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15349 n10640 c_6_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15348 n10835 p_6_4_pi2j n10640 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15347 n10835 c_5_5_cout n10638 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15346 vdd c_6_4_a n10638 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15345 n10638 p_6_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15344 c_8_3_cin n10835 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15343 n10836 n10838 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15342 c_8_2_a c_6_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15341 c_8_1_a c_6_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15340 n11190 n11193 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15339 c_6_3_cout n11191 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15338 n11404 c_6_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15337 vdd c_6_3_b n11404 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15336 n11191 c_6_3_cin n11404 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15335 n11191 c_6_3_a n11410 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15334 n11410 c_6_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15333 c_6_3_s2_s c_6_3_cin n11190 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15332 vdd c_6_3_s1_s n11193 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15331 c_6_3_s1_s c_6_3_a n11408 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15330 n11408 c_6_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15329 n11200 p_6_2_d2j n11201 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15328 n11201 p_6_2_d2jbar n11202 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15327 n11202 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15326 vdd a_2 n11200 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15325 vdd p_6_3_t_s n11196 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15324 n11196 p_6_1_n2j c_6_3_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15323 vdd n11201 n11198 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15322 n11198 n11199 p_6_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15321 n11199 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15320 vdd n11624 n11414 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15319 n11412 p_6_1_n2j c_6_2_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15318 vdd p_6_2_t_s n11412 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15317 vdd a_0 n11415 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15316 n11416 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15315 n11627 p_6_2_d2j n11416 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15314 n11415 p_6_2_d2jbar n11627 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15313 n11624 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15312 n11414 n11627 p_6_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15311 n11409 c_6_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15310 c_6_2_s1_s c_6_2_b n11409 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15309 vdd c_6_2_s1_s n11620 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15308 c_6_2_s2_s c_5_3_cout n11407 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15307 n11406 c_6_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15306 n11617 c_6_2_b n11406 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15305 n11617 c_5_3_cout n11405 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15304 vdd c_6_2_a n11405 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15303 n11405 c_6_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15302 c_8_1_cin n11617 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15301 n11407 n11620 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15300 c_6_2_sum c_6_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15299 c_6_1_sum c_6_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15298 n11986 n11981 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15297 c_6_1_cout n11985 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15296 n11979 c_6_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15295 vdd p_6_1_pi2j n11979 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15294 n11985 c_6_1_cin n11979 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15293 n11985 c_6_1_a n11983 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15292 n11983 p_6_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15291 c_6_1_s2_s c_6_1_cin n11986 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15290 vdd c_6_1_s1_s n11981 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15289 c_6_1_s1_s c_6_1_a n11982 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15288 n11982 p_6_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15287 n11997 p_6_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15286 vdd a_0 n11997 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15285 vdd p_6_1_t_s n11991 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15284 n11991 p_6_1_n2j p_6_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15283 vdd n11997 n11993 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15282 n11993 n11995 p_6_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15281 n11995 p_6_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15280 n12139 c_5_1_sum cl4_6_s1_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15279 vdd n12357 n12139 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15278 p_8 cl4_6_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15277 n12348 c_5_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15276 vdd n12357 n12348 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15275 n12345 n12348 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15274 n12342 c_5_1_cout n12138 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15273 n12138 c_5_2_sum n12342 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15272 n12137 c_5_2_sum n12138 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_15271 vdd c_5_1_cout n12137 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_15270 n12138 c_5_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15269 vdd n12357 n12138 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15268 n12339 n12342 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15267 n12136 c_5_2_sum cl4_6_s2_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15266 vdd c_5_1_cout n12136 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15265 n12338 cl4_6_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_15264 n12135 n12345 cl4_6_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15263 vdd n12338 n12135 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15262 p_9 cl4_6_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15261 n209 p_5_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15260 c_5_33_s1_s c_5_31_a n209 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15259 vdd c_5_33_s1_s n205 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15258 c_5_33_s2_s c_5_32_cin n207 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15257 n203 p_5_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15256 n204 c_5_31_a n203 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15255 n204 c_5_32_cin n202 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15254 vdd p_5_33_pi2j n202 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15253 n202 c_5_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15252 c_6_32_cin n204 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15251 n207 n205 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15250 c_6_31_a c_5_33_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15249 n215 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15248 vdd p_5_33_t_s n211 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15247 n211 p_5_1_n2j p_5_33_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15246 vdd n215 n210 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15245 n210 n213 p_5_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15244 n213 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15243 vdd n552 n359 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15242 n358 p_5_1_n2j p_5_32_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15241 vdd p_5_32_t_s n358 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15240 vdd a_30 n360 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15239 n361 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15238 n554 p_5_2_d2j n361 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15237 n360 p_5_2_d2jbar n554 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15236 n552 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15235 n359 n554 p_5_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15234 n357 c_5_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15233 c_5_32_s1_s p_5_32_pi2j n357 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15232 vdd c_5_32_s1_s n549 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15231 c_5_32_s2_s c_5_32_cin n355 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15230 n356 c_5_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15229 n544 p_5_32_pi2j n356 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15228 n544 c_5_32_cin n354 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15227 vdd c_5_31_a n354 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15226 n354 p_5_32_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15225 c_6_31_cin n544 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15224 n355 n549 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15223 c_6_30_a c_5_32_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15222 c_6_29_a c_5_31_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15221 n903 n902 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15220 c_5_31_cout n906 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15219 n897 c_5_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15218 vdd p_5_31_pi2j n897 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15217 n906 c_5_31_cin n897 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15216 n906 c_5_31_a n904 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15215 n904 p_5_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15214 c_5_31_s2_s c_5_31_cin n903 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15213 vdd c_5_31_s1_s n902 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15212 c_5_31_s1_s c_5_31_a n900 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15211 n900 p_5_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15210 n913 p_5_2_d2j n911 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15209 n911 p_5_2_d2jbar n914 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15208 n914 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15207 vdd a_30 n913 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15206 vdd p_5_31_t_s n908 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15205 n908 p_5_1_n2j p_5_31_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15204 vdd n911 n907 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15203 n907 n912 p_5_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15202 n912 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15201 vdd n1312 n1081 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15200 n1080 p_5_1_n2j p_5_30_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15199 vdd p_5_30_t_s n1080 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15198 vdd a_28 n1082 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15197 n1083 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15196 n1314 p_5_2_d2j n1083 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15195 n1082 p_5_2_d2jbar n1314 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15194 n1312 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15193 n1081 n1314 p_5_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15192 n1079 c_5_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15191 c_5_30_s1_s p_5_30_pi2j n1079 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15190 vdd c_5_30_s1_s n1308 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15189 c_5_30_s2_s c_4_31_cout n1078 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15188 n1077 c_5_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15187 n1305 p_5_30_pi2j n1077 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15186 n1305 c_4_31_cout n1076 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15185 vdd c_5_30_a n1076 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15184 n1076 p_5_30_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15183 c_6_29_cin n1305 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15182 n1078 n1308 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15181 c_6_28_a c_5_30_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15180 c_6_27_a c_5_29_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15179 n1685 n1684 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15178 c_5_29_cout n1687 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15177 n1677 c_5_29_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15176 vdd p_5_29_pi2j n1677 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15175 n1687 c_5_29_cin n1677 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15174 n1687 c_5_29_a n1686 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15173 n1686 p_5_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15172 c_5_29_s2_s c_5_29_cin n1685 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15171 vdd c_5_29_s1_s n1684 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15170 c_5_29_s1_s c_5_29_a n1682 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15169 n1682 p_5_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15168 n1694 p_5_2_d2j n1693 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15167 n1693 p_5_2_d2jbar n1696 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15166 n1696 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15165 vdd a_28 n1694 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15164 vdd p_5_29_t_s n1689 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15163 n1689 p_5_1_n2j p_5_29_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15162 vdd n1693 n1690 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15161 n1690 n1695 p_5_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15160 n1695 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15159 vdd n2065 n1852 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15158 n1853 p_5_1_n2j p_5_28_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15157 vdd p_5_28_t_s n1853 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15156 vdd a_26 n1854 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15155 n1855 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15154 n2067 p_5_2_d2j n1855 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15153 n1854 p_5_2_d2jbar n2067 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15152 n2065 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15151 n1852 n2067 p_5_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15150 n1681 c_5_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15149 c_5_28_s1_s p_5_28_pi2j n1681 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15148 vdd c_5_28_s1_s n1851 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15147 c_5_28_s2_s c_4_29_cout n1850 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15146 n1680 c_5_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15145 n2057 p_5_28_pi2j n1680 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15144 n2057 c_4_29_cout n1849 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15143 vdd c_5_28_a n1849 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15142 n1849 p_5_28_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15141 c_6_27_cin n2057 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15140 n1850 n1851 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15139 c_6_26_a c_5_28_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15138 c_6_25_a c_5_27_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15137 n2212 n2491 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15136 c_5_27_cout n2498 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15135 n2490 c_5_27_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15134 vdd c_5_27_b n2490 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15133 n2498 c_5_27_cin n2490 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15132 n2498 c_5_27_a n2499 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15131 n2499 c_5_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15130 c_5_27_s2_s c_5_27_cin n2212 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15129 vdd c_5_27_s1_s n2491 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15128 c_5_27_s1_s c_5_27_a n2497 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15127 n2497 c_5_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15126 n2214 p_5_2_d2j n2501 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15125 n2501 p_5_2_d2jbar n2216 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15124 n2216 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15123 vdd a_26 n2214 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15122 vdd p_5_27_t_s n2213 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15121 n2213 p_5_1_n2j c_5_27_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15120 vdd n2501 n2504 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15119 n2504 n2505 p_5_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15118 n2505 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15117 vdd n2680 n2502 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15116 n2503 p_5_1_n2j p_5_26_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15115 vdd p_5_26_t_s n2503 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15114 vdd a_24 n2507 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15113 n2508 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15112 n2681 p_5_2_d2j n2508 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15111 n2507 p_5_2_d2jbar n2681 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15110 n2680 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15109 n2502 n2681 p_5_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15108 n2496 c_5_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15107 c_5_26_s1_s p_5_26_pi2j n2496 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15106 vdd c_5_26_s1_s n2679 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15105 c_5_26_s2_s c_4_27_cout n2678 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15104 n2495 c_5_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15103 n2868 p_5_26_pi2j n2495 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15102 n2868 c_4_27_cout n2676 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15101 vdd c_5_26_a n2676 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15100 n2676 p_5_26_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15099 c_6_25_cin n2868 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15098 n2678 n2679 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15097 c_6_24_a c_5_26_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15096 c_6_23_a c_5_25_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15095 n3038 n3039 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15094 c_5_25_cout n3284 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15093 n3277 c_5_25_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15092 vdd c_5_25_b n3277 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15091 n3284 c_5_25_cin n3277 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15090 n3284 c_5_25_a n3285 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15089 n3285 c_5_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15088 c_5_25_s2_s c_5_25_cin n3038 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15087 vdd c_5_25_s1_s n3039 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15086 c_5_25_s1_s c_5_25_a n3283 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15085 n3283 c_5_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15084 n3043 p_5_2_d2j n3042 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15083 n3042 p_5_2_d2jbar n3044 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15082 n3044 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15081 vdd a_24 n3043 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15080 vdd p_5_25_t_s n3041 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15079 n3041 p_5_1_n2j c_5_25_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15078 vdd n3042 n3040 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15077 n3040 n3288 p_5_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15076 n3288 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15075 vdd n3481 n3287 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15074 n3286 p_5_1_n2j c_5_24_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15073 vdd p_5_24_t_s n3286 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15072 vdd a_22 n3290 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15071 n3291 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15070 n3482 p_5_2_d2j n3291 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15069 n3290 p_5_2_d2jbar n3482 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15068 n3481 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15067 n3287 n3482 p_5_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15066 n3281 c_5_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15065 c_5_24_s1_s c_5_24_b n3281 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15064 vdd c_5_24_s1_s n3480 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15063 c_5_24_s2_s c_4_25_cout n3476 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15062 n3280 c_5_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15061 n3474 c_5_24_b n3280 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15060 n3474 c_4_25_cout n3276 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15059 vdd c_5_24_a n3276 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15058 n3276 c_5_24_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15057 c_6_23_cin n3474 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15056 n3476 n3480 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15055 c_6_22_a c_5_24_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15054 c_6_21_a c_5_23_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15053 n3872 n3875 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15052 c_5_23_cout n3873 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15051 n4060 c_5_23_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15050 vdd c_5_23_b n4060 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15049 n3873 c_5_23_cin n4060 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15048 n3873 c_5_23_a n3871 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15047 n3871 c_5_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15046 c_5_23_s2_s c_5_23_cin n3872 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15045 vdd c_5_23_s1_s n3875 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15044 c_5_23_s1_s c_5_23_a n3869 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15043 n3869 c_5_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15042 n3881 p_5_2_d2j n3879 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15041 n3879 p_5_2_d2jbar n3882 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15040 n3882 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15039 vdd a_22 n3881 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15038 vdd p_5_23_t_s n3877 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15037 n3877 p_5_1_n2j c_5_23_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15036 vdd n3879 n3876 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15035 n3876 n3880 p_5_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15034 n3880 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15033 vdd n4291 n4066 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15032 n4065 p_5_1_n2j p_5_22_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15031 vdd p_5_22_t_s n4065 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15030 vdd a_20 n4067 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15029 n4068 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_15028 n4293 p_5_2_d2j n4068 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15027 n4067 p_5_2_d2jbar n4293 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_15026 n4291 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15025 n4066 n4293 p_5_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_15024 n4064 c_5_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15023 c_5_22_s1_s p_5_22_pi2j n4064 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15022 vdd c_5_22_s1_s n4289 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15021 c_5_22_s2_s c_4_23_cout n4062 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15020 n4063 c_5_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15019 n4283 p_5_22_pi2j n4063 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15018 n4283 c_4_23_cout n4059 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15017 vdd c_5_22_a n4059 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15016 n4059 p_5_22_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15015 c_6_21_cin n4283 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15014 n4062 n4289 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15013 c_6_20_a c_5_22_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15012 c_6_19_a c_5_21_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15011 n4652 n4647 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_15010 c_5_21_cout n4650 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_15009 n4644 c_5_21_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15008 vdd p_5_21_pi2j n4644 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15007 n4650 c_5_21_cin n4644 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15006 n4650 c_5_21_a n4653 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15005 n4653 p_5_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15004 c_5_21_s2_s c_5_21_cin n4652 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_15003 vdd c_5_21_s1_s n4647 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_15002 c_5_21_s1_s c_5_21_a n4648 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15001 n4648 p_5_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_15000 n4660 p_5_2_d2j n4658 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14999 n4658 p_5_2_d2jbar n4661 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14998 n4661 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14997 vdd a_20 n4660 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14996 vdd p_5_21_t_s n4655 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14995 n4655 p_5_1_n2j p_5_21_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14994 vdd n4658 n4654 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14993 n4654 n4659 p_5_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14992 n4659 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14991 vdd n5037 n4824 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14990 n4823 p_5_1_n2j p_5_20_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14989 vdd p_5_20_t_s n4823 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14988 vdd a_18 n4825 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14987 n4826 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14986 n5039 p_5_2_d2j n4826 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14985 n4825 p_5_2_d2jbar n5039 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14984 n5037 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14983 n4824 n5039 p_5_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14982 n4822 c_5_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14981 c_5_20_s1_s p_5_20_pi2j n4822 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14980 vdd c_5_20_s1_s n5035 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14979 c_5_20_s2_s c_4_21_cout n4821 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14978 n4820 c_5_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14977 n5029 p_5_20_pi2j n4820 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14976 n5029 c_4_21_cout n4819 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14975 vdd c_5_20_a n4819 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14974 n4819 p_5_20_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14973 c_6_19_cin n5029 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14972 n4821 n5035 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14971 c_6_18_a c_5_20_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14970 c_6_17_a c_5_19_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14969 n5412 n5411 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14968 c_5_19_cout n5415 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14967 n5404 c_5_19_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14966 vdd p_5_19_pi2j n5404 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14965 n5415 c_5_19_cin n5404 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14964 n5415 c_5_19_a n5413 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14963 n5413 p_5_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14962 c_5_19_s2_s c_5_19_cin n5412 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14961 vdd c_5_19_s1_s n5411 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14960 c_5_19_s1_s c_5_19_a n5409 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14959 n5409 p_5_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14958 n5421 p_5_2_d2j n5420 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14957 n5420 p_5_2_d2jbar n5423 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14956 n5423 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14955 vdd a_18 n5421 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14954 vdd p_5_19_t_s n5416 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14953 n5416 p_5_1_n2j p_5_19_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14952 vdd n5420 n5417 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14951 n5417 n5422 p_5_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14950 n5422 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14949 vdd n5792 n5579 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14948 n5578 p_5_1_n2j p_5_18_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14947 vdd p_5_18_t_s n5578 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14946 vdd a_16 n5580 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14945 n5581 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14944 n5791 p_5_2_d2j n5581 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14943 n5580 p_5_2_d2jbar n5791 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14942 n5792 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14941 n5579 n5791 p_5_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14940 n5407 c_5_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14939 c_5_18_s1_s p_5_18_pi2j n5407 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14938 vdd c_5_18_s1_s n5577 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14937 c_5_18_s2_s c_4_19_cout n5576 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14936 n5408 c_5_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14935 n5782 p_5_18_pi2j n5408 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14934 n5782 c_4_19_cout n5575 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14933 vdd c_5_18_a n5575 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14932 n5575 p_5_18_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14931 c_6_17_cin n5782 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14930 n5576 n5577 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14929 c_6_16_a c_5_18_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14928 c_6_15_a c_5_17_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14927 n6207 n6199 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14926 c_5_17_cout n6209 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14925 n6198 c_5_17_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14924 vdd p_5_17_pi2j n6198 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14923 n6209 c_5_17_cin n6198 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14922 n6209 c_5_17_a n6208 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14921 n6208 p_5_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14920 c_5_17_s2_s c_5_17_cin n6207 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14919 vdd c_5_17_s1_s n6199 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14918 c_5_17_s1_s c_5_17_a n6204 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14917 n6204 p_5_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14916 n5913 p_5_2_d2j n6210 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14915 n6210 p_5_2_d2jbar n5915 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14914 n5915 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14913 vdd a_16 n5913 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14912 vdd p_5_17_t_s n6213 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14911 n6213 p_5_1_n2j p_5_17_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14910 vdd n6210 n6214 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14909 n6214 n6216 p_5_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14908 n6216 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14907 vdd n6572 n6211 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14906 n6212 p_5_1_n2j p_5_16_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14905 vdd p_5_16_t_s n6212 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14904 vdd a_14 n6218 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14903 n6219 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14902 n6380 p_5_2_d2j n6219 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14901 n6218 p_5_2_d2jbar n6380 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14900 n6572 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14899 n6211 n6380 p_5_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14898 n6203 c_5_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14897 c_5_16_s1_s p_5_16_pi2j n6203 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14896 vdd c_5_16_s1_s n6379 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14895 c_5_16_s2_s c_4_17_cout n6378 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14894 n6202 c_5_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14893 n6565 p_5_16_pi2j n6202 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14892 n6565 c_4_17_cout n6376 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14891 vdd c_5_16_a n6376 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14890 n6376 p_5_16_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14889 c_6_15_cin n6565 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14888 n6378 n6379 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14887 c_6_14_a c_5_16_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14886 c_6_13_a c_5_15_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14885 n6739 n6740 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14884 c_5_15_cout n6987 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14883 n6979 c_5_15_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14882 vdd c_5_15_b n6979 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14881 n6987 c_5_15_cin n6979 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14880 n6987 c_5_15_a n6984 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14879 n6984 c_5_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14878 c_5_15_s2_s c_5_15_cin n6739 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14877 vdd c_5_15_s1_s n6740 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14876 c_5_15_s1_s c_5_15_a n6985 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14875 n6985 c_5_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14874 n6744 p_5_2_d2j n6743 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14873 n6743 p_5_2_d2jbar n6745 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14872 n6745 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14871 vdd a_14 n6744 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14870 vdd p_5_15_t_s n6742 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14869 n6742 p_5_1_n2j c_5_15_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14868 vdd n6743 n6741 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14867 n6741 n6990 p_5_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14866 n6990 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14865 vdd n7177 n6989 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14864 n6988 p_5_1_n2j p_5_14_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14863 vdd p_5_14_t_s n6988 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14862 vdd a_12 n6992 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14861 n6993 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14860 n7178 p_5_2_d2j n6993 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14859 n6992 p_5_2_d2jbar n7178 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14858 n7177 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14857 n6989 n7178 p_5_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14856 n6983 c_5_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14855 c_5_14_s1_s p_5_14_pi2j n6983 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14854 vdd c_5_14_s1_s n7176 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14853 c_5_14_s2_s c_4_15_cout n7172 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14852 n6982 c_5_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14851 n7171 p_5_14_pi2j n6982 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14850 n7171 c_4_15_cout n6978 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14849 vdd c_5_14_a n6978 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14848 n6978 p_5_14_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14847 c_6_13_cin n7171 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14846 n7172 n7176 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14845 c_6_12_a c_5_14_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14844 c_6_11_a c_5_13_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14843 n7540 n7544 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14842 c_5_13_cout n7542 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14841 n7753 c_5_13_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14840 vdd c_5_13_b n7753 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14839 n7542 c_5_13_cin n7753 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14838 n7542 c_5_13_a n7758 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14837 n7758 c_5_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14836 c_5_13_s2_s c_5_13_cin n7540 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14835 vdd c_5_13_s1_s n7544 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14834 c_5_13_s1_s c_5_13_a n7759 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14833 n7759 c_5_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14832 n7549 p_5_2_d2j n7547 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14831 n7547 p_5_2_d2jbar n7550 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14830 n7550 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14829 vdd a_12 n7549 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14828 vdd p_5_13_t_s n7546 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14827 n7546 p_5_1_n2j c_5_13_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14826 vdd n7547 n7545 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14825 n7545 n7548 p_5_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14824 n7548 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14823 vdd n7973 n7761 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14822 n7760 p_5_1_n2j c_5_12_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14821 vdd p_5_12_t_s n7760 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14820 vdd a_10 n7763 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14819 n7764 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14818 n7975 p_5_2_d2j n7764 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14817 n7763 p_5_2_d2jbar n7975 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14816 n7973 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14815 n7761 n7975 p_5_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14814 n7757 c_5_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14813 c_5_12_s1_s c_5_12_b n7757 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14812 vdd c_5_12_s1_s n7972 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14811 c_5_12_s2_s c_4_13_cout n7755 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14810 n7756 c_5_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14809 n7967 c_5_12_b n7756 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14808 n7967 c_4_13_cout n7752 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14807 vdd c_5_12_a n7752 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14806 n7752 c_5_12_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14805 c_6_11_cin n7967 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14804 n7755 n7972 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14803 c_6_10_a c_5_12_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14802 c_6_9_a c_5_11_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14801 n8339 n8335 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14800 c_5_11_cout n8340 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14799 n8332 c_5_11_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14798 vdd p_5_11_pi2j n8332 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14797 n8340 c_5_11_cin n8332 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14796 n8340 c_5_11_a n8338 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14795 n8338 p_5_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14794 c_5_11_s2_s c_5_11_cin n8339 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14793 vdd c_5_11_s1_s n8335 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14792 c_5_11_s1_s c_5_11_a n8336 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14791 n8336 p_5_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14790 n8348 p_5_2_d2j n8346 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14789 n8346 p_5_2_d2jbar n8349 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14788 n8349 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14787 vdd a_10 n8348 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14786 vdd p_5_11_t_s n8343 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14785 n8343 p_5_1_n2j p_5_11_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14784 vdd n8346 n8342 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14783 n8342 n8347 p_5_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14782 n8347 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14781 vdd n8726 n8513 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14780 n8512 p_5_1_n2j p_5_10_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14779 vdd p_5_10_t_s n8512 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14778 vdd a_8 n8514 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14777 n8515 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14776 n8728 p_5_2_d2j n8515 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14775 n8514 p_5_2_d2jbar n8728 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14774 n8726 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14773 n8513 n8728 p_5_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14772 n8511 c_5_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14771 c_5_10_s1_s p_5_10_pi2j n8511 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14770 vdd c_5_10_s1_s n8722 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14769 c_5_10_s2_s c_4_11_cout n8510 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14768 n8509 c_5_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14767 n8718 p_5_10_pi2j n8509 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14766 n8718 c_4_11_cout n8508 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14765 vdd c_5_10_a n8508 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14764 n8508 p_5_10_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14763 c_6_9_cin n8718 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14762 n8510 n8722 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14761 c_6_8_a c_5_10_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14760 c_6_7_a c_5_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14759 n9100 n9099 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14758 c_5_9_cout n9103 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14757 n9092 c_5_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14756 vdd p_5_9_pi2j n9092 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14755 n9103 c_5_9_cin n9092 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14754 n9103 c_5_9_a n9101 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14753 n9101 p_5_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14752 c_5_9_s2_s c_5_9_cin n9100 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14751 vdd c_5_9_s1_s n9099 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14750 c_5_9_s1_s c_5_9_a n9097 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14749 n9097 p_5_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14748 n9109 p_5_2_d2j n9108 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14747 n9108 p_5_2_d2jbar n9111 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14746 n9111 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14745 vdd a_8 n9109 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14744 vdd p_5_9_t_s n9104 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14743 n9104 p_5_1_n2j p_5_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14742 vdd n9108 n9105 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14741 n9105 n9110 p_5_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14740 n9110 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14739 vdd n9471 n9254 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14738 n9253 p_5_1_n2j p_5_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14737 vdd p_5_8_t_s n9253 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14736 vdd a_6 n9255 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14735 n9256 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14734 n9470 p_5_2_d2j n9256 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14733 n9255 p_5_2_d2jbar n9470 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14732 n9471 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14731 n9254 n9470 p_5_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14730 n9095 c_5_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14729 c_5_8_s1_s p_5_8_pi2j n9095 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14728 vdd c_5_8_s1_s n9459 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14727 c_5_8_s2_s c_4_9_cout n9252 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14726 n9096 c_5_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14725 n9461 p_5_8_pi2j n9096 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14724 n9461 c_4_9_cout n9251 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14723 vdd c_5_8_a n9251 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14722 n9251 p_5_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14721 c_6_7_cin n9461 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14720 n9252 n9459 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14719 c_6_6_a c_5_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14718 c_6_5_a c_5_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14717 n9891 n9887 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14716 c_5_7_cout n9892 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14715 n9882 c_5_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14714 vdd p_5_7_pi2j n9882 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14713 n9892 c_5_7_cin n9882 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14712 n9892 c_5_7_a n9890 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14711 n9890 p_5_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14710 c_5_7_s2_s c_5_7_cin n9891 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14709 vdd c_5_7_s1_s n9887 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14708 c_5_7_s1_s c_5_7_a n9888 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14707 n9888 p_5_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14706 n9591 p_5_2_d2j n9894 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14705 n9894 p_5_2_d2jbar n9593 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14704 n9593 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14703 vdd a_6 n9591 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14702 vdd p_5_7_t_s n9897 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14701 n9897 p_5_1_n2j p_5_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14700 vdd n9894 n9898 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14699 n9898 n9900 p_5_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14698 n9900 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14697 vdd n10245 n9895 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14696 n9896 p_5_1_n2j p_5_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14695 vdd p_5_6_t_s n9896 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14694 vdd a_4 n9902 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14693 n9903 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14692 n10244 p_5_2_d2j n9903 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14691 n9902 p_5_2_d2jbar n10244 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14690 n10245 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14689 n9895 n10244 p_5_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14688 n9886 c_5_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14687 c_5_6_s1_s p_5_6_pi2j n9886 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14686 vdd c_5_6_s1_s n10042 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14685 c_5_6_s2_s c_4_7_cout n10041 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14684 n9885 c_5_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14683 n10237 p_5_6_pi2j n9885 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14682 n10237 c_4_7_cout n10040 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14681 vdd c_5_6_a n10040 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14680 n10040 p_5_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14679 c_6_5_cin n10237 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14678 n10041 n10042 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14677 c_6_4_a c_5_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14676 c_6_3_a c_5_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14675 n10413 n10415 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14674 c_5_5_cout n10662 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14673 n10656 c_5_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14672 vdd c_5_5_b n10656 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14671 n10662 c_5_5_cin n10656 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14670 n10662 c_5_5_a n10663 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14669 n10663 c_5_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14668 c_5_5_s2_s c_5_5_cin n10413 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14667 vdd c_5_5_s1_s n10415 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14666 c_5_5_s1_s c_5_5_a n10661 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14665 n10661 c_5_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14664 n10418 p_5_2_d2j n10665 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14663 n10665 p_5_2_d2jbar n10419 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14662 n10419 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14661 vdd a_4 n10418 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14660 vdd p_5_5_t_s n10417 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14659 n10417 p_5_1_n2j c_5_5_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14658 vdd n10665 n10416 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14657 n10416 n10668 p_5_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14656 n10668 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14655 vdd n10851 n10667 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14654 n10666 p_5_1_n2j p_5_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14653 vdd p_5_4_t_s n10666 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14652 vdd a_2 n10670 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14651 n10671 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14650 n10852 p_5_2_d2j n10671 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14649 n10670 p_5_2_d2jbar n10852 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14648 n10851 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14647 n10667 n10852 p_5_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14646 n10660 c_5_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14645 c_5_4_s1_s p_5_4_pi2j n10660 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14644 vdd c_5_4_s1_s n10850 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14643 c_5_4_s2_s c_4_5_cout n10847 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14642 n10659 c_5_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14641 n10845 p_5_4_pi2j n10659 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14640 n10845 c_4_5_cout n10655 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14639 vdd c_5_4_a n10655 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14638 n10655 p_5_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14637 c_6_3_cin n10845 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14636 n10847 n10850 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14635 c_6_2_a c_5_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14634 c_6_1_a c_5_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14633 n11205 n11209 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14632 c_5_3_cout n11207 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14631 n11418 c_5_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14630 vdd c_5_3_b n11418 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14629 n11207 c_5_3_cin n11418 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14628 n11207 c_5_3_a n11424 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14627 n11424 c_5_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14626 c_5_3_s2_s c_5_3_cin n11205 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14625 vdd c_5_3_s1_s n11209 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14624 c_5_3_s1_s c_5_3_a n11423 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14623 n11423 c_5_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14622 n11214 p_5_2_d2j n11212 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14621 n11212 p_5_2_d2jbar n11215 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14620 n11215 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14619 vdd a_2 n11214 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14618 vdd p_5_3_t_s n11211 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14617 n11211 p_5_1_n2j c_5_3_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14616 vdd n11212 n11210 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14615 n11210 n11213 p_5_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14614 n11213 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14613 vdd n11636 n11426 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14612 n11425 p_5_1_n2j c_5_2_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14611 vdd p_5_2_t_s n11425 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14610 vdd a_0 n11428 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14609 n11429 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14608 n11638 p_5_2_d2j n11429 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14607 n11428 p_5_2_d2jbar n11638 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14606 n11636 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14605 n11426 n11638 p_5_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14604 n11422 c_5_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14603 c_5_2_s1_s c_5_2_b n11422 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14602 vdd c_5_2_s1_s n11635 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14601 c_5_2_s2_s c_4_3_cout n11420 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14600 n11421 c_5_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14599 n11629 c_5_2_b n11421 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14598 n11629 c_4_3_cout n11417 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14597 vdd c_5_2_a n11417 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14596 n11417 c_5_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14595 c_6_1_cin n11629 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14594 n11420 n11635 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14593 c_5_2_sum c_5_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14592 c_5_1_sum c_5_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14591 n12006 n12001 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14590 c_5_1_cout n12004 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14589 n11998 c_5_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14588 vdd p_5_1_pi2j n11998 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14587 n12004 c_5_1_cin n11998 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14586 n12004 c_5_1_a n12007 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14585 n12007 p_5_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14584 c_5_1_s2_s c_5_1_cin n12006 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14583 vdd c_5_1_s1_s n12001 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14582 c_5_1_s1_s c_5_1_a n12002 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14581 n12002 p_5_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14580 n12014 p_5_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14579 vdd a_0 n12014 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14578 vdd p_5_1_t_s n12010 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14577 n12010 p_5_1_n2j p_5_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14576 vdd n12014 n12009 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14575 n12009 n12015 p_5_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14574 n12015 p_5_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14573 n12144 c_4_1_sum cl4_5_s1_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14572 vdd n12375 n12144 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14571 p_6 cl4_5_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14570 n12364 c_4_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14569 vdd n12375 n12364 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14568 n12363 n12364 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14567 n12361 c_4_1_cout n12143 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14566 n12143 c_4_2_sum n12361 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14565 n12142 c_4_2_sum n12143 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_14564 vdd c_4_1_cout n12142 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_14563 n12143 c_4_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14562 vdd n12375 n12143 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14561 n12357 n12361 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14560 n12141 c_4_2_sum cl4_5_s2_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14559 vdd c_4_1_cout n12141 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14558 n12356 cl4_5_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_14557 n12140 n12363 cl4_5_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14556 vdd n12356 n12140 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14555 p_7 cl4_5_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14554 n222 p_4_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14553 c_4_33_s1_s c_4_31_a n222 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14552 vdd c_4_33_s1_s n223 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14551 c_4_33_s2_s c_4_32_cin n221 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14550 n219 p_4_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14549 n220 c_4_31_a n219 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14548 n220 c_4_32_cin n216 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14547 vdd p_4_33_pi2j n216 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14546 n216 c_4_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14545 c_5_32_cin n220 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14544 n221 n223 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14543 c_5_31_a c_4_33_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14542 n229 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14541 vdd p_4_33_t_s n218 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14540 n218 p_4_1_n2j p_4_33_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14539 vdd n229 n225 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14538 n225 n228 p_4_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14537 n228 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14536 vdd n565 n367 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14535 n365 p_4_1_n2j p_4_32_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14534 vdd p_4_32_t_s n365 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14533 vdd a_30 n368 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14532 n369 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14531 n568 p_4_2_d2j n369 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14530 n368 p_4_2_d2jbar n568 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14529 n565 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14528 n367 n568 p_4_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14527 n366 c_4_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14526 c_4_32_s1_s p_4_32_pi2j n366 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14525 vdd c_4_32_s1_s n561 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14524 c_4_32_s2_s c_4_32_cin n364 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14523 n363 c_4_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14522 n558 p_4_32_pi2j n363 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14521 n558 c_4_32_cin n362 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14520 vdd c_4_31_a n362 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14519 n362 p_4_32_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14518 c_5_31_cin n558 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14517 n364 n561 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14516 c_5_30_a c_4_32_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14515 c_5_29_a c_4_31_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14514 n923 n922 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14513 c_4_31_cout n925 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14512 n916 c_4_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14511 vdd p_4_31_pi2j n916 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14510 n925 c_4_31_cin n916 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14509 n925 c_4_31_a n924 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14508 n924 p_4_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14507 c_4_31_s2_s c_4_31_cin n923 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14506 vdd c_4_31_s1_s n922 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14505 c_4_31_s1_s c_4_31_a n919 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14504 n919 p_4_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14503 n931 p_4_2_d2j n929 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14502 n929 p_4_2_d2jbar n930 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14501 n930 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14500 vdd a_30 n931 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14499 vdd p_4_31_t_s n920 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14498 n920 p_4_1_n2j p_4_31_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14497 vdd n929 n926 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14496 n926 n932 p_4_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14495 n932 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14494 vdd n1328 n1089 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14493 n1088 p_4_1_n2j p_4_30_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14492 vdd p_4_30_t_s n1088 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14491 vdd a_28 n1090 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14490 n1091 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14489 n1331 p_4_2_d2j n1091 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14488 n1090 p_4_2_d2jbar n1331 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14487 n1328 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14486 n1089 n1331 p_4_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14485 n1087 c_4_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14484 c_4_30_s1_s p_4_30_pi2j n1087 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14483 vdd c_4_30_s1_s n1325 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14482 c_4_30_s2_s c_3_31_cout n1085 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14481 n1086 c_4_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14480 n1318 p_4_30_pi2j n1086 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14479 n1318 c_3_31_cout n1084 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14478 vdd c_4_30_a n1084 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14477 n1084 p_4_30_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14476 c_5_29_cin n1318 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14475 n1085 n1325 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14474 c_5_28_a c_4_30_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14473 c_5_27_a c_4_29_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14472 n1708 n1704 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14471 c_4_29_cout n1709 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14470 n1698 c_4_29_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14469 vdd p_4_29_pi2j n1698 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14468 n1709 c_4_29_cin n1698 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14467 n1709 c_4_29_a n1707 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14466 n1707 p_4_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14465 c_4_29_s2_s c_4_29_cin n1708 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14464 vdd c_4_29_s1_s n1704 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14463 c_4_29_s1_s c_4_29_a n1705 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14462 n1705 p_4_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14461 n1715 p_4_2_d2j n1714 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14460 n1714 p_4_2_d2jbar n1713 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14459 n1713 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14458 vdd a_28 n1715 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14457 vdd p_4_29_t_s n1703 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14456 n1703 p_4_1_n2j p_4_29_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14455 vdd n1714 n1710 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14454 n1710 n1716 p_4_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14453 n1716 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14452 vdd n2082 n1860 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14451 n1858 p_4_1_n2j p_4_28_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14450 vdd p_4_28_t_s n1858 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14449 vdd a_26 n1862 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14448 n1861 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14447 n2081 p_4_2_d2j n1861 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14446 n1862 p_4_2_d2jbar n2081 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14445 n2082 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14444 n1860 n2081 p_4_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14443 n1702 c_4_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14442 c_4_28_s1_s p_4_28_pi2j n1702 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14441 vdd c_4_28_s1_s n1859 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14440 c_4_28_s2_s c_3_29_cout n1857 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14439 n1701 c_4_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14438 n2071 p_4_28_pi2j n1701 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14437 n2071 c_3_29_cout n1856 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14436 vdd c_4_28_a n1856 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14435 n1856 p_4_28_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14434 c_5_27_cin n2071 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14433 n1857 n1859 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14432 c_5_26_a c_4_28_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14431 c_5_25_a c_4_27_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14430 n2220 n2511 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14429 c_4_27_cout n2521 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14428 n2510 c_4_27_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14427 vdd c_4_27_b n2510 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14426 n2521 c_4_27_cin n2510 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14425 n2521 c_4_27_a n2520 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14424 n2520 c_4_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14423 c_4_27_s2_s c_4_27_cin n2220 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14422 vdd c_4_27_s1_s n2511 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14421 c_4_27_s1_s c_4_27_a n2519 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14420 n2519 c_4_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14419 n2222 p_4_2_d2j n2522 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14418 n2522 p_4_2_d2jbar n2221 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14417 n2221 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14416 vdd a_26 n2222 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14415 vdd p_4_27_t_s n2219 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14414 n2219 p_4_1_n2j c_4_27_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14413 vdd n2522 n2524 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14412 n2524 n2526 p_4_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14411 n2526 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14410 vdd n2688 n2525 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14409 n2516 p_4_1_n2j p_4_26_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14408 vdd p_4_26_t_s n2516 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14407 vdd a_24 n2527 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14406 n2528 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14405 n2691 p_4_2_d2j n2528 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14404 n2527 p_4_2_d2jbar n2691 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14403 n2688 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14402 n2525 n2691 p_4_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14401 n2517 c_4_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14400 c_4_26_s1_s p_4_26_pi2j n2517 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14399 vdd c_4_26_s1_s n2687 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14398 c_4_26_s2_s c_3_27_cout n2686 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14397 n2515 c_4_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14396 n2883 p_4_26_pi2j n2515 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14395 n2883 c_3_27_cout n2684 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14394 vdd c_4_26_a n2684 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14393 n2684 p_4_26_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14392 c_5_25_cin n2883 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14391 n2686 n2687 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14390 c_5_24_a c_4_26_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14389 c_5_23_a c_4_25_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14388 n3048 n3049 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14387 c_4_25_cout n3302 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14386 n3293 c_4_25_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14385 vdd c_4_25_b n3293 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14384 n3302 c_4_25_cin n3293 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14383 n3302 c_4_25_a n3301 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14382 n3301 c_4_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14381 c_4_25_s2_s c_4_25_cin n3048 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14380 vdd c_4_25_s1_s n3049 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14379 c_4_25_s1_s c_4_25_a n3300 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14378 n3300 c_4_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14377 n3053 p_4_2_d2j n3051 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14376 n3051 p_4_2_d2jbar n3052 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14375 n3052 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14374 vdd a_24 n3053 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14373 vdd p_4_25_t_s n3047 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14372 n3047 p_4_1_n2j c_4_25_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14371 vdd n3051 n3050 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14370 n3050 n3305 p_4_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14369 n3305 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14368 vdd n3492 n3304 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14367 n3297 p_4_1_n2j c_4_24_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14366 vdd p_4_24_t_s n3297 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14365 vdd a_22 n3306 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14364 n3307 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14363 n3495 p_4_2_d2j n3307 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14362 n3306 p_4_2_d2jbar n3495 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14361 n3492 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14360 n3304 n3495 p_4_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14359 n3298 c_4_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14358 c_4_24_s1_s c_4_24_b n3298 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14357 vdd c_4_24_s1_s n3489 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14356 c_4_24_s2_s c_3_25_cout n3488 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14355 n3296 c_4_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14354 n3485 c_4_24_b n3296 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14353 n3485 c_3_25_cout n3292 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14352 vdd c_4_24_a n3292 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14351 n3292 c_4_24_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14350 c_5_23_cin n3485 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14349 n3488 n3489 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14348 c_5_22_a c_4_24_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14347 c_5_21_a c_4_23_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14346 n3889 n3892 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14345 c_4_23_cout n3891 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14344 n4070 c_4_23_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14343 vdd c_4_23_b n4070 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14342 n3891 c_4_23_cin n4070 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14341 n3891 c_4_23_a n3888 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14340 n3888 c_4_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14339 c_4_23_s2_s c_4_23_cin n3889 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14338 vdd c_4_23_s1_s n3892 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14337 c_4_23_s1_s c_4_23_a n3887 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14336 n3887 c_4_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14335 n3897 p_4_2_d2j n3895 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14334 n3895 p_4_2_d2jbar n3896 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14333 n3896 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14332 vdd a_22 n3897 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14331 vdd p_4_23_t_s n3886 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14330 n3886 p_4_1_n2j c_4_23_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14329 vdd n3895 n3893 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14328 n3893 n3898 p_4_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14327 n3898 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14326 vdd n4306 n4076 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14325 n4074 p_4_1_n2j p_4_22_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14324 vdd p_4_22_t_s n4074 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14323 vdd a_20 n4077 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14322 n4078 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14321 n4309 p_4_2_d2j n4078 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14320 n4077 p_4_2_d2jbar n4309 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14319 n4306 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14318 n4076 n4309 p_4_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14317 n4075 c_4_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14316 c_4_22_s1_s p_4_22_pi2j n4075 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14315 vdd c_4_22_s1_s n4301 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14314 c_4_22_s2_s c_3_23_cout n4073 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14313 n4072 c_4_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14312 n4298 p_4_22_pi2j n4072 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14311 n4298 c_3_23_cout n4069 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14310 vdd c_4_22_a n4069 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14309 n4069 p_4_22_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14308 c_5_21_cin n4298 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14307 n4073 n4301 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14306 c_5_20_a c_4_22_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14305 c_5_19_a c_4_21_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14304 n4672 n4667 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14303 c_4_21_cout n4671 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14302 n4663 c_4_21_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14301 vdd p_4_21_pi2j n4663 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14300 n4671 c_4_21_cin n4663 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14299 n4671 c_4_21_a n4669 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14298 n4669 p_4_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14297 c_4_21_s2_s c_4_21_cin n4672 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14296 vdd c_4_21_s1_s n4667 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14295 c_4_21_s1_s c_4_21_a n4668 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14294 n4668 p_4_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14293 n4678 p_4_2_d2j n4676 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14292 n4676 p_4_2_d2jbar n4677 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14291 n4677 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14290 vdd a_20 n4678 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14289 vdd p_4_21_t_s n4666 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14288 n4666 p_4_1_n2j p_4_21_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14287 vdd n4676 n4673 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14286 n4673 n4679 p_4_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14285 n4679 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14284 vdd n5052 n4832 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14283 n4831 p_4_1_n2j p_4_20_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14282 vdd p_4_20_t_s n4831 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14281 vdd a_18 n4833 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14280 n4834 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14279 n5055 p_4_2_d2j n4834 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14278 n4833 p_4_2_d2jbar n5055 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14277 n5052 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14276 n4832 n5055 p_4_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14275 n4830 c_4_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14274 c_4_20_s1_s p_4_20_pi2j n4830 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14273 vdd c_4_20_s1_s n5048 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14272 c_4_20_s2_s c_3_21_cout n4828 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14271 n4829 c_4_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14270 n5042 p_4_20_pi2j n4829 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14269 n5042 c_3_21_cout n4827 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14268 vdd c_4_20_a n4827 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14267 n4827 p_4_20_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14266 c_5_19_cin n5042 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14265 n4828 n5048 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14264 c_5_18_a c_4_20_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14263 c_5_17_a c_4_19_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14262 n5435 n5431 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14261 c_4_19_cout n5436 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14260 n5425 c_4_19_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14259 vdd p_4_19_pi2j n5425 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14258 n5436 c_4_19_cin n5425 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14257 n5436 c_4_19_a n5434 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14256 n5434 p_4_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14255 c_4_19_s2_s c_4_19_cin n5435 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14254 vdd c_4_19_s1_s n5431 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14253 c_4_19_s1_s c_4_19_a n5432 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14252 n5432 p_4_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14251 n5442 p_4_2_d2j n5441 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14250 n5441 p_4_2_d2jbar n5440 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14249 n5440 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14248 vdd a_18 n5442 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14247 vdd p_4_19_t_s n5430 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14246 n5430 p_4_1_n2j p_4_19_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14245 vdd n5441 n5437 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14244 n5437 n5443 p_4_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14243 n5443 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14242 vdd n5806 n5586 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14241 n5584 p_4_1_n2j p_4_18_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14240 vdd p_4_18_t_s n5584 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14239 vdd a_16 n5587 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14238 n5588 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14237 n5808 p_4_2_d2j n5588 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14236 n5587 p_4_2_d2jbar n5808 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14235 n5806 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14234 n5586 n5808 p_4_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14233 n5429 c_4_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14232 c_4_18_s1_s p_4_18_pi2j n5429 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14231 vdd c_4_18_s1_s n5585 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14230 c_4_18_s2_s c_3_19_cout n5583 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14229 n5428 c_4_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14228 n5799 p_4_18_pi2j n5428 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14227 n5799 c_3_19_cout n5582 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14226 vdd c_4_18_a n5582 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14225 n5582 p_4_18_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14224 c_5_17_cin n5799 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14223 n5583 n5585 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14222 c_5_16_a c_4_18_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14221 c_5_15_a c_4_17_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14220 n6231 n6222 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14219 c_4_17_cout n6233 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14218 n6221 c_4_17_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14217 vdd p_4_17_pi2j n6221 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14216 n6233 c_4_17_cin n6221 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14215 n6233 c_4_17_a n6232 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14214 n6232 p_4_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14213 c_4_17_s2_s c_4_17_cin n6231 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14212 vdd c_4_17_s1_s n6222 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14211 c_4_17_s1_s c_4_17_a n6229 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14210 n6229 p_4_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14209 n5919 p_4_2_d2j n6234 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14208 n6234 p_4_2_d2jbar n5918 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14207 n5918 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14206 vdd a_16 n5919 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14205 vdd p_4_17_t_s n6227 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14204 n6227 p_4_1_n2j p_4_17_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14203 vdd n6234 n6235 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14202 n6235 n6239 p_4_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14201 n6239 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14200 vdd n6585 n6236 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14199 n6228 p_4_1_n2j p_4_16_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14198 vdd p_4_16_t_s n6228 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14197 vdd a_14 n6240 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14196 n6241 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14195 n6389 p_4_2_d2j n6241 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14194 n6240 p_4_2_d2jbar n6389 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14193 n6585 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14192 n6236 n6389 p_4_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14191 n6226 c_4_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14190 c_4_16_s1_s p_4_16_pi2j n6226 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14189 vdd c_4_16_s1_s n6386 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14188 c_4_16_s2_s c_3_17_cout n6385 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14187 n6225 c_4_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14186 n6580 p_4_16_pi2j n6225 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14185 n6580 c_3_17_cout n6383 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14184 vdd c_4_16_a n6383 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14183 n6383 p_4_16_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14182 c_5_15_cin n6580 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14181 n6385 n6386 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14180 c_5_14_a c_4_16_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14179 c_5_13_a c_4_15_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14178 n6749 n6750 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14177 c_4_15_cout n7003 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14176 n6995 c_4_15_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14175 vdd c_4_15_b n6995 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14174 n7003 c_4_15_cin n6995 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14173 n7003 c_4_15_a n7004 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14172 n7004 c_4_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14171 c_4_15_s2_s c_4_15_cin n6749 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14170 vdd c_4_15_s1_s n6750 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14169 c_4_15_s1_s c_4_15_a n7001 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14168 n7001 c_4_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14167 n6754 p_4_2_d2j n6752 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14166 n6752 p_4_2_d2jbar n6753 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14165 n6753 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14164 vdd a_14 n6754 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14163 vdd p_4_15_t_s n6748 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14162 n6748 p_4_1_n2j c_4_15_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14161 vdd n6752 n6751 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14160 n6751 n7007 p_4_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14159 n7007 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14158 vdd n7187 n7006 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14157 n7002 p_4_1_n2j p_4_14_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14156 vdd p_4_14_t_s n7002 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14155 vdd a_12 n7008 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14154 n7009 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14153 n7190 p_4_2_d2j n7009 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14152 n7008 p_4_2_d2jbar n7190 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14151 n7187 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14150 n7006 n7190 p_4_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14149 n6999 c_4_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14148 c_4_14_s1_s p_4_14_pi2j n6999 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14147 vdd c_4_14_s1_s n7184 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14146 c_4_14_s2_s c_3_15_cout n7183 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14145 n6998 c_4_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14144 n7181 p_4_14_pi2j n6998 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14143 n7181 c_3_15_cout n6994 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14142 vdd c_4_14_a n6994 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14141 n6994 p_4_14_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14140 c_5_13_cin n7181 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14139 n7183 n7184 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14138 c_5_12_a c_4_14_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14137 c_5_11_a c_4_13_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14136 n7555 n7558 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14135 c_4_13_cout n7556 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14134 n7766 c_4_13_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14133 vdd c_4_13_b n7766 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14132 n7556 c_4_13_cin n7766 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14131 n7556 c_4_13_a n7772 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14130 n7772 c_4_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14129 c_4_13_s2_s c_4_13_cin n7555 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14128 vdd c_4_13_s1_s n7558 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14127 c_4_13_s1_s c_4_13_a n7773 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14126 n7773 c_4_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14125 n7562 p_4_2_d2j n7560 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14124 n7560 p_4_2_d2jbar n7561 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14123 n7561 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14122 vdd a_12 n7562 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14121 vdd p_4_13_t_s n7554 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14120 n7554 p_4_1_n2j c_4_13_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14119 vdd n7560 n7559 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14118 n7559 n7563 p_4_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14117 n7563 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14116 vdd n7987 n7775 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14115 n7770 p_4_1_n2j c_4_12_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14114 vdd p_4_12_t_s n7770 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14113 vdd a_10 n7776 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14112 n7777 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14111 n7990 p_4_2_d2j n7777 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14110 n7776 p_4_2_d2jbar n7990 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14109 n7987 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14108 n7775 n7990 p_4_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14107 n7771 c_4_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14106 c_4_12_s1_s c_4_12_b n7771 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14105 vdd c_4_12_s1_s n7983 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14104 c_4_12_s2_s c_3_13_cout n7769 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14103 n7768 c_4_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14102 n7978 c_4_12_b n7768 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14101 n7978 c_3_13_cout n7765 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14100 vdd c_4_12_a n7765 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14099 n7765 c_4_12_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14098 c_5_11_cin n7978 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14097 n7769 n7983 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14096 c_5_10_a c_4_12_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14095 c_5_9_a c_4_11_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14094 n8359 n8355 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14093 c_4_11_cout n8360 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14092 n8351 c_4_11_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14091 vdd p_4_11_pi2j n8351 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14090 n8360 c_4_11_cin n8351 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14089 n8360 c_4_11_a n8358 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14088 n8358 p_4_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14087 c_4_11_s2_s c_4_11_cin n8359 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14086 vdd c_4_11_s1_s n8355 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14085 c_4_11_s1_s c_4_11_a n8356 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14084 n8356 p_4_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14083 n8366 p_4_2_d2j n8364 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14082 n8364 p_4_2_d2jbar n8365 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14081 n8365 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14080 vdd a_10 n8366 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14079 vdd p_4_11_t_s n8354 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14078 n8354 p_4_1_n2j p_4_11_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14077 vdd n8364 n8361 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14076 n8361 n8367 p_4_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14075 n8367 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14074 vdd n8741 n8521 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14073 n8520 p_4_1_n2j p_4_10_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14072 vdd p_4_10_t_s n8520 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14071 vdd a_8 n8522 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14070 n8523 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14069 n8744 p_4_2_d2j n8523 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14068 n8522 p_4_2_d2jbar n8744 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14067 n8741 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14066 n8521 n8744 p_4_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14065 n8519 c_4_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14064 c_4_10_s1_s p_4_10_pi2j n8519 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14063 vdd c_4_10_s1_s n8738 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14062 c_4_10_s2_s c_3_11_cout n8517 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14061 n8518 c_4_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14060 n8731 p_4_10_pi2j n8518 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14059 n8731 c_3_11_cout n8516 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14058 vdd c_4_10_a n8516 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14057 n8516 p_4_10_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14056 c_5_9_cin n8731 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14055 n8517 n8738 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14054 c_5_8_a c_4_10_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14053 c_5_7_a c_4_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14052 n9123 n9119 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14051 c_4_9_cout n9124 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14050 n9113 c_4_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14049 vdd p_4_9_pi2j n9113 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14048 n9124 c_4_9_cin n9113 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14047 n9124 c_4_9_a n9122 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14046 n9122 p_4_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14045 c_4_9_s2_s c_4_9_cin n9123 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14044 vdd c_4_9_s1_s n9119 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14043 c_4_9_s1_s c_4_9_a n9120 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14042 n9120 p_4_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14041 n9130 p_4_2_d2j n9129 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14040 n9129 p_4_2_d2jbar n9128 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14039 n9128 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14038 vdd a_8 n9130 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14037 vdd p_4_9_t_s n9118 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14036 n9118 p_4_1_n2j p_4_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14035 vdd n9129 n9125 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14034 n9125 n9131 p_4_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14033 n9131 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14032 vdd n9486 n9260 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14031 n9259 p_4_1_n2j p_4_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14030 vdd p_4_8_t_s n9259 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14029 vdd a_6 n9261 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14028 n9262 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_14027 n9488 p_4_2_d2j n9262 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14026 n9261 p_4_2_d2jbar n9488 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_14025 n9486 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14024 n9260 n9488 p_4_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_14023 n9117 c_4_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14022 c_4_8_s1_s p_4_8_pi2j n9117 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14021 vdd c_4_8_s1_s n9474 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14020 c_4_8_s2_s c_3_9_cout n9258 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_14019 n9116 c_4_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14018 n9479 p_4_8_pi2j n9116 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14017 n9479 c_3_9_cout n9257 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14016 vdd c_4_8_a n9257 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14015 n9257 p_4_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14014 c_5_7_cin n9479 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14013 n9258 n9474 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14012 c_5_6_a c_4_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14011 c_5_5_a c_4_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14010 n9915 n9912 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14009 c_4_7_cout n9917 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_14008 n9905 c_4_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_14007 vdd p_4_7_pi2j n9905 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14006 n9917 c_4_7_cin n9905 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14005 n9917 c_4_7_a n9914 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14004 n9914 p_4_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14003 c_4_7_s2_s c_4_7_cin n9915 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14002 vdd c_4_7_s1_s n9912 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_14001 c_4_7_s1_s c_4_7_a n9913 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_14000 n9913 p_4_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13999 n9597 p_4_2_d2j n9918 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13998 n9918 p_4_2_d2jbar n9596 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13997 n9596 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13996 vdd a_6 n9597 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13995 vdd p_4_7_t_s n9910 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13994 n9910 p_4_1_n2j p_4_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13993 vdd n9918 n9919 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13992 n9919 n9923 p_4_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13991 n9923 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13990 vdd n10259 n9920 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13989 n9911 p_4_1_n2j p_4_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13988 vdd p_4_6_t_s n9911 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13987 vdd a_4 n9924 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13986 n9925 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13985 n10257 p_4_2_d2j n9925 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13984 n9924 p_4_2_d2jbar n10257 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13983 n10259 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13982 n9920 n10257 p_4_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13981 n9909 c_4_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13980 c_4_6_s1_s p_4_6_pi2j n9909 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13979 vdd c_4_6_s1_s n10047 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13978 c_4_6_s2_s c_3_7_cout n10046 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13977 n9908 c_4_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13976 n10252 p_4_6_pi2j n9908 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13975 n10252 c_3_7_cout n10045 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13974 vdd c_4_6_a n10045 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13973 n10045 p_4_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13972 c_5_5_cin n10252 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13971 n10046 n10047 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13970 c_5_4_a c_4_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13969 c_5_3_a c_4_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13968 n10424 n10425 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13967 c_4_5_cout n10682 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13966 n10673 c_4_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13965 vdd c_4_5_b n10673 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13964 n10682 c_4_5_cin n10673 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13963 n10682 c_4_5_a n10681 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13962 n10681 c_4_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13961 c_4_5_s2_s c_4_5_cin n10424 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13960 vdd c_4_5_s1_s n10425 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13959 c_4_5_s1_s c_4_5_a n10680 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13958 n10680 c_4_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13957 n10428 p_4_2_d2j n10683 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13956 n10683 p_4_2_d2jbar n10427 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13955 n10427 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13954 vdd a_4 n10428 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13953 vdd p_4_5_t_s n10423 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13952 n10423 p_4_1_n2j c_4_5_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13951 vdd n10683 n10426 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13950 n10426 n10686 p_4_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13949 n10686 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13948 vdd n10861 n10685 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13947 n10677 p_4_1_n2j p_4_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13946 vdd p_4_4_t_s n10677 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13945 vdd a_2 n10687 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13944 n10688 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13943 n10864 p_4_2_d2j n10688 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13942 n10687 p_4_2_d2jbar n10864 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13941 n10861 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13940 n10685 n10864 p_4_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13939 n10678 c_4_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13938 c_4_4_s1_s p_4_4_pi2j n10678 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13937 vdd c_4_4_s1_s n10860 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13936 c_4_4_s2_s c_3_5_cout n10857 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13935 n10676 c_4_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13934 n10855 p_4_4_pi2j n10676 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13933 n10855 c_3_5_cout n10672 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13932 vdd c_4_4_a n10672 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13931 n10672 p_4_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13930 c_5_3_cin n10855 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13929 n10857 n10860 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13928 c_5_2_a c_4_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13927 c_5_1_a c_4_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13926 n11220 n11223 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13925 c_4_3_cout n11221 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13924 n11431 c_4_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13923 vdd c_4_3_b n11431 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13922 n11221 c_4_3_cin n11431 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13921 n11221 c_4_3_a n11437 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13920 n11437 c_4_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13919 c_4_3_s2_s c_4_3_cin n11220 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13918 vdd c_4_3_s1_s n11223 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13917 c_4_3_s1_s c_4_3_a n11438 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13916 n11438 c_4_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13915 n11227 p_4_2_d2j n11225 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13914 n11225 p_4_2_d2jbar n11226 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13913 n11226 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13912 vdd a_2 n11227 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13911 vdd p_4_3_t_s n11219 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13910 n11219 p_4_1_n2j c_4_3_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13909 vdd n11225 n11224 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13908 n11224 n11228 p_4_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13907 n11228 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13906 vdd n11650 n11440 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13905 n11435 p_4_1_n2j c_4_2_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13904 vdd p_4_2_t_s n11435 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13903 vdd a_0 n11441 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13902 n11442 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13901 n11653 p_4_2_d2j n11442 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13900 n11441 p_4_2_d2jbar n11653 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13899 n11650 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13898 n11440 n11653 p_4_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13897 n11436 c_4_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13896 c_4_2_s1_s c_4_2_b n11436 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13895 vdd c_4_2_s1_s n11646 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13894 c_4_2_s2_s c_3_3_cout n11434 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13893 n11433 c_4_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13892 n11643 c_4_2_b n11433 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13891 n11643 c_3_3_cout n11430 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13890 vdd c_4_2_a n11430 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13889 n11430 c_4_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13888 c_5_1_cin n11643 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13887 n11434 n11646 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13886 c_4_2_sum c_4_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13885 c_4_1_sum c_4_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13884 n12026 n12024 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13883 c_4_1_cout n12025 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13882 n12018 c_4_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13881 vdd p_4_1_pi2j n12018 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13880 n12025 c_4_1_cin n12018 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13879 n12025 c_4_1_a n12027 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13878 n12027 p_4_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13877 c_4_1_s2_s c_4_1_cin n12026 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13876 vdd c_4_1_s1_s n12024 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13875 c_4_1_s1_s c_4_1_a n12021 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13874 n12021 p_4_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13873 n12035 p_4_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13872 vdd a_0 n12035 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13871 vdd p_4_1_t_s n12022 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13870 n12022 p_4_1_n2j p_4_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13869 vdd n12035 n12029 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13868 n12029 n12034 p_4_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13867 n12034 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13866 n12149 c_3_1_sum cl4_4_s1_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13865 vdd n12392 n12149 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13864 p_4 cl4_4_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13863 n12381 c_3_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13862 vdd n12392 n12381 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13861 n12380 n12381 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13860 n12377 c_3_1_cout n12147 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13859 n12147 c_3_2_sum n12377 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13858 n12148 c_3_2_sum n12147 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_13857 vdd c_3_1_cout n12148 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_13856 n12147 c_3_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13855 vdd n12392 n12147 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13854 n12375 n12377 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13853 n12146 c_3_2_sum cl4_4_s2_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13852 vdd c_3_1_cout n12146 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13851 n12372 cl4_4_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_13850 n12145 n12380 cl4_4_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13849 vdd n12372 n12145 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13848 p_5 cl4_4_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13847 n237 p_3_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13846 c_3_33_s1_s c_3_31_a n237 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13845 vdd c_3_33_s1_s n238 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13844 c_3_33_s2_s c_3_32_cin n231 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13843 n232 p_3_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13842 n230 c_3_31_a n232 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13841 n230 c_3_32_cin n234 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13840 vdd p_3_33_pi2j n234 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13839 n234 c_3_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13838 c_4_32_cin n230 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13837 n231 n238 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13836 c_4_31_a c_3_33_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13835 n243 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13834 vdd p_3_33_t_s n236 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13833 n236 p_3_1_n2j p_3_33_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13832 vdd n243 n242 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13831 n242 n240 p_3_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13830 n240 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13829 vdd n578 n375 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13828 n374 p_3_1_n2j p_3_32_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13827 vdd p_3_32_t_s n374 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13826 vdd a_30 n376 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13825 n377 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13824 n580 p_3_2_d2j n377 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13823 n376 p_3_2_d2jbar n580 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13822 n578 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13821 n375 n580 p_3_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13820 n373 c_3_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13819 c_3_32_s1_s p_3_32_pi2j n373 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13818 vdd c_3_32_s1_s n574 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13817 c_3_32_s2_s c_3_32_cin n372 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13816 n370 c_3_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13815 n569 p_3_32_pi2j n370 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13814 n569 c_3_32_cin n371 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13813 vdd c_3_31_a n371 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13812 n371 p_3_32_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13811 c_4_31_cin n569 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13810 n372 n574 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13809 c_4_30_a c_3_32_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13808 c_4_29_a c_3_31_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13807 n935 n944 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13806 c_3_31_cout n936 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13805 n938 c_3_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13804 vdd p_3_31_pi2j n938 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13803 n936 c_3_31_cin n938 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13802 n936 c_3_31_a n934 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13801 n934 p_3_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13800 c_3_31_s2_s c_3_31_cin n935 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13799 vdd c_3_31_s1_s n944 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13798 c_3_31_s1_s c_3_31_a n941 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13797 n941 p_3_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13796 n950 p_3_2_d2j n948 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13795 n948 p_3_2_d2jbar n949 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13794 n949 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13793 vdd a_30 n950 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13792 vdd p_3_31_t_s n940 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13791 n940 p_3_1_n2j p_3_31_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13790 vdd n948 n947 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13789 n947 n945 p_3_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13788 n945 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13787 vdd n1343 n1097 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13786 n1096 p_3_1_n2j p_3_30_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13785 vdd p_3_30_t_s n1096 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13784 vdd a_28 n1098 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13783 n1099 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13782 n1346 p_3_2_d2j n1099 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13781 n1098 p_3_2_d2jbar n1346 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13780 n1343 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13779 n1097 n1346 p_3_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13778 n1095 c_3_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13777 c_3_30_s1_s p_3_30_pi2j n1095 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13776 vdd c_3_30_s1_s n1338 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13775 c_3_30_s2_s c_2_31_cout n1092 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13774 n1093 c_3_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13773 n1333 p_3_30_pi2j n1093 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13772 n1333 c_2_31_cout n1094 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13771 vdd c_3_30_a n1094 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13770 n1094 p_3_30_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13769 c_4_29_cin n1333 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13768 n1092 n1338 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13767 c_4_28_a c_3_30_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13766 c_4_27_a c_3_29_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13765 n1720 n1728 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13764 c_3_29_cout n1721 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13763 n1723 c_3_29_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13762 vdd p_3_29_pi2j n1723 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13761 n1721 c_3_29_cin n1723 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13760 n1721 c_3_29_a n1719 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13759 n1719 p_3_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13758 c_3_29_s2_s c_3_29_cin n1720 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13757 vdd c_3_29_s1_s n1728 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13756 c_3_29_s1_s c_3_29_a n1729 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13755 n1729 p_3_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13754 n1736 p_3_2_d2j n1734 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13753 n1734 p_3_2_d2jbar n1735 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13752 n1735 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13751 vdd a_28 n1736 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13750 vdd p_3_29_t_s n1726 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13749 n1726 p_3_1_n2j p_3_29_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13748 vdd n1734 n1733 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13747 n1733 n1731 p_3_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13746 n1731 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13745 vdd n2093 n1867 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13744 n1865 p_3_1_n2j p_3_28_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13743 vdd p_3_28_t_s n1865 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13742 vdd a_26 n1868 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13741 n1869 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13740 n2095 p_3_2_d2j n1869 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13739 n1868 p_3_2_d2jbar n2095 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13738 n2093 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13737 n1867 n2095 p_3_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13736 n1725 c_3_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13735 c_3_28_s1_s p_3_28_pi2j n1725 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13734 vdd c_3_28_s1_s n1866 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13733 c_3_28_s2_s c_2_29_cout n1863 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13732 n1718 c_3_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13731 n2085 p_3_28_pi2j n1718 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13730 n2085 c_2_29_cout n1864 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13729 vdd c_3_28_a n1864 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13728 n1864 p_3_28_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13727 c_4_27_cin n2085 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13726 n1863 n1866 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13725 c_4_26_a c_3_28_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13724 c_4_25_a c_3_27_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13723 n2226 n2531 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13722 c_3_27_cout n2534 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13721 n2535 c_3_27_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13720 vdd c_3_27_b n2535 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13719 n2534 c_3_27_cin n2535 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13718 n2534 c_3_27_a n2533 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13717 n2533 c_3_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13716 c_3_27_s2_s c_3_27_cin n2226 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13715 vdd c_3_27_s1_s n2531 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13714 c_3_27_s1_s c_3_27_a n2540 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13713 n2540 c_3_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13712 n2229 p_3_2_d2j n2542 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13711 n2542 p_3_2_d2jbar n2228 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13710 n2228 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13709 vdd a_26 n2229 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13708 vdd p_3_27_t_s n2227 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13707 n2227 p_3_1_n2j c_3_27_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13706 vdd n2542 n2545 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13705 n2545 n2543 p_3_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13704 n2543 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13703 vdd n2696 n2546 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13702 n2541 p_3_1_n2j p_3_26_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13701 vdd p_3_26_t_s n2541 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13700 vdd a_24 n2547 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13699 n2548 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13698 n2698 p_3_2_d2j n2548 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13697 n2547 p_3_2_d2jbar n2698 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13696 n2696 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13695 n2546 n2698 p_3_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13694 n2538 c_3_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13693 c_3_26_s1_s p_3_26_pi2j n2538 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13692 vdd c_3_26_s1_s n2695 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13691 c_3_26_s2_s c_2_27_cout n2693 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13690 n2532 c_3_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13689 n2892 p_3_26_pi2j n2532 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13688 n2892 c_2_27_cout n2692 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13687 vdd c_3_26_a n2692 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13686 n2692 p_3_26_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13685 c_4_25_cin n2892 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13684 n2693 n2695 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13683 c_4_24_a c_3_26_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13682 c_4_23_a c_3_25_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13681 n3054 n3058 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13680 c_3_25_cout n3310 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13679 n3312 c_3_25_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13678 vdd c_3_25_b n3312 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13677 n3310 c_3_25_cin n3312 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13676 n3310 c_3_25_a n3311 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13675 n3311 c_3_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13674 c_3_25_s2_s c_3_25_cin n3054 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13673 vdd c_3_25_s1_s n3058 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13672 c_3_25_s1_s c_3_25_a n3317 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13671 n3317 c_3_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13670 n3062 p_3_2_d2j n3060 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13669 n3060 p_3_2_d2jbar n3061 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13668 n3061 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13667 vdd a_24 n3062 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13666 vdd p_3_25_t_s n3057 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13665 n3057 p_3_1_n2j c_3_25_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13664 vdd n3060 n3059 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13663 n3059 n3320 p_3_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13662 n3320 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13661 vdd n3503 n3321 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13660 n3318 p_3_1_n2j c_3_24_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13659 vdd p_3_24_t_s n3318 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13658 vdd a_22 n3322 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13657 n3323 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13656 n3505 p_3_2_d2j n3323 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13655 n3322 p_3_2_d2jbar n3505 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13654 n3503 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13653 n3321 n3505 p_3_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13652 n3315 c_3_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13651 c_3_24_s1_s c_3_24_b n3315 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13650 vdd c_3_24_s1_s n3500 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13649 c_3_24_s2_s c_2_25_cout n3497 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13648 n3309 c_3_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13647 n3496 c_3_24_b n3309 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13646 n3496 c_2_25_cout n3308 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13645 vdd c_3_24_a n3308 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13644 n3308 c_3_24_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13643 c_4_23_cin n3496 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13642 n3497 n3500 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13641 c_4_22_a c_3_24_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13640 c_4_21_a c_3_23_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13639 n3900 n3908 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13638 c_3_23_cout n3901 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13637 n4082 c_3_23_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13636 vdd c_3_23_b n4082 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13635 n3901 c_3_23_cin n4082 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13634 n3901 c_3_23_a n3899 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13633 n3899 c_3_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13632 c_3_23_s2_s c_3_23_cin n3900 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13631 vdd c_3_23_s1_s n3908 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13630 c_3_23_s1_s c_3_23_a n3905 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13629 n3905 c_3_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13628 n3914 p_3_2_d2j n3912 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13627 n3912 p_3_2_d2jbar n3913 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13626 n3913 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13625 vdd a_22 n3914 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13624 vdd p_3_23_t_s n3906 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13623 n3906 p_3_1_n2j c_3_23_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13622 vdd n3912 n3911 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13621 n3911 n3909 p_3_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13620 n3909 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13619 vdd n4320 n4086 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13618 n4085 p_3_1_n2j p_3_22_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13617 vdd p_3_22_t_s n4085 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13616 vdd a_20 n4087 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13615 n4088 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13614 n4322 p_3_2_d2j n4088 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13613 n4087 p_3_2_d2jbar n4322 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13612 n4320 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13611 n4086 n4322 p_3_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13610 n4084 c_3_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13609 c_3_22_s1_s p_3_22_pi2j n4084 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13608 vdd c_3_22_s1_s n4315 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13607 c_3_22_s2_s c_2_23_cout n4081 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13606 n4079 c_3_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13605 n4310 p_3_22_pi2j n4079 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13604 n4310 c_2_23_cout n4080 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13603 vdd c_3_22_a n4080 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13602 n4080 p_3_22_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13601 c_4_21_cin n4310 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13600 n4081 n4315 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13599 c_4_20_a c_3_22_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13598 c_4_19_a c_3_21_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13597 n4682 n4688 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13596 c_3_21_cout n4683 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13595 n4685 c_3_21_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13594 vdd p_3_21_pi2j n4685 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13593 n4683 c_3_21_cin n4685 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13592 n4683 c_3_21_a n4681 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13591 n4681 p_3_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13590 c_3_21_s2_s c_3_21_cin n4682 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13589 vdd c_3_21_s1_s n4688 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13588 c_3_21_s1_s c_3_21_a n4689 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13587 n4689 p_3_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13586 n4697 p_3_2_d2j n4695 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13585 n4695 p_3_2_d2jbar n4696 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13584 n4696 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13583 vdd a_20 n4697 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13582 vdd p_3_21_t_s n4687 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13581 n4687 p_3_1_n2j p_3_21_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13580 vdd n4695 n4694 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13579 n4694 n4692 p_3_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13578 n4692 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13577 vdd n5066 n4840 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13576 n4839 p_3_1_n2j p_3_20_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13575 vdd p_3_20_t_s n4839 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13574 vdd a_18 n4841 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13573 n4842 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13572 n5068 p_3_2_d2j n4842 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13571 n4841 p_3_2_d2jbar n5068 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13570 n5066 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13569 n4840 n5068 p_3_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13568 n4838 c_3_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13567 c_3_20_s1_s p_3_20_pi2j n4838 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13566 vdd c_3_20_s1_s n5061 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13565 c_3_20_s2_s c_2_21_cout n4835 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13564 n4836 c_3_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13563 n5058 p_3_20_pi2j n4836 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13562 n5058 c_2_21_cout n4837 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13561 vdd c_3_20_a n4837 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13560 n4837 p_3_20_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13559 c_4_19_cin n5058 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13558 n4835 n5061 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13557 c_4_18_a c_3_20_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13556 c_4_17_a c_3_19_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13555 n5446 n5455 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13554 c_3_19_cout n5448 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13553 n5450 c_3_19_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13552 vdd p_3_19_pi2j n5450 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13551 n5448 c_3_19_cin n5450 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13550 n5448 c_3_19_a n5447 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13549 n5447 p_3_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13548 c_3_19_s2_s c_3_19_cin n5446 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13547 vdd c_3_19_s1_s n5455 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13546 c_3_19_s1_s c_3_19_a n5456 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13545 n5456 p_3_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13544 n5463 p_3_2_d2j n5461 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13543 n5461 p_3_2_d2jbar n5462 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13542 n5462 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13541 vdd a_18 n5463 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13540 vdd p_3_19_t_s n5454 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13539 n5454 p_3_1_n2j p_3_19_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13538 vdd n5461 n5460 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13537 n5460 n5458 p_3_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13536 n5458 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13535 vdd n5820 n5593 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13534 n5591 p_3_1_n2j p_3_18_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13533 vdd p_3_18_t_s n5591 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13532 vdd a_16 n5594 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13531 n5595 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13530 n5822 p_3_2_d2j n5595 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13529 n5594 p_3_2_d2jbar n5822 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13528 n5820 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13527 n5593 n5822 p_3_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13526 n5452 c_3_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13525 c_3_18_s1_s p_3_18_pi2j n5452 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13524 vdd c_3_18_s1_s n5592 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13523 c_3_18_s2_s c_2_19_cout n5590 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13522 n5445 c_3_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13521 n5812 p_3_18_pi2j n5445 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13520 n5812 c_2_19_cout n5589 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13519 vdd c_3_18_a n5589 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13518 n5589 p_3_18_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13517 c_4_17_cin n5812 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13516 n5590 n5592 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13515 c_4_16_a c_3_18_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13514 c_4_15_a c_3_17_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13513 n6245 n6243 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13512 c_3_17_cout n6247 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13511 n6249 c_3_17_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13510 vdd p_3_17_pi2j n6249 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13509 n6247 c_3_17_cin n6249 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13508 n6247 c_3_17_a n6246 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13507 n6246 p_3_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13506 c_3_17_s2_s c_3_17_cin n6245 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13505 vdd c_3_17_s1_s n6243 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13504 c_3_17_s1_s c_3_17_a n6255 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13503 n6255 p_3_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13502 n5924 p_3_2_d2j n6257 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13501 n6257 p_3_2_d2jbar n5923 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13500 n5923 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13499 vdd a_16 n5924 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13498 vdd p_3_17_t_s n6252 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13497 n6252 p_3_1_n2j p_3_17_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13496 vdd n6257 n6260 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13495 n6260 n6258 p_3_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13494 n6258 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13493 vdd n6597 n6261 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13492 n6253 p_3_1_n2j p_3_16_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13491 vdd p_3_16_t_s n6253 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13490 vdd a_14 n6262 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13489 n6263 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13488 n6395 p_3_2_d2j n6263 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13487 n6262 p_3_2_d2jbar n6395 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13486 n6597 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13485 n6261 n6395 p_3_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13484 n6251 c_3_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13483 c_3_16_s1_s p_3_16_pi2j n6251 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13482 vdd c_3_16_s1_s n6393 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13481 c_3_16_s2_s c_2_17_cout n6391 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13480 n6244 c_3_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13479 n6592 p_3_16_pi2j n6244 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13478 n6592 c_2_17_cout n6390 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13477 vdd c_3_16_a n6390 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13476 n6390 p_3_16_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13475 c_4_15_cin n6592 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13474 n6391 n6393 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13473 c_4_14_a c_3_16_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13472 c_4_13_a c_3_15_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13471 n6755 n6759 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13470 c_3_15_cout n7012 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13469 n7013 c_3_15_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13468 vdd c_3_15_b n7013 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13467 n7012 c_3_15_cin n7013 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13466 n7012 c_3_15_a n7014 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13465 n7014 c_3_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13464 c_3_15_s2_s c_3_15_cin n6755 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13463 vdd c_3_15_s1_s n6759 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13462 c_3_15_s1_s c_3_15_a n7019 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13461 n7019 c_3_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13460 n6763 p_3_2_d2j n6761 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13459 n6761 p_3_2_d2jbar n6762 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13458 n6762 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13457 vdd a_14 n6763 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13456 vdd p_3_15_t_s n6758 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13455 n6758 p_3_1_n2j c_3_15_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13454 vdd n6761 n6760 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13453 n6760 n7021 p_3_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13452 n7021 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13451 vdd n7197 n7023 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13450 n7020 p_3_1_n2j p_3_14_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13449 vdd p_3_14_t_s n7020 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13448 vdd a_12 n7024 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13447 n7025 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13446 n7199 p_3_2_d2j n7025 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13445 n7024 p_3_2_d2jbar n7199 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13444 n7197 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13443 n7023 n7199 p_3_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13442 n7017 c_3_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13441 c_3_14_s1_s p_3_14_pi2j n7017 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13440 vdd c_3_14_s1_s n7194 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13439 c_3_14_s2_s c_2_15_cout n7192 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13438 n7011 c_3_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13437 n7191 p_3_14_pi2j n7011 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13436 n7191 c_2_15_cout n7010 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13435 vdd c_3_14_a n7010 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13434 n7010 p_3_14_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13433 c_4_13_cin n7191 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13432 n7192 n7194 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13431 c_4_12_a c_3_14_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13430 c_4_11_a c_3_13_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13429 n7564 n7571 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13428 c_3_13_cout n7565 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13427 n7781 c_3_13_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13426 vdd c_3_13_b n7781 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13425 n7565 c_3_13_cin n7781 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13424 n7565 c_3_13_a n7782 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13423 n7782 c_3_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13422 c_3_13_s2_s c_3_13_cin n7564 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13421 vdd c_3_13_s1_s n7571 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13420 c_3_13_s1_s c_3_13_a n7785 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13419 n7785 c_3_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13418 n7576 p_3_2_d2j n7574 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13417 n7574 p_3_2_d2jbar n7575 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13416 n7575 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13415 vdd a_12 n7576 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13414 vdd p_3_13_t_s n7569 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13413 n7569 p_3_1_n2j c_3_13_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13412 vdd n7574 n7573 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13411 n7573 n7572 p_3_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13410 n7572 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13409 vdd n8000 n7788 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13408 n7786 p_3_1_n2j c_3_12_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13407 vdd p_3_12_t_s n7786 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13406 vdd a_10 n7789 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13405 n7790 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13404 n8002 p_3_2_d2j n7790 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13403 n7789 p_3_2_d2jbar n8002 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13402 n8000 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13401 n7788 n8002 p_3_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13400 n7784 c_3_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13399 c_3_12_s1_s c_3_12_b n7784 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13398 vdd c_3_12_s1_s n7996 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13397 c_3_12_s2_s c_2_13_cout n7780 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13396 n7778 c_3_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13395 n7993 c_3_12_b n7778 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13394 n7993 c_2_13_cout n7779 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13393 vdd c_3_12_a n7779 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13392 n7779 c_3_12_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13391 c_4_11_cin n7993 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13390 n7780 n7996 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13389 c_4_10_a c_3_12_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13388 c_4_9_a c_3_11_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13387 n8370 n8377 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13386 c_3_11_cout n8372 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13385 n8373 c_3_11_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13384 vdd p_3_11_pi2j n8373 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13383 n8372 c_3_11_cin n8373 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13382 n8372 c_3_11_a n8369 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13381 n8369 p_3_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13380 c_3_11_s2_s c_3_11_cin n8370 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13379 vdd c_3_11_s1_s n8377 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13378 c_3_11_s1_s c_3_11_a n8378 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13377 n8378 p_3_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13376 n8385 p_3_2_d2j n8383 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13375 n8383 p_3_2_d2jbar n8384 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13374 n8384 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13373 vdd a_10 n8385 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13372 vdd p_3_11_t_s n8376 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13371 n8376 p_3_1_n2j p_3_11_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13370 vdd n8383 n8382 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13369 n8382 n8380 p_3_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13368 n8380 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13367 vdd n8755 n8529 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13366 n8528 p_3_1_n2j p_3_10_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13365 vdd p_3_10_t_s n8528 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13364 vdd a_8 n8530 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13363 n8531 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13362 n8757 p_3_2_d2j n8531 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13361 n8530 p_3_2_d2jbar n8757 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13360 n8755 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13359 n8529 n8757 p_3_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13358 n8527 c_3_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13357 c_3_10_s1_s p_3_10_pi2j n8527 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13356 vdd c_3_10_s1_s n8750 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13355 c_3_10_s2_s c_2_11_cout n8524 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13354 n8525 c_3_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13353 n8745 p_3_10_pi2j n8525 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13352 n8745 c_2_11_cout n8526 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13351 vdd c_3_10_a n8526 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13350 n8526 p_3_10_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13349 c_4_9_cin n8745 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13348 n8524 n8750 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13347 c_4_8_a c_3_10_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13346 c_4_7_a c_3_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13345 n9135 n9143 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13344 c_3_9_cout n9136 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13343 n9138 c_3_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13342 vdd p_3_9_pi2j n9138 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13341 n9136 c_3_9_cin n9138 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13340 n9136 c_3_9_a n9134 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13339 n9134 p_3_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13338 c_3_9_s2_s c_3_9_cin n9135 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13337 vdd c_3_9_s1_s n9143 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13336 c_3_9_s1_s c_3_9_a n9144 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13335 n9144 p_3_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13334 n9151 p_3_2_d2j n9149 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13333 n9149 p_3_2_d2jbar n9150 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13332 n9150 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13331 vdd a_8 n9151 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13330 vdd p_3_9_t_s n9142 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13329 n9142 p_3_1_n2j p_3_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13328 vdd n9149 n9148 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13327 n9148 n9146 p_3_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13326 n9146 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13325 vdd n9501 n9266 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13324 n9265 p_3_1_n2j p_3_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13323 vdd p_3_8_t_s n9265 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13322 vdd a_6 n9267 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13321 n9268 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13320 n9503 p_3_2_d2j n9268 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13319 n9267 p_3_2_d2jbar n9503 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13318 n9501 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13317 n9266 n9503 p_3_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13316 n9140 c_3_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13315 c_3_8_s1_s p_3_8_pi2j n9140 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13314 vdd c_3_8_s1_s n9493 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13313 c_3_8_s2_s c_2_9_cout n9264 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13312 n9133 c_3_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13311 n9491 p_3_8_pi2j n9133 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13310 n9491 c_2_9_cout n9263 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13309 vdd c_3_8_a n9263 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13308 n9263 p_3_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13307 c_4_7_cin n9491 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13306 n9264 n9493 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13305 c_4_6_a c_3_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13304 c_4_5_a c_3_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13303 n9928 n9939 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13302 c_3_7_cout n9930 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13301 n9932 c_3_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13300 vdd p_3_7_pi2j n9932 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13299 n9930 c_3_7_cin n9932 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13298 n9930 c_3_7_a n9929 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13297 n9929 p_3_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13296 c_3_7_s2_s c_3_7_cin n9928 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13295 vdd c_3_7_s1_s n9939 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13294 c_3_7_s1_s c_3_7_a n9940 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13293 n9940 p_3_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13292 n9602 p_3_2_d2j n9941 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13291 n9941 p_3_2_d2jbar n9601 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13290 n9601 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13289 vdd a_6 n9602 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13288 vdd p_3_7_t_s n9937 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13287 n9937 p_3_1_n2j p_3_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13286 vdd n9941 n9944 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13285 n9944 n9942 p_3_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13284 n9942 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13283 vdd n10272 n9945 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13282 n9935 p_3_1_n2j p_3_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13281 vdd p_3_6_t_s n9935 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13280 vdd a_4 n9946 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13279 n9947 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13278 n10271 p_3_2_d2j n9947 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13277 n9946 p_3_2_d2jbar n10271 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13276 n10272 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13275 n9945 n10271 p_3_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13274 n9934 c_3_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13273 c_3_6_s1_s p_3_6_pi2j n9934 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13272 vdd c_3_6_s1_s n10052 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13271 c_3_6_s2_s c_2_7_cout n10050 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13270 n9927 c_3_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13269 n10265 p_3_6_pi2j n9927 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13268 n10265 c_2_7_cout n10051 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13267 vdd c_3_6_a n10051 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13266 n10051 p_3_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13265 c_4_5_cin n10265 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13264 n10050 n10052 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13263 c_4_4_a c_3_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13262 c_4_3_a c_3_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13261 n10430 n10434 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13260 c_3_5_cout n10692 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13259 n10693 c_3_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13258 vdd c_3_5_b n10693 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13257 n10692 c_3_5_cin n10693 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13256 n10692 c_3_5_a n10691 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13255 n10691 c_3_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13254 c_3_5_s2_s c_3_5_cin n10430 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13253 vdd c_3_5_s1_s n10434 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13252 c_3_5_s1_s c_3_5_a n10698 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13251 n10698 c_3_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13250 n10437 p_3_2_d2j n10702 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13249 n10702 p_3_2_d2jbar n10436 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13248 n10436 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13247 vdd a_4 n10437 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13246 vdd p_3_5_t_s n10433 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13245 n10433 p_3_1_n2j c_3_5_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13244 vdd n10702 n10435 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13243 n10435 n10701 p_3_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13242 n10701 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13241 vdd n10871 n10703 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13240 n10699 p_3_1_n2j p_3_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13239 vdd p_3_4_t_s n10699 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13238 vdd a_2 n10704 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13237 n10705 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13236 n10873 p_3_2_d2j n10705 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13235 n10704 p_3_2_d2jbar n10873 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13234 n10871 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13233 n10703 n10873 p_3_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13232 n10696 c_3_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13231 c_3_4_s1_s p_3_4_pi2j n10696 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13230 vdd c_3_4_s1_s n10870 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13229 c_3_4_s2_s c_2_5_cout n10866 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13228 n10689 c_3_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13227 n10865 p_3_4_pi2j n10689 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13226 n10865 c_2_5_cout n10690 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13225 vdd c_3_4_a n10690 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13224 n10690 p_3_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13223 c_4_3_cin n10865 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13222 n10866 n10870 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13221 c_4_2_a c_3_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13220 c_4_1_a c_3_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13219 n11229 n11236 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13218 c_3_3_cout n11230 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13217 n11446 c_3_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13216 vdd c_3_3_b n11446 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13215 n11230 c_3_3_cin n11446 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13214 n11230 c_3_3_a n11447 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13213 n11447 c_3_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13212 c_3_3_s2_s c_3_3_cin n11229 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13211 vdd c_3_3_s1_s n11236 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13210 c_3_3_s1_s c_3_3_a n11450 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13209 n11450 c_3_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13208 n11241 p_3_2_d2j n11239 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13207 n11239 p_3_2_d2jbar n11240 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13206 n11240 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13205 vdd a_2 n11241 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13204 vdd p_3_3_t_s n11234 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13203 n11234 p_3_1_n2j c_3_3_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13202 vdd n11239 n11238 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13201 n11238 n11237 p_3_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13200 n11237 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13199 vdd n11663 n11453 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13198 n11451 p_3_1_n2j c_3_2_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13197 vdd p_3_2_t_s n11451 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13196 vdd a_0 n11454 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13195 n11455 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13194 n11665 p_3_2_d2j n11455 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13193 n11454 p_3_2_d2jbar n11665 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13192 n11663 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13191 n11453 n11665 p_3_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13190 n11449 c_3_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13189 c_3_2_s1_s c_3_2_b n11449 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13188 vdd c_3_2_s1_s n11659 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13187 c_3_2_s2_s c_2_3_cout n11445 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13186 n11443 c_3_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13185 n11656 c_3_2_b n11443 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13184 n11656 c_2_3_cout n11444 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13183 vdd c_3_2_a n11444 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13182 n11444 c_3_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13181 c_4_1_cin n11656 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13180 n11445 n11659 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13179 c_3_2_sum c_3_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13178 c_3_1_sum c_3_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13177 n12038 n12046 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13176 c_3_1_cout n12039 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13175 n12041 c_3_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13174 vdd p_3_1_pi2j n12041 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13173 n12039 c_3_1_cin n12041 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13172 n12039 c_3_1_a n12037 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13171 n12037 p_3_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13170 c_3_1_s2_s c_3_1_cin n12038 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13169 vdd c_3_1_s1_s n12046 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13168 c_3_1_s1_s c_3_1_a n12047 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13167 n12047 p_3_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13166 n12054 p_3_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13165 vdd a_0 n12054 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13164 vdd p_3_1_t_s n12044 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13163 n12044 p_3_1_n2j p_3_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13162 vdd n12054 n12051 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13161 n12051 n12050 p_3_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13160 n12050 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13159 n12154 c_2_1_sum cl4_3_s1_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13158 vdd n12406 n12154 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13157 p_2 cl4_3_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13156 n12397 c_2_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13155 vdd n12406 n12397 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13154 n12398 n12397 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13153 n12394 c_2_1_cout n12153 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13152 n12153 c_2_2_sum n12394 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13151 n12152 c_2_2_sum n12153 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_13150 vdd c_2_1_cout n12152 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_13149 n12153 c_2_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13148 vdd n12406 n12153 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13147 n12392 n12394 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13146 n12151 c_2_2_sum cl4_3_s2_s vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13145 vdd c_2_1_cout n12151 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13144 n12390 cl4_3_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_13143 n12150 n12398 cl4_3_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13142 vdd n12390 n12150 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13141 p_3 cl4_3_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13140 c_3_31_a c_2_33_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13139 n245 n251 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13138 c_3_32_cin n248 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13137 n244 c_2_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13136 vdd p_2_33_pi2j n244 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13135 n248 vss n244 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13134 n248 c_2_31_a n246 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13133 n246 p_2_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13132 c_2_33_s2_s vss n245 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13131 vdd c_2_33_s1_s n251 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13130 c_2_33_s1_s c_2_31_a n252 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13129 n252 p_2_33_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13128 n258 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13127 vdd p_2_33_t_s n249 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13126 n249 p_2_1_n2j p_2_33_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13125 vdd n258 n254 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13124 n254 n255 p_2_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13123 n255 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13122 vdd n586 n380 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13121 n379 p_2_1_n2j c_2_32_b vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13120 vdd p_2_32_t_s n379 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13119 vdd a_30 n382 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13118 n381 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13117 n590 p_2_2_d2j n381 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13116 n382 p_2_2_d2jbar n590 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13115 n586 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13114 n380 n590 p_2_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13113 vdd c_2_32_s1_s c_3_30_a vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_13112 n583 c_2_32_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13111 vdd c_2_31_a n583 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13110 c_3_31_cin n583 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13109 c_2_32_s1_s c_2_32_b n378 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13108 n378 c_2_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13107 c_3_29_a c_2_31_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13106 n953 n958 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13105 c_2_31_cout n955 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13104 n951 c_2_31_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13103 vdd p_2_31_pi2j n951 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13102 n955 vss n951 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13101 n955 c_2_31_a n952 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13100 n952 p_2_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13099 c_2_31_s2_s vss n953 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13098 vdd c_2_31_s1_s n958 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13097 c_2_31_s1_s c_2_31_a n960 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13096 n960 p_2_31_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13095 n966 p_2_2_d2j n968 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13094 n968 p_2_2_d2jbar n967 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13093 n967 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13092 vdd a_30 n966 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13091 vdd p_2_31_t_s n957 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13090 n957 p_2_1_n2j p_2_31_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13089 vdd n968 n962 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13088 n962 n963 p_2_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13087 n963 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13086 vdd n1354 n1102 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13085 n1101 p_2_1_n2j p_2_30_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13084 vdd p_2_30_t_s n1101 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13083 vdd a_28 n1104 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13082 n1103 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13081 n1355 p_2_2_d2j n1103 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13080 n1104 p_2_2_d2jbar n1355 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13079 n1354 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13078 n1102 n1355 p_2_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13077 vdd c_2_30_s1_s c_3_28_a vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_13076 n1349 p_2_30_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13075 vdd c_2_30_a n1349 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13074 c_3_29_cin n1349 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13073 c_2_30_s1_s p_2_30_pi2j n1100 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13072 n1100 c_2_30_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13071 c_3_27_a c_2_29_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13070 n1740 n1745 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13069 c_2_29_cout n1739 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13068 n1737 c_2_29_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13067 vdd p_2_29_pi2j n1737 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13066 n1739 p_18_1_c2j n1737 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13065 n1739 c_2_29_a n1738 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13064 n1738 p_2_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13063 c_2_29_s2_s p_18_1_c2j n1740 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13062 vdd c_2_29_s1_s n1745 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13061 c_2_29_s1_s c_2_29_a n1747 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13060 n1747 p_2_29_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13059 n1755 p_2_2_d2j n1754 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13058 n1754 p_2_2_d2jbar n1753 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13057 n1753 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13056 vdd a_28 n1755 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13055 vdd p_2_29_t_s n1744 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13054 n1744 p_2_1_n2j p_2_29_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13053 vdd n1754 n1750 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13052 n1750 n1751 p_2_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13051 n1751 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13050 vdd n2104 n1871 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13049 n1870 p_2_1_n2j p_2_28_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13048 vdd p_2_28_t_s n1870 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13047 vdd a_26 n1872 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13046 n1873 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13045 n2106 p_2_2_d2j n1873 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13044 n1872 p_2_2_d2jbar n2106 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13043 n2104 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13042 n1871 n2106 p_2_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13041 vdd c_2_28_s1_s c_3_26_a vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_13040 n2099 p_2_28_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13039 vdd c_2_28_a n2099 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13038 c_3_27_cin n2099 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13037 c_2_28_s1_s p_2_28_pi2j n1743 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13036 n1743 c_2_28_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13035 c_3_25_a c_2_27_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13034 n2233 n2551 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13033 c_2_27_cout n2552 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13032 n2549 n2555 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13031 vdd c_2_27_b n2549 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13030 n2552 p_17_1_c2j n2549 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13029 n2552 n2555 n2553 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_13028 n2553 c_2_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13027 c_2_27_s2_s p_17_1_c2j n2233 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_13026 vdd c_2_27_s1_s n2551 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_13025 c_2_27_s1_s n2555 n2559 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13024 n2559 c_2_27_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13023 n2236 p_2_2_d2j n2561 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13022 n2561 p_2_2_d2jbar n2237 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13021 n2237 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13020 vdd a_26 n2236 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13019 vdd p_2_27_t_s n2234 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13018 n2234 p_2_1_n2j c_2_27_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13017 vdd n2561 n2563 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13016 n2563 n2560 p_2_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13015 n2560 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13014 vdd n2700 n2564 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13013 n2557 p_2_1_n2j c_2_26_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13012 vdd p_2_26_t_s n2557 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13011 vdd a_24 n2566 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13010 n2565 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_13009 n2701 p_2_2_d2j n2565 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13008 n2566 p_2_2_d2jbar n2701 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_13007 n2700 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13006 n2564 n2701 p_2_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_13005 vdd c_2_26_s1_s c_3_24_a vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_13004 n2905 c_2_26_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13003 vdd c_2_26_a n2905 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13002 c_3_25_cin n2905 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_13001 c_2_26_s1_s c_2_26_b n2556 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_13000 n2556 c_2_26_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12999 c_3_23_a c_2_25_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12998 n3063 n3065 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12997 c_2_25_cout n3325 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12996 n3324 c_2_25_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12995 vdd c_2_25_b n3324 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12994 n3325 p_16_1_c2j n3324 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12993 n3325 c_2_25_a n3326 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12992 n3326 c_2_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12991 c_2_25_s2_s p_16_1_c2j n3063 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12990 vdd c_2_25_s1_s n3065 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12989 c_2_25_s1_s c_2_25_a n3332 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12988 n3332 c_2_25_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12987 n3069 p_2_2_d2j n3071 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12986 n3071 p_2_2_d2jbar n3070 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12985 n3070 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12984 vdd a_24 n3069 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12983 vdd p_2_25_t_s n3066 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12982 n3066 p_2_1_n2j c_2_25_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12981 vdd n3071 n3067 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12980 n3067 n3334 p_2_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12979 n3334 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12978 vdd n3511 n3335 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12977 n3331 p_2_1_n2j c_2_24_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12976 vdd p_2_24_t_s n3331 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12975 vdd a_22 n3337 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12974 n3336 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12973 n3514 p_2_2_d2j n3336 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12972 n3337 p_2_2_d2jbar n3514 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12971 n3511 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12970 n3335 n3514 p_2_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12969 vdd c_2_24_s1_s c_3_22_a vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_12968 n3508 c_2_24_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12967 vdd c_2_24_a n3508 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12966 c_3_23_cin n3508 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12965 c_2_24_s1_s c_2_24_b n3329 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12964 n3329 c_2_24_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12963 c_3_21_a c_2_23_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12962 n3916 n3921 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12961 c_2_23_cout n3917 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12960 n4089 c_2_23_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12959 vdd c_2_23_b n4089 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12958 n3917 p_15_1_c2j n4089 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12957 n3917 c_2_23_a n3915 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12956 n3915 c_2_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12955 c_2_23_s2_s p_15_1_c2j n3916 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12954 vdd c_2_23_s1_s n3921 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12953 c_2_23_s1_s c_2_23_a n3922 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12952 n3922 c_2_23_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12951 n3928 p_2_2_d2j n3930 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12950 n3930 p_2_2_d2jbar n3929 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12949 n3929 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12948 vdd a_22 n3928 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12947 vdd p_2_23_t_s n3920 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12946 n3920 p_2_1_n2j c_2_23_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12945 vdd n3930 n3924 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12944 n3924 n3925 p_2_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12943 n3925 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12942 vdd n4329 n4093 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12941 n4092 p_2_1_n2j c_2_22_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12940 vdd p_2_22_t_s n4092 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12939 vdd a_20 n4095 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12938 n4094 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12937 n4333 p_2_2_d2j n4094 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12936 n4095 p_2_2_d2jbar n4333 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12935 n4329 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12934 n4093 n4333 p_2_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12933 vdd c_2_22_s1_s c_3_20_a vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_12932 n4325 c_2_22_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12931 vdd c_2_22_a n4325 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12930 c_3_21_cin n4325 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12929 c_2_22_s1_s c_2_22_b n4091 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12928 n4091 c_2_22_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12927 c_3_19_a c_2_21_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12926 n4700 n4705 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12925 c_2_21_cout n4702 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12924 n4698 c_2_21_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12923 vdd p_2_21_pi2j n4698 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12922 n4702 p_14_1_c2j n4698 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12921 n4702 c_2_21_a n4699 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12920 n4699 p_2_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12919 c_2_21_s2_s p_14_1_c2j n4700 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12918 vdd c_2_21_s1_s n4705 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12917 c_2_21_s1_s c_2_21_a n4707 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12916 n4707 p_2_21_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12915 n4713 p_2_2_d2j n4715 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12914 n4715 p_2_2_d2jbar n4714 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12913 n4714 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12912 vdd a_20 n4713 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12911 vdd p_2_21_t_s n4704 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12910 n4704 p_2_1_n2j p_2_21_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12909 vdd n4715 n4709 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12908 n4709 n4710 p_2_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12907 n4710 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12906 vdd n5075 n4845 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12905 n4844 p_2_1_n2j p_2_20_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12904 vdd p_2_20_t_s n4844 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12903 vdd a_18 n4847 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12902 n4846 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12901 n5078 p_2_2_d2j n4846 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12900 n4847 p_2_2_d2jbar n5078 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12899 n5075 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12898 n4845 n5078 p_2_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12897 vdd c_2_20_s1_s c_3_18_a vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_12896 n5071 p_2_20_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12895 vdd c_2_20_a n5071 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12894 c_3_19_cin n5071 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12893 c_2_20_s1_s p_2_20_pi2j n4843 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12892 n4843 c_2_20_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12891 c_3_17_a c_2_19_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12890 n5465 n5472 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12889 c_2_19_cout n5467 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12888 n5464 c_2_19_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12887 vdd p_2_19_pi2j n5464 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12886 n5467 p_12_1_c2j n5464 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12885 n5467 c_2_19_a n5466 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12884 n5466 p_2_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12883 c_2_19_s2_s p_12_1_c2j n5465 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12882 vdd c_2_19_s1_s n5472 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12881 c_2_19_s1_s c_2_19_a n5473 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12880 n5473 p_2_19_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12879 n5482 p_2_2_d2j n5481 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12878 n5481 p_2_2_d2jbar n5480 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12877 n5480 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12876 vdd a_18 n5482 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12875 vdd p_2_19_t_s n5471 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12874 n5471 p_2_1_n2j p_2_19_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12873 vdd n5481 n5477 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12872 n5477 n5478 p_2_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12871 n5478 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12870 vdd n5830 n5597 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12869 n5596 p_2_1_n2j p_2_18_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12868 vdd p_2_18_t_s n5596 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12867 vdd a_16 n5599 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12866 n5598 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12865 n5833 p_2_2_d2j n5598 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12864 n5599 p_2_2_d2jbar n5833 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12863 n5830 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12862 n5597 n5833 p_2_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12861 vdd c_2_18_s1_s c_3_16_a vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_12860 n5825 p_2_18_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12859 vdd c_2_18_a n5825 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12858 c_3_17_cin n5825 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12857 c_2_18_s1_s p_2_18_pi2j n5470 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12856 n5470 c_2_18_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12855 c_3_15_a c_2_17_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12854 n6266 n6265 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12853 c_2_17_cout n6268 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12852 n6264 c_2_17_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12851 vdd p_2_17_pi2j n6264 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12850 n6268 p_11_1_c2j n6264 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12849 n6268 c_2_17_a n6267 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12848 n6267 p_2_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12847 c_2_17_s2_s p_11_1_c2j n6266 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12846 vdd c_2_17_s1_s n6265 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12845 c_2_17_s1_s c_2_17_a n6276 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12844 n6276 p_2_17_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12843 n5928 p_2_2_d2j n6278 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12842 n6278 p_2_2_d2jbar n5929 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12841 n5929 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12840 vdd a_16 n5928 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12839 vdd p_2_17_t_s n6274 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12838 n6274 p_2_1_n2j p_2_17_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12837 vdd n6278 n6280 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12836 n6280 n6277 p_2_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12835 n6277 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12834 vdd n6609 n6281 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12833 n6272 p_2_1_n2j p_2_16_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12832 vdd p_2_16_t_s n6272 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12831 vdd a_14 n6283 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12830 n6284 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12829 n6397 p_2_2_d2j n6284 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12828 n6283 p_2_2_d2jbar n6397 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12827 n6609 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12826 n6281 n6397 p_2_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12825 vdd c_2_16_s1_s c_3_14_a vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_12824 n6604 p_2_16_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12823 vdd c_2_16_a n6604 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12822 c_3_15_cin n6604 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12821 c_2_16_s1_s p_2_16_pi2j n6271 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12820 n6271 c_2_16_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12819 c_3_13_a c_2_15_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12818 n6764 n6766 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12817 c_2_15_cout n7028 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12816 n7026 c_2_15_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12815 vdd c_2_15_b n7026 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12814 n7028 p_10_1_c2j n7026 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12813 n7028 c_2_15_a n7027 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12812 n7027 c_2_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12811 c_2_15_s2_s p_10_1_c2j n6764 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12810 vdd c_2_15_s1_s n6766 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12809 c_2_15_s1_s c_2_15_a n7034 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12808 n7034 c_2_15_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12807 n6770 p_2_2_d2j n6772 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12806 n6772 p_2_2_d2jbar n6771 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12805 n6771 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12804 vdd a_14 n6770 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12803 vdd p_2_15_t_s n6767 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12802 n6767 p_2_1_n2j c_2_15_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12801 vdd n6772 n6768 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12800 n6768 n7036 p_2_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12799 n7036 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12798 vdd n7205 n7037 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12797 n7032 p_2_1_n2j p_2_14_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12796 vdd p_2_14_t_s n7032 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12795 vdd a_12 n7039 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12794 n7038 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12793 n7208 p_2_2_d2j n7038 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12792 n7039 p_2_2_d2jbar n7208 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12791 n7205 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12790 n7037 n7208 p_2_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12789 vdd c_2_14_s1_s c_3_12_a vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_12788 n7202 p_2_14_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12787 vdd c_2_14_a n7202 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12786 c_3_13_cin n7202 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12785 c_2_14_s1_s p_2_14_pi2j n7031 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12784 n7031 c_2_14_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12783 c_3_11_a c_2_13_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12782 n7577 n7582 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12781 c_2_13_cout n7578 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12780 n7791 c_2_13_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12779 vdd c_2_13_b n7791 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12778 n7578 p_9_1_c2j n7791 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12777 n7578 c_2_13_a n7792 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12776 n7792 c_2_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12775 c_2_13_s2_s p_9_1_c2j n7577 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12774 vdd c_2_13_s1_s n7582 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12773 c_2_13_s1_s c_2_13_a n7795 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12772 n7795 c_2_13_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12771 n7587 p_2_2_d2j n7589 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12770 n7589 p_2_2_d2jbar n7588 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12769 n7588 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12768 vdd a_12 n7587 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12767 vdd p_2_13_t_s n7581 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12766 n7581 p_2_1_n2j c_2_13_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12765 vdd n7589 n7584 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12764 n7584 n7585 p_2_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12763 n7585 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12762 vdd n8008 n7798 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12761 n7796 p_2_1_n2j c_2_12_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12760 vdd p_2_12_t_s n7796 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12759 vdd a_10 n7800 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12758 n7799 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12757 n8012 p_2_2_d2j n7799 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12756 n7800 p_2_2_d2jbar n8012 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12755 n8008 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12754 n7798 n8012 p_2_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12753 vdd c_2_12_s1_s c_3_10_a vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_12752 n8005 c_2_12_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12751 vdd c_2_12_a n8005 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12750 c_3_11_cin n8005 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12749 c_2_12_s1_s c_2_12_b n7794 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12748 n7794 c_2_12_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12747 c_3_9_a c_2_11_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12746 n8388 n8394 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12745 c_2_11_cout n8390 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12744 n8386 c_2_11_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12743 vdd p_2_11_pi2j n8386 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12742 n8390 p_8_1_c2j n8386 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12741 n8390 c_2_11_a n8387 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12740 n8387 p_2_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12739 c_2_11_s2_s p_8_1_c2j n8388 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12738 vdd c_2_11_s1_s n8394 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12737 c_2_11_s1_s c_2_11_a n8396 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12736 n8396 p_2_11_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12735 n8401 p_2_2_d2j n8403 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12734 n8403 p_2_2_d2jbar n8402 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12733 n8402 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12732 vdd a_10 n8401 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12731 vdd p_2_11_t_s n8393 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12730 n8393 p_2_1_n2j p_2_11_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12729 vdd n8403 n8397 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12728 n8397 n8398 p_2_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12727 n8398 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12726 vdd n8764 n8534 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12725 n8533 p_2_1_n2j p_2_10_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12724 vdd p_2_10_t_s n8533 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12723 vdd a_8 n8536 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12722 n8535 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12721 n8767 p_2_2_d2j n8535 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12720 n8536 p_2_2_d2jbar n8767 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12719 n8764 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12718 n8534 n8767 p_2_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12717 vdd c_2_10_s1_s c_3_8_a vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12716 n8760 p_2_10_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12715 vdd c_2_10_a n8760 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12714 c_3_9_cin n8760 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12713 c_2_10_s1_s p_2_10_pi2j n8532 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12712 n8532 c_2_10_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12711 c_3_7_a c_2_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12710 n9153 n9160 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12709 c_2_9_cout n9155 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12708 n9152 c_2_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12707 vdd p_2_9_pi2j n9152 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12706 n9155 p_6_1_c2j n9152 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12705 n9155 c_2_9_a n9154 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12704 n9154 p_2_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12703 c_2_9_s2_s p_6_1_c2j n9153 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12702 vdd c_2_9_s1_s n9160 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12701 c_2_9_s1_s c_2_9_a n9161 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12700 n9161 p_2_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12699 n9170 p_2_2_d2j n9169 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12698 n9169 p_2_2_d2jbar n9168 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12697 n9168 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12696 vdd a_8 n9170 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12695 vdd p_2_9_t_s n9159 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12694 n9159 p_2_1_n2j p_2_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12693 vdd n9169 n9165 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12692 n9165 n9166 p_2_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12691 n9166 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12690 vdd n9511 n9270 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12689 n9269 p_2_1_n2j p_2_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12688 vdd p_2_8_t_s n9269 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12687 vdd a_6 n9272 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12686 n9271 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12685 n9514 p_2_2_d2j n9271 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12684 n9272 p_2_2_d2jbar n9514 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12683 n9511 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12682 n9270 n9514 p_2_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12681 vdd c_2_8_s1_s c_3_6_a vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12680 n9506 p_2_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12679 vdd c_2_8_a n9506 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12678 c_3_7_cin n9506 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12677 c_2_8_s1_s p_2_8_pi2j n9158 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12676 n9158 c_2_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12675 c_3_5_a c_2_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12674 n9950 n9957 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12673 c_2_7_cout n9949 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12672 n9948 c_2_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12671 vdd p_2_7_pi2j n9948 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12670 n9949 p_5_1_c2j n9948 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12669 n9949 c_2_7_a n9951 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12668 n9951 p_2_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12667 c_2_7_s2_s p_5_1_c2j n9950 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12666 vdd c_2_7_s1_s n9957 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12665 c_2_7_s1_s c_2_7_a n9959 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12664 n9959 p_2_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12663 n9606 p_2_2_d2j n9961 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12662 n9961 p_2_2_d2jbar n9607 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12661 n9607 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12660 vdd a_6 n9606 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12659 vdd p_2_7_t_s n9956 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12658 n9956 p_2_1_n2j p_2_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12657 vdd n9961 n9964 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12656 n9964 n9962 p_2_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12655 n9962 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12654 vdd n10284 n9965 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12653 n9955 p_2_1_n2j p_2_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12652 vdd p_2_6_t_s n9955 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12651 vdd a_4 n9968 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12650 n9967 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12649 n10283 p_2_2_d2j n9967 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12648 n9968 p_2_2_d2jbar n10283 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12647 n10284 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12646 n9965 n10283 p_2_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12645 vdd c_2_6_s1_s c_3_4_a vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12644 n10278 p_2_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12643 vdd c_2_6_a n10278 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12642 c_3_5_cin n10278 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12641 c_2_6_s1_s p_2_6_pi2j n9954 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12640 n9954 c_2_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12639 c_3_3_a c_2_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12638 n10439 n10441 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12637 c_2_5_cout n10708 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12636 n10706 c_2_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12635 vdd c_2_5_b n10706 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12634 n10708 p_4_1_c2j n10706 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12633 n10708 c_2_5_a n10707 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12632 n10707 c_2_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12631 c_2_5_s2_s p_4_1_c2j n10439 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12630 vdd c_2_5_s1_s n10441 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12629 c_2_5_s1_s c_2_5_a n10714 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12628 n10714 c_2_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12627 n10445 p_2_2_d2j n10715 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12626 n10715 p_2_2_d2jbar n10446 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12625 n10446 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12624 vdd a_4 n10445 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12623 vdd p_2_5_t_s n10442 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12622 n10442 p_2_1_n2j c_2_5_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12621 vdd n10715 n10443 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12620 n10443 n10716 p_2_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12619 n10716 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12618 vdd n10876 n10718 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12617 n10712 p_2_1_n2j p_2_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12616 vdd p_2_4_t_s n10712 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12615 vdd a_2 n10720 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12614 n10719 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12613 n10879 p_2_2_d2j n10719 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12612 n10720 p_2_2_d2jbar n10879 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12611 n10876 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12610 n10718 n10879 p_2_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12609 vdd c_2_4_s1_s c_3_2_a vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12608 n11026 p_2_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12607 vdd c_2_4_a n11026 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12606 c_3_3_cin n11026 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12605 c_2_4_s1_s p_2_4_pi2j n10711 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12604 n10711 c_2_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12603 c_3_1_a c_2_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12602 n11242 n11247 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12601 c_2_3_cout n11243 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12600 n11456 c_2_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12599 vdd c_2_3_b n11456 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12598 n11243 p_3_1_c2j n11456 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12597 n11243 c_2_3_a n11457 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12596 n11457 c_2_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12595 c_2_3_s2_s p_3_1_c2j n11242 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_12594 vdd c_2_3_s1_s n11247 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12593 c_2_3_s1_s c_2_3_a n11460 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12592 n11460 c_2_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12591 n11252 p_2_2_d2j n11254 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12590 n11254 p_2_2_d2jbar n11253 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12589 n11253 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12588 vdd a_2 n11252 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12587 vdd p_2_3_t_s n11246 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12586 n11246 p_2_1_n2j c_2_3_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12585 vdd n11254 n11249 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12584 n11249 n11250 p_2_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12583 n11250 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12582 vdd n11671 n11463 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12581 n11461 p_2_1_n2j c_2_2_b vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12580 vdd p_2_2_t_s n11461 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12579 vdd a_0 n11465 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12578 n11464 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12577 n11675 p_2_2_d2j n11464 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12576 n11465 p_2_2_d2jbar n11675 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12575 n11671 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12574 n11463 n11675 p_2_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12573 vdd c_2_2_s1_s c_2_2_sum vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_12572 n11668 c_2_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12571 vdd c_2_2_a n11668 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12570 c_3_1_cin n11668 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12569 c_2_2_s1_s c_2_2_b n11459 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12568 n11459 c_2_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12567 c_2_1_sum c_2_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12566 n12057 n12064 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12565 c_2_1_cout n12056 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12564 n12055 c_2_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12563 vdd p_2_1_pi2j n12055 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12562 n12056 n12067 n12055 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12561 n12056 c_2_1_a n12058 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12560 n12058 p_2_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12559 c_2_1_s2_s n12067 n12057 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12558 vdd c_2_1_s1_s n12064 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_12557 c_2_1_s1_s c_2_1_a n12065 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12556 n12065 p_2_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12555 n12069 n12067 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12554 n12068 n12069 p_2_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12553 vdd n12073 n12068 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12552 n12063 p_2_1_n2j p_2_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12551 vdd p_2_1_t_s n12063 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12550 vdd a_0 n12073 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12549 n12073 p_2_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12548 n12156 n12416 cl4_2_s1_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12547 vdd p_1_2_c2j n12156 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12546 p_0 cl4_2_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12545 n12410 n12416 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12544 vdd p_1_2_c2j n12410 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12543 n12411 n12410 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12542 vdd p_1_2_pi2j n12407 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_12541 n12407 n12416 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12540 vdd p_1_2_c2j n12407 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12539 n12406 n12407 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_12538 n12155 n12411 cl4_2_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12537 vdd p_1_2_pi2j n12155 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_12536 p_1 cl4_2_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_12535 p_1_33_a a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12534 vdd p_1_33_t_s n257 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12533 n257 d_0_n2j c_2_31_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12532 vdd p_1_33_a n260 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12531 n260 n261 p_1_33_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12530 n261 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12529 vdd d_0_n2j n383 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12528 vdd n592 n384 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12527 n592 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12526 vdd a_30 n385 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12525 n595 d_0_d2j n386 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12524 n386 a_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12523 n385 d_0_d2jbar n595 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12522 n383 p_1_32_t_s c_2_30_a vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12521 n384 n595 p_1_32_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12520 n973 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12519 n969 n973 p_1_31_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12518 vdd p_1_31_a n969 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12517 n965 d_0_n2j c_2_29_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12516 vdd p_1_31_t_s n965 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12515 vdd a_30 n974 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12514 n972 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12513 p_1_31_a d_0_d2jbar n972 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12512 n974 d_0_d2j p_1_31_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12511 vdd d_0_n2j n1105 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12510 vdd n1359 n1106 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12509 n1359 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12508 vdd a_28 n1107 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12507 n1362 d_0_d2j n1108 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12506 n1108 a_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12505 n1107 d_0_d2jbar n1362 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12504 n1105 p_1_30_t_s c_2_28_a vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12503 n1106 n1362 p_1_30_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12502 n1759 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12501 n1757 n1759 p_1_29_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12500 vdd p_1_29_a n1757 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12499 n1752 d_0_n2j n2555 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12498 vdd p_1_29_t_s n1752 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12497 vdd a_28 n1760 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12496 n1761 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12495 p_1_29_a d_0_d2jbar n1761 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12494 n1760 d_0_d2j p_1_29_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12493 vdd d_0_n2j n1874 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12492 vdd n2110 n1875 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12491 n2110 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12490 vdd a_26 n1876 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12489 n2112 d_0_d2j n1877 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12488 n1877 a_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12487 n1876 d_0_d2jbar n2112 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12486 n1874 p_1_28_t_s c_2_26_a vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12485 n1875 n2112 p_1_28_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12484 n2568 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12483 n2572 n2568 p_1_27_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12482 vdd p_1_27_a n2572 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12481 n2235 d_0_n2j c_2_25_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12480 vdd p_1_27_t_s n2235 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12479 vdd a_26 n2241 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12478 n2240 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12477 p_1_27_a d_0_d2jbar n2240 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12476 n2241 d_0_d2j p_1_27_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12475 vdd d_0_n2j n2569 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12474 vdd n2704 n2570 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12473 n2704 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12472 vdd a_24 n2573 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12471 n2707 d_0_d2j n2574 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12470 n2574 a_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12469 n2573 d_0_d2jbar n2707 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12468 n2569 p_1_26_t_s c_2_24_a vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12467 n2570 n2707 p_1_26_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12466 n3338 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12465 n3072 n3338 p_1_25_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12464 vdd p_1_25_a n3072 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12463 n3068 d_0_n2j c_2_23_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12462 vdd p_1_25_t_s n3068 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12461 vdd a_24 n3076 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12460 n3075 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12459 p_1_25_a d_0_d2jbar n3075 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12458 n3076 d_0_d2j p_1_25_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12457 vdd d_0_n2j n3339 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12456 vdd n3515 n3340 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12455 n3515 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12454 vdd a_22 n3341 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12453 n3518 d_0_d2j n3342 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12452 n3342 a_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12451 n3341 d_0_d2jbar n3518 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12450 n3339 p_1_24_t_s c_2_22_a vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12449 n3340 n3518 p_1_24_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12448 n3935 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12447 n3931 n3935 p_1_23_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12446 vdd p_1_23_a n3931 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12445 n3927 d_0_n2j c_2_21_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12444 vdd p_1_23_t_s n3927 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12443 vdd a_22 n3936 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12442 n3934 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12441 p_1_23_a d_0_d2jbar n3934 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12440 n3936 d_0_d2j p_1_23_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12439 vdd d_0_n2j n4096 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12438 vdd n4335 n4097 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12437 n4335 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12436 vdd a_20 n4098 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12435 n4338 d_0_d2j n4099 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12434 n4099 a_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12433 n4098 d_0_d2jbar n4338 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12432 n4096 p_1_22_t_s c_2_20_a vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12431 n4097 n4338 p_1_22_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12430 n4720 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12429 n4716 n4720 p_1_21_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12428 vdd p_1_21_a n4716 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12427 n4712 d_0_n2j c_2_19_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12426 vdd p_1_21_t_s n4712 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12425 vdd a_20 n4721 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12424 n4719 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12423 p_1_21_a d_0_d2jbar n4719 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12422 n4721 d_0_d2j p_1_21_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12421 vdd d_0_n2j n4848 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12420 vdd n5081 n4849 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12419 n5081 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12418 vdd a_18 n4850 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12417 n5084 d_0_d2j n4851 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12416 n4851 a_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12415 n4850 d_0_d2jbar n5084 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12414 n4848 p_1_20_t_s c_2_18_a vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12413 n4849 n5084 p_1_20_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12412 n5486 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12411 n5484 n5486 p_1_19_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12410 vdd p_1_19_a n5484 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12409 n5479 d_0_n2j c_2_17_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12408 vdd p_1_19_t_s n5479 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12407 vdd a_18 n5487 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12406 n5488 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12405 p_1_19_a d_0_d2jbar n5488 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12404 n5487 d_0_d2j p_1_19_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12403 vdd d_0_n2j n5600 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12402 vdd n5838 n5601 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12401 n5838 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12400 vdd a_16 n5602 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12399 n5836 d_0_d2j n5603 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12398 n5603 a_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12397 n5602 d_0_d2jbar n5836 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12396 n5600 p_1_18_t_s c_2_16_a vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12395 n5601 n5836 p_1_18_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12394 n6286 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12393 n6290 n6286 p_1_17_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12392 vdd p_1_17_a n6290 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12391 n6282 d_0_n2j c_2_15_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12390 vdd p_1_17_t_s n6282 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12389 vdd a_16 n5933 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12388 n5932 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12387 p_1_17_a d_0_d2jbar n5932 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12386 n5933 d_0_d2j p_1_17_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12385 vdd d_0_n2j n6287 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12384 vdd n6613 n6288 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12383 n6613 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12382 vdd a_14 n6291 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12381 n6402 d_0_d2j n6292 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12380 n6292 a_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12379 n6291 d_0_d2jbar n6402 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12378 n6287 p_1_16_t_s c_2_14_a vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12377 n6288 n6402 p_1_16_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12376 n7040 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12375 n6773 n7040 p_1_15_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12374 vdd p_1_15_a n6773 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12373 n6769 d_0_n2j c_2_13_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12372 vdd p_1_15_t_s n6769 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12371 vdd a_14 n6777 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12370 n6776 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12369 p_1_15_a d_0_d2jbar n6776 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12368 n6777 d_0_d2j p_1_15_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12367 vdd d_0_n2j n7041 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12366 vdd n7209 n7042 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12365 n7209 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12364 vdd a_12 n7043 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12363 n7212 d_0_d2j n7044 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12362 n7044 a_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12361 n7043 d_0_d2jbar n7212 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12360 n7041 p_1_14_t_s c_2_12_a vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12359 n7042 n7212 p_1_14_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12358 n7801 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12357 n7590 n7801 p_1_13_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12356 vdd p_1_13_a n7590 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12355 n7586 d_0_n2j c_2_11_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12354 vdd p_1_13_t_s n7586 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12353 vdd a_12 n7594 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12352 n7593 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12351 p_1_13_a d_0_d2jbar n7593 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12350 n7594 d_0_d2j p_1_13_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12349 vdd d_0_n2j n7802 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12348 vdd n8014 n7803 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12347 n8014 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12346 vdd a_10 n7804 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12345 n8017 d_0_d2j n7805 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12344 n7805 a_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12343 n7804 d_0_d2jbar n8017 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12342 n7802 p_1_12_t_s c_2_10_a vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12341 n7803 n8017 p_1_12_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12340 n8408 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12339 n8404 n8408 p_1_11_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12338 vdd p_1_11_a n8404 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12337 n8400 d_0_n2j c_2_9_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12336 vdd p_1_11_t_s n8400 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12335 vdd a_10 n8409 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12334 n8407 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12333 p_1_11_a d_0_d2jbar n8407 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12332 n8409 d_0_d2j p_1_11_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12331 vdd d_0_n2j n8537 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12330 vdd n8770 n8538 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12329 n8770 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12328 vdd a_8 n8539 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12327 n8773 d_0_d2j n8540 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12326 n8540 a_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12325 n8539 d_0_d2jbar n8773 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12324 n8537 p_1_10_t_s c_2_8_a vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12323 n8538 n8773 p_1_10_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12322 n9174 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12321 n9172 n9174 p_1_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12320 vdd p_1_9_a n9172 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12319 n9167 d_0_n2j c_2_7_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12318 vdd p_1_9_t_s n9167 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12317 vdd a_8 n9175 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12316 n9176 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12315 p_1_9_a d_0_d2jbar n9176 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12314 n9175 d_0_d2j p_1_9_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12313 vdd d_0_n2j n9273 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12312 vdd n9519 n9274 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12311 n9519 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12310 vdd a_6 n9275 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12309 n9517 d_0_d2j n9276 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12308 n9276 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12307 n9275 d_0_d2jbar n9517 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12306 n9273 p_1_8_t_s c_2_6_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12305 n9274 n9517 p_1_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12304 n9969 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12303 n9974 n9969 p_1_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12302 vdd p_1_7_a n9974 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12301 n9966 d_0_n2j c_2_5_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12300 vdd p_1_7_t_s n9966 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12299 vdd a_6 n9611 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12298 n9610 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12297 p_1_7_a d_0_d2jbar n9610 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12296 n9611 d_0_d2j p_1_7_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12295 vdd d_0_n2j n9971 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12294 vdd n10289 n9972 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12293 n10289 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12292 vdd a_4 n9976 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12291 n10287 d_0_d2j n9977 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12290 n9977 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12289 n9976 d_0_d2jbar n10287 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12288 n9971 p_1_6_t_s c_2_4_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12287 n9972 n10287 p_1_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12286 n10722 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12285 n10447 n10722 p_1_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12284 vdd p_1_5_a n10447 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12283 n10444 d_0_n2j c_2_3_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12282 vdd p_1_5_t_s n10444 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12281 vdd a_4 n10450 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12280 n10449 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12279 p_1_5_a d_0_d2jbar n10449 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12278 n10450 d_0_d2j p_1_5_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12277 vdd d_0_n2j n10723 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12276 vdd n10880 n10724 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12275 n10880 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12274 vdd a_2 n10725 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12273 n10883 d_0_d2j n10726 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12272 n10726 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12271 n10725 d_0_d2jbar n10883 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12270 n10723 p_1_4_t_s c_2_2_a vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12269 n10724 n10883 p_1_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12268 n11466 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12267 n11255 n11466 p_1_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12266 vdd p_1_3_a n11255 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12265 n11251 d_0_n2j c_2_1_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12264 vdd p_1_3_t_s n11251 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12263 vdd a_2 n11259 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12262 n11258 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12261 p_1_3_a d_0_d2jbar n11258 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12260 n11259 d_0_d2j p_1_3_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12259 vdd d_0_n2j n11467 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12258 vdd n11677 n11468 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12257 n11677 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12256 vdd a_0 n11469 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12255 n11680 d_0_d2j n11470 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12254 n11470 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12253 n11469 d_0_d2jbar n11680 vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12252 n11467 p_1_2_t_s p_1_2_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_12251 n11468 n11680 p_1_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12250 n12077 d_0_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12249 vdd a_0 n12077 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_12248 vdd p_1_1_t_s n12072 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12247 n12072 d_0_n2j n12416 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12246 vdd n12077 n12075 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12245 n12075 n12076 p_1_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12244 n12076 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_12243 n978 n1366 n979 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12242 n979 b_31 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12241 vdd b_31 n976 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12240 n976 n1373 n975 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12239 n975 n1367 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12238 vdd b_29 n979 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12237 n979 n1367 n978 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12236 n978 n1373 n979 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12235 n979 b_30 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12234 vdd p_18_2_d2j p_18_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_12233 p_18_1_c2j n976 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12232 vdd n978 p_18_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12231 p_18_2_d2j n1370 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12230 n1366 b_31 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12229 vdd n1366 n1109 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12228 n1109 b_31 n1370 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12227 n1367 b_29 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12226 n1370 n1367 n1109 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12225 n1109 b_29 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12224 n1370 n1373 n1109 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12223 n1373 b_30 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12222 n1109 b_30 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12221 n1766 n2114 n1767 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12220 n1767 b_29 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12219 vdd b_29 n1764 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12218 n1764 n2121 n1763 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12217 n1763 n2118 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12216 vdd b_27 n1767 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12215 n1767 n2118 n1766 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12214 n1766 n2121 n1767 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12213 n1767 b_28 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12212 vdd p_17_2_d2j p_17_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_12211 p_17_1_c2j n1764 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12210 vdd n1766 p_17_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12209 p_17_2_d2j n2128 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12208 n2114 b_29 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12207 vdd n2114 n1765 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12206 n1765 b_29 n2128 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12205 n2118 b_27 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12204 n2128 n2118 n1765 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12203 n1765 b_27 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12202 n2128 n2121 n1765 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12201 n2121 b_28 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12200 n1765 b_28 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12199 n2578 n2915 n2579 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12198 n2579 b_27 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12197 vdd b_27 n2576 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12196 n2576 n2921 n2575 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12195 n2575 n2917 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12194 vdd b_25 n2579 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12193 n2579 n2917 n2578 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12192 n2578 n2921 n2579 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12191 n2579 b_26 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12190 vdd p_16_2_d2j p_16_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_12189 p_16_1_c2j n2576 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12188 vdd n2578 p_16_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12187 p_16_2_d2j n2927 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12186 n2915 b_27 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12185 vdd n2915 n2577 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12184 n2577 b_27 n2927 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12183 n2917 b_25 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12182 n2927 n2917 n2577 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12181 n2577 b_25 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12180 n2927 n2921 n2577 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12179 n2921 b_26 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12178 n2577 b_26 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12177 n3080 n3521 n3081 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12176 n3081 b_25 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12175 vdd b_25 n3078 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12174 n3078 n3660 n3077 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12173 n3077 n3657 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12172 vdd b_23 n3081 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12171 n3081 n3657 n3080 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12170 n3080 n3660 n3081 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12169 n3081 b_24 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12168 vdd p_15_2_d2j p_15_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_12167 p_15_1_c2j n3078 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12166 vdd n3080 p_15_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12165 p_15_2_d2j n3668 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12164 n3521 b_25 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12163 vdd n3521 n3343 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12162 n3343 b_25 n3668 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12161 n3657 b_23 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12160 n3668 n3657 n3343 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12159 n3343 b_23 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12158 n3668 n3660 n3343 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12157 n3660 b_24 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12156 n3343 b_24 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12155 n3941 n4342 n3940 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12154 n3940 b_23 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12153 vdd b_23 n3938 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12152 n3938 n4349 n3937 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12151 n3937 n4344 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12150 vdd b_21 n3940 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12149 n3940 n4344 n3941 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12148 n3941 n4349 n3940 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12147 n3940 b_22 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12146 vdd p_14_2_d2j p_14_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_12145 p_14_1_c2j n3938 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12144 vdd n3941 p_14_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12143 p_14_2_d2j n4346 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12142 n4342 b_23 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12141 vdd n4342 n4100 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12140 n4100 b_23 n4346 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12139 n4344 b_21 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12138 n4346 n4344 n4100 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12137 n4100 b_21 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12136 n4346 n4349 n4100 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12135 n4349 b_22 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12134 n4100 b_22 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12133 n4725 n5088 n4726 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12132 n4726 b_21 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12131 vdd b_21 n4723 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12130 n4723 n5092 n4722 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12129 n4722 n5089 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12128 vdd b_19 n4726 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12127 n4726 n5089 n4725 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12126 n4725 n5092 n4726 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12125 n4726 b_20 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12124 vdd p_12_2_d2j p_12_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_12123 p_12_1_c2j n4723 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12122 vdd n4725 p_12_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12121 p_12_2_d2j n5093 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12120 n5088 b_21 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12119 vdd n5088 n4852 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12118 n4852 b_21 n5093 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12117 n5089 b_19 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12116 n5093 n5089 n4852 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12115 n4852 b_19 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12114 n5093 n5092 n4852 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12113 n5092 b_20 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12112 n4852 b_20 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12111 n5493 n5840 n5494 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12110 n5494 b_19 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12109 vdd b_19 n5491 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12108 n5491 n5846 n5490 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12107 n5490 n5844 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12106 vdd b_17 n5494 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12105 n5494 n5844 n5493 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12104 n5493 n5846 n5494 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12103 n5494 b_18 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12102 vdd p_11_2_d2j p_11_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_12101 p_11_1_c2j n5491 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12100 vdd n5493 p_11_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12099 p_11_2_d2j n5854 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12098 n5840 b_19 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12097 vdd n5840 n5492 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12096 n5492 b_19 n5854 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12095 n5844 b_17 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12094 n5854 n5844 n5492 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12093 n5492 b_17 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12092 n5854 n5846 n5492 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12091 n5846 b_18 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12090 n5492 b_18 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12089 n6296 n6616 n6297 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12088 n6297 b_17 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12087 vdd b_17 n6294 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12086 n6294 n6623 n6293 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12085 n6293 n6618 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12084 vdd b_15 n6297 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12083 n6297 n6618 n6296 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12082 n6296 n6623 n6297 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12081 n6297 b_16 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12080 vdd p_10_2_d2j p_10_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_12079 p_10_1_c2j n6294 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12078 vdd n6296 p_10_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12077 p_10_2_d2j n6628 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12076 n6616 b_17 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12075 vdd n6616 n6295 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12074 n6295 b_17 n6628 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12073 n6618 b_15 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12072 n6628 n6618 n6295 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12071 n6295 b_15 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12070 n6628 n6623 n6295 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12069 n6623 b_16 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12068 n6295 b_16 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12067 n7048 n7214 n7049 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12066 n7049 b_15 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12065 vdd b_15 n7046 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12064 n7046 n7371 n7045 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12063 n7045 n7367 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12062 vdd b_13 n7049 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12061 n7049 n7367 n7048 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12060 n7048 n7371 n7049 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12059 n7049 b_14 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12058 vdd p_9_2_d2j p_9_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_12057 p_9_1_c2j n7046 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12056 vdd n7048 p_9_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12055 p_9_2_d2j n7377 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12054 n7214 b_15 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12053 vdd n7214 n7047 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12052 n7047 b_15 n7377 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12051 n7367 b_13 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12050 n7377 n7367 n7047 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12049 n7047 b_13 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12048 n7377 n7371 n7047 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12047 n7371 b_14 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12046 n7047 b_14 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12045 n7598 n8020 n7599 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12044 n7599 b_13 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12043 vdd b_13 n7596 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12042 n7596 n8027 n7595 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12041 n7595 n8023 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12040 vdd b_11 n7599 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12039 n7599 n8023 n7598 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12038 n7598 n8027 n7599 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12037 n7599 b_12 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12036 vdd p_8_2_d2j p_8_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_12035 p_8_1_c2j n7596 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12034 vdd n7598 p_8_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12033 p_8_2_d2j n8024 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12032 n8020 b_13 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12031 vdd n8020 n7806 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12030 n7806 b_13 n8024 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12029 n8023 b_11 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12028 n8024 n8023 n7806 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12027 n7806 b_11 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12026 n8024 n8027 n7806 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12025 n8027 b_12 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12024 n7806 b_12 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12023 n8413 n8778 n8414 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12022 n8414 b_11 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12021 vdd b_11 n8411 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12020 n8411 n8781 n8410 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12019 n8410 n8775 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12018 vdd b_9 n8414 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12017 n8414 n8775 n8413 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12016 n8413 n8781 n8414 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12015 n8414 b_10 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12014 vdd p_6_2_d2j p_6_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_12013 p_6_1_c2j n8411 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12012 vdd n8413 p_6_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12011 p_6_2_d2j n8782 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12010 n8778 b_11 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12009 vdd n8778 n8541 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12008 n8541 b_11 n8782 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12007 n8775 b_9 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12006 n8782 n8775 n8541 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12005 n8541 b_9 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12004 n8782 n8781 n8541 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12003 n8781 b_10 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12002 n8541 b_10 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_12001 n9180 n9525 n9181 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_12000 n9181 b_9 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11999 vdd b_9 n9179 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11998 n9179 n9528 n9178 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11997 n9178 n9526 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11996 vdd b_7 n9181 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11995 n9181 n9526 n9180 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11994 n9180 n9528 n9181 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11993 n9181 b_8 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11992 vdd p_5_2_d2j p_5_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_11991 p_5_1_c2j n9179 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11990 vdd n9180 p_5_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11989 p_5_2_d2j n9529 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11988 n9525 b_9 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11987 vdd n9525 n9277 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11986 n9277 b_9 n9529 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11985 n9526 b_7 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11984 n9529 n9526 n9277 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11983 n9277 b_7 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11982 n9529 n9528 n9277 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11981 n9528 b_8 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11980 n9277 b_8 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11979 n9981 n10293 n9982 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11978 n9982 b_7 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11977 vdd b_7 n9979 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11976 n9979 n10300 n9978 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11975 n9978 n10298 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11974 vdd b_5 n9982 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11973 n9982 n10298 n9981 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11972 n9981 n10300 n9982 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11971 n9982 b_6 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11970 vdd p_4_2_d2j p_4_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_11969 p_4_1_c2j n9979 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11968 vdd n9981 p_4_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11967 p_4_2_d2j n10305 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11966 n10293 b_7 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11965 vdd n10293 n9980 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11964 n9980 b_7 n10305 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11963 n10298 b_5 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11962 n10305 n10298 n9980 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11961 n9980 b_5 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11960 n10305 n10300 n9980 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11959 n10300 b_6 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11958 n9980 b_6 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11957 n10730 n10885 n10731 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11956 n10731 b_5 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11955 vdd b_5 n10728 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11954 n10728 n11042 n10727 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11953 n10727 n11038 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11952 vdd b_3 n10731 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11951 n10731 n11038 n10730 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11950 n10730 n11042 n10731 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11949 n10731 b_4 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11948 vdd p_3_2_d2j p_3_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_11947 p_3_1_c2j n10728 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11946 vdd n10730 p_3_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11945 p_3_2_d2j n11048 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11944 n10885 b_5 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11943 vdd n10885 n10729 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11942 n10729 b_5 n11048 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11941 n11038 b_3 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11940 n11048 n11038 n10729 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11939 n10729 b_3 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11938 n11048 n11042 n10729 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11937 n11042 b_4 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11936 n10729 b_4 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11935 n11263 n11683 n11264 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11934 n11264 b_3 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11933 vdd b_3 n11261 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11932 n11261 n11690 n11260 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11931 n11260 n11685 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11930 vdd b_1 n11264 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11929 n11264 n11685 n11263 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11928 n11263 n11690 n11264 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11927 n11264 b_2 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11926 vdd p_2_2_d2j p_2_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_11925 n12067 n11261 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11924 vdd n11263 p_2_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11923 p_2_2_d2j n11687 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11922 n11683 b_3 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11921 vdd n11683 n11471 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11920 n11471 b_3 n11687 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11919 n11685 b_1 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11918 n11687 n11685 n11471 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11917 n11471 b_1 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11916 n11687 n11690 n11471 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11915 n11690 b_2 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11914 n11471 b_2 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11913 n12157 b_0 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11912 n12430 b_0 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11911 n12427 n12430 n12157 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11910 n12157 vss vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11909 n12427 n12423 n12157 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11908 n12423 vss vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11907 n12157 b_1 n12427 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11906 vdd n12421 n12157 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11905 n12421 b_1 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11904 d_0_d2j n12427 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11903 vdd n12083 d_0_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11902 p_1_2_c2j n12080 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11901 vdd d_0_d2j d_0_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11900 n12082 b_0 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11899 n12083 n12430 n12082 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11898 n12082 n12423 n12083 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11897 vdd vss n12082 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11896 n12079 n12423 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11895 n12080 n12430 n12079 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11894 vdd b_1 n12080 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11893 n12082 b_1 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_11892 n12083 n12421 n12082 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_11891 c_18_1_sum cla_cell0_0_a n12163 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11890 n12163 c_18_1_sum cla_cell0_0_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11889 vss n12163 p_30 vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_11888 vss cla_cell0_0_a n12160 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11887 n12160 c_18_1_sum n12161 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11886 vss n12161 cla_cell0_0_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11885 c_18_2_sum c_18_1_cout n11787 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11884 n11787 c_18_2_sum c_18_1_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11883 vss n11787 cla_cell0_1_p vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11882 vss c_18_1_cout n11692 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11881 n11692 c_18_2_sum n11783 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11880 vss n11783 cla_cell0_1_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11879 vss n11479 cla_cell0_2_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11878 n11480 c_18_2_cout n11479 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11877 vss c_18_3_sum n11480 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11876 c_18_2_cout c_18_3_sum n11481 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11875 n11481 c_18_2_cout c_18_3_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11874 cla_cell0_2_p n11481 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11873 vss cla_cell0_2_p cla_cell0_2_pn vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11872 c_18_4_sum c_18_3_cout n11059 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11871 n11059 c_18_4_sum c_18_3_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11870 vss n11059 cla_cell1_3_p1 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11869 vss c_18_3_cout n10896 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11868 n10896 c_18_4_sum n11270 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11867 vss n11270 cla_cell0_3_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11866 c_18_4_cout c_18_5_sum n10899 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11865 n10899 c_18_4_cout c_18_5_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11864 vss n10899 cla_cell3_4_p1 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11863 vss c_18_5_sum n10895 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11862 n10895 c_18_4_cout n10893 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11861 vss n10893 cla_cell0_4_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11860 vss n10461 cla_cell0_5_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11859 n10075 c_18_6_sum n10461 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11858 vss c_18_5_cout n10075 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11857 c_18_6_sum c_18_5_cout n10465 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11856 n10465 c_18_6_sum c_18_5_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11855 cla_cell1_5_p1 n10465 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11854 vss cla_cell1_5_p1 cla_cell7_5_p vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11853 vss n10073 cla_cell1_6_tsg vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11852 n10074 c_18_6_cout n10073 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11851 vss c_18_7_sum n10074 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11850 c_18_6_cout c_18_7_sum n10079 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11849 n10079 c_18_6_cout c_18_7_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11848 cla_cell0_6_p n10079 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11847 vss cla_cell0_6_p cla_cell7_6_p vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11846 vss n9630 cla_cell0_7_g vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_11845 n9288 c_18_8_sum n9630 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11844 vss c_18_7_cout n9288 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11843 c_18_8_sum c_18_7_cout n9634 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11842 n9634 c_18_8_sum c_18_7_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11841 cla_cell0_7_p n9634 vss vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_11840 vss cla_cell0_7_p cla_cell0_7_pn vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11839 vss n9289 cla_cell0_8_g vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_11838 n9287 c_18_8_cout n9289 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11837 vss c_18_9_sum n9287 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11836 c_18_8_cout c_18_9_sum n9292 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11835 n9292 c_18_8_cout c_18_9_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11834 cla_cell0_8_p n9292 vss vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_11833 vss cla_cell0_8_p cla_cell7_8_p vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11832 c_18_10_sum c_18_9_cout n8869 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11831 n8869 c_18_10_sum c_18_9_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11830 vss n8869 cla_cell0_9_p vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_11829 vss c_18_9_cout n8788 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11828 n8788 c_18_10_sum n8862 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11827 vss n8862 cla_cell0_9_g vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_11826 c_18_10_cout c_18_11_sum n8561 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11825 n8561 c_18_10_cout c_18_11_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11824 vss n8561 cla_cell0_10_p vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11823 vss c_18_11_sum n8558 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11822 n8558 c_18_10_cout n8557 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11821 vss n8557 cla_cell0_10_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11820 c_18_12_sum c_18_11_cout n8132 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11819 n8132 c_18_12_sum c_18_11_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11818 vss n8132 cla_cell0_11_p vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11817 vss c_18_11_cout n8031 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11816 n8031 c_18_12_sum n8126 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11815 vss n8126 cla_cell0_11_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11814 c_18_12_cout c_18_13_sum n7820 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11813 n7820 c_18_12_cout c_18_13_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11812 vss n7820 cla_cell0_12_p vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11811 vss c_18_13_sum n7816 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11810 n7816 c_18_12_cout n7815 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11809 vss n7815 cla_cell0_12_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11808 c_18_14_sum c_18_13_cout n7393 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11807 n7393 c_18_14_sum c_18_13_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11806 vss n7393 cla_cell0_13_p vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11805 vss c_18_13_cout n7228 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11804 n7228 c_18_14_sum n7604 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11803 vss n7604 cla_cell0_13_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11802 c_18_14_cout c_18_15_sum n7230 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11801 n7230 c_18_14_cout c_18_15_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11800 vss n7230 cla_cell0_14_p vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11799 vss c_18_15_sum n7227 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11798 n7227 c_18_14_cout n7059 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11797 vss n7059 cla_cell0_14_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11796 c_18_16_sum c_18_15_cout n6799 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11795 n6799 c_18_16_sum c_18_15_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11794 vss n6799 cla_cell1_15_p1 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11793 vss c_18_15_cout n6416 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11792 n6416 c_18_16_sum n6795 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11791 vss n6795 cla_cell0_15_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11790 c_18_16_cout c_18_17_sum n6419 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11789 n6419 c_18_16_cout c_18_17_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11788 vss n6419 cla_cell5_16_p1 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11787 vss c_18_17_sum n6414 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11786 n6414 c_18_16_cout n6415 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11785 vss n6415 cla_cell1_16_sg vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11784 vss n5946 cla_cell0_17_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11783 n5622 c_18_18_sum n5946 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11782 vss c_18_17_cout n5622 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11781 c_18_18_sum c_18_17_cout n5950 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11780 n5950 c_18_18_sum c_18_17_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11779 cla_cell0_17_p n5950 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11778 vss cla_cell0_17_p cla_cell0_17_pn vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11777 vss n5620 cla_cell1_18_tsg vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11776 n5621 c_18_18_cout n5620 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11775 vss c_18_19_sum n5621 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11774 c_18_18_cout c_18_19_sum n5625 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11773 n5625 c_18_18_cout c_18_19_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11772 cla_cell0_18_p n5625 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11771 vss cla_cell0_18_p cla_cell7_18_p vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11770 vss n5173 cla_cell0_19_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11769 n4868 c_18_20_sum n5173 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11768 vss c_18_19_cout n4868 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11767 c_18_20_sum c_18_19_cout n5180 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11766 n5180 c_18_20_sum c_18_19_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11765 cla_cell0_19_p n5180 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11764 vss cla_cell0_19_p cla_cell0_19_pn vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11763 vss n4866 cla_cell0_20_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11762 n4867 c_18_20_cout n4866 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11761 vss c_18_21_sum n4867 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11760 c_18_20_cout c_18_21_sum n4871 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11759 n4871 c_18_20_cout c_18_21_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11758 cla_cell0_20_p n4871 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11757 vss cla_cell0_20_p cla_cell0_20_pn vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11756 vss n4437 cla_cell0_21_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11755 n4355 c_18_22_sum n4437 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11754 vss c_18_21_cout n4355 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11753 c_18_22_sum c_18_21_cout n4441 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11752 n4441 c_18_22_sum c_18_21_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11751 cla_cell0_21_p n4441 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11750 vss cla_cell0_21_p cla_cell0_21_pn vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11749 vss n4122 cla_cell0_22_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11748 n4120 c_18_22_cout n4122 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11747 vss c_18_23_sum n4120 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11746 c_18_22_cout c_18_23_sum n4126 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11745 n4126 c_18_22_cout c_18_23_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11744 cla_cell0_22_p n4126 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11743 vss cla_cell0_22_p cla_cell0_22_pn vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11742 vss n3683 cla_cell0_23_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11741 n3533 c_18_24_sum n3683 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11740 vss c_18_23_cout n3533 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11739 c_18_24_sum c_18_23_cout n3689 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11738 n3689 c_18_24_sum c_18_23_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11737 cla_cell0_23_p n3689 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11736 vss cla_cell0_23_p cla_cell0_23_pn vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11735 vss n3349 cla_cell0_24_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11734 n3532 c_18_24_cout n3349 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11733 vss c_18_25_sum n3532 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11732 c_18_24_cout c_18_25_sum n3351 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11731 n3351 c_18_24_cout c_18_25_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11730 cla_cell0_24_p n3351 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11729 vss cla_cell0_24_p cla_cell0_24_pn vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11728 vss n3093 cla_cell0_25_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11727 n2729 c_18_26_sum n3093 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11726 vss c_18_25_cout n2729 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11725 c_18_26_sum c_18_25_cout n3097 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11724 n3097 c_18_26_sum c_18_25_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11723 cla_cell1_25_p1 n3097 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11722 vss cla_cell1_25_p1 cla_cell0_25_pn vss TN L=0.18U W=1.08U 
+ AS=0.3888P AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11721 vss n2727 cla_cell1_26_tsg vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11720 n2728 c_18_26_cout n2727 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11719 vss c_18_27_sum n2728 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11718 c_18_26_cout c_18_27_sum n2732 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11717 n2732 c_18_26_cout c_18_27_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11716 cla_cell0_26_p n2732 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11715 vss cla_cell0_26_p cla_cell7_26_p vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11714 vss n2261 cla_cell0_27_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11713 n1895 c_18_28_sum n2261 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11712 vss c_18_27_cout n1895 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11711 c_18_28_sum c_18_27_cout n2266 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11710 n2266 c_18_28_sum c_18_27_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11709 cla_cell0_27_p n2266 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11708 vss cla_cell0_27_p cla_cell7_27_p vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11707 vss n1896 cla_cell3_28_g1 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11706 n1894 c_18_28_cout n1896 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11705 vss c_18_29_sum n1894 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11704 c_18_28_cout c_18_29_sum n1899 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11703 n1899 c_18_28_cout c_18_29_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11702 cla_cell0_28_p n1899 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11701 vss cla_cell0_28_p cla_cell7_28_p vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11700 vss n1447 cla_cell0_29_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11699 n1130 c_18_30_sum n1447 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11698 vss c_18_29_cout n1130 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11697 c_18_30_sum c_18_29_cout n1455 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11696 n1455 c_18_30_sum c_18_29_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11695 cla_cell0_29_p n1455 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11694 vss cla_cell0_29_p cla_cell0_29_pn vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11693 vss n1131 cla_cell0_30_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11692 n1129 c_18_30_cout n1131 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11691 vss c_18_31_sum n1129 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11690 c_18_30_cout c_18_31_sum n1135 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11689 n1135 c_18_30_cout c_18_31_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11688 cla_cell0_30_p n1135 vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11687 vss cla_cell0_30_p cla_cell0_30_pn vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11686 vss n689 cla_cell0_31_g vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_11685 n604 c_18_32_sum n689 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11684 vss c_18_31_cout n604 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11683 c_18_32_sum c_18_31_cout n694 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11682 n694 c_18_32_sum c_18_31_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11681 cla_cell0_31_p n694 vss vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_11680 vss cla_cell0_31_p cla_cell0_31_pn vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11679 vss n394 cla_cell0_32_g vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_11678 n392 c_18_32_cout n394 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11677 vss cla_cell0_32_a n392 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11676 c_18_32_cout cla_cell0_32_a n398 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11675 n398 c_18_32_cout cla_cell0_32_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11674 cla_cell0_32_p n398 vss vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_11673 vss cla_cell0_32_p cla_cell0_32_pn vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11672 cla_cell0_32_a cla_cell0_33_a n46 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11671 n46 cla_cell0_32_a cla_cell0_33_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11670 vss n46 cla_cell0_33_p vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_11669 vss cla_cell0_33_a n4 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11668 n4 cla_cell0_32_a n41 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11667 vss n41 cla_cell0_33_g vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_11666 vss cla_cell0_0_g n11691 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_11665 n11691 cla_cell0_1_p cla_cell1_1_co vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_11664 cla_cell1_1_co cla_cell0_1_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11663 cla_cell1_2_ng cla_cell0_2_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11662 vss cla_cell0_2_p cla_cell1_2_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11661 vss cla_cell0_2_g n10894 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11660 n10894 cla_cell1_3_p1 cla_cell1_3_g vss TN L=0.18U W=1.62U 
+ AS=0.5832P AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11659 cla_cell1_3_g cla_cell0_3_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11658 vss cla_cell1_3_p1 n10892 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11657 n10892 cla_cell0_2_p n11054 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11656 n11054 cla_cell0_2_p n10892 vss TN L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_11655 vss cla_cell0_4_g n10072 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11654 n10072 cla_cell1_5_p1 cla_cell2_5_tsg vss TN L=0.18U W=1.62U 
+ AS=0.5832P AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11653 cla_cell2_5_tsg cla_cell0_5_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11652 vss cla_cell1_5_p1 n10069 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11651 n10069 cla_cell3_4_p1 cla_cell2_5_tsp vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11650 cla_cell2_5_tsp cla_cell3_4_p1 n10069 vss TN L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_11649 cla_cell1_6_ng cla_cell1_6_tsg vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11648 vss cla_cell0_6_p cla_cell1_6_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11647 vss cla_cell1_6_tsg n9285 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11646 n9285 cla_cell0_7_p cla_cell1_7_g vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11645 cla_cell1_7_g cla_cell0_7_g vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11644 n9283 cla_cell0_6_p cla_cell2_7_pl vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11643 vss cla_cell0_7_p n9283 vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_11642 cla_cell1_8_ng cla_cell0_8_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11641 vss cla_cell0_8_p cla_cell1_8_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11640 vss cla_cell0_8_g n8787 vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_11639 n8787 cla_cell0_9_p cla_cell1_9_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11638 cla_cell1_9_g cla_cell0_9_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11637 vss cla_cell0_9_p n8786 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11636 n8786 cla_cell0_8_p cla_cell2_9_sp vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11635 cla_cell2_9_sp cla_cell0_8_p n8786 vss TN L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_11634 cla_cell1_10_ng cla_cell0_10_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11633 vss cla_cell0_10_p cla_cell1_10_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11632 vss cla_cell0_10_g n8030 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11631 n8030 cla_cell0_11_p cla_cell1_11_g vss TN L=0.18U W=1.62U 
+ AS=0.5832P AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11630 cla_cell1_11_g cla_cell0_11_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11629 vss cla_cell0_11_p n8029 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11628 n8029 cla_cell0_10_p n8124 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11627 n8124 cla_cell0_10_p n8029 vss TN L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_11626 vss cla_cell0_12_g n7226 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11625 n7226 cla_cell0_13_p cla_cell1_13_g vss TN L=0.18U W=1.62U 
+ AS=0.5832P AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11624 cla_cell1_13_g cla_cell0_13_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11623 vss cla_cell0_13_p n7224 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11622 n7224 cla_cell0_12_p cla_cell2_13_tsp vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11621 cla_cell2_13_tsp cla_cell0_12_p n7224 vss TN L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_11620 cla_cell1_14_ng cla_cell0_14_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11619 vss cla_cell0_14_p cla_cell1_14_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11618 vss cla_cell0_14_g n6413 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11617 n6413 cla_cell1_15_p1 cla_cell2_15_gl vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11616 cla_cell2_15_gl cla_cell0_15_g vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11615 n6412 cla_cell0_14_p cla_cell2_15_pl vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11614 vss cla_cell1_15_p1 n6412 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11613 vss cla_cell1_16_sg n5619 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11612 n5619 cla_cell0_17_p cla_cell1_17_g vss TN L=0.18U W=1.62U 
+ AS=0.5832P AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11611 cla_cell1_17_g cla_cell0_17_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11610 vss cla_cell0_17_p n5856 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11609 n5856 cla_cell5_16_p1 cla_cell2_17_tsp vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11608 cla_cell2_17_tsp cla_cell5_16_p1 n5856 vss TN L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_11607 cla_cell1_18_ng cla_cell1_18_tsg vss vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11606 vss cla_cell0_18_p cla_cell1_18_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11605 vss cla_cell1_18_tsg n4864 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11604 n4864 cla_cell0_19_p cla_cell1_19_g vss TN L=0.18U W=1.62U 
+ AS=0.5832P AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11603 cla_cell1_19_g cla_cell0_19_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11602 vss cla_cell0_19_p n5096 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11601 n5096 cla_cell0_18_p n5172 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11600 n5172 cla_cell0_18_p n5096 vss TN L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_11599 vss cla_cell0_20_g n4354 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11598 n4354 cla_cell0_21_p cla_cell1_21_g vss TN L=0.18U W=1.62U 
+ AS=0.5832P AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11597 cla_cell1_21_g cla_cell0_21_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11596 vss cla_cell0_21_p n4353 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11595 n4353 cla_cell0_20_p cla_cell2_21_tsp vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11594 cla_cell2_21_tsp cla_cell0_20_p n4353 vss TN L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_11593 cla_cell1_22_ng cla_cell0_22_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11592 vss cla_cell0_22_p cla_cell1_22_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11591 vss cla_cell0_22_g n3531 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11590 n3531 cla_cell0_23_p cla_cell1_23_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11589 cla_cell1_23_g cla_cell0_23_g vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11588 n3529 cla_cell0_22_p cla_cell2_23_pl vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11587 vss cla_cell0_23_p n3529 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11586 cla_cell1_24_ng cla_cell0_24_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11585 vss cla_cell0_24_p cla_cell1_24_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11584 vss cla_cell0_24_g n2726 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11583 n2726 cla_cell1_25_p1 cla_cell4_25_gl vss TN L=0.18U W=1.62U 
+ AS=0.5832P AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11582 cla_cell4_25_gl cla_cell0_25_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11581 vss cla_cell1_25_p1 n2723 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11580 n2723 cla_cell0_24_p cla_cell2_25_sp vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11579 cla_cell2_25_sp cla_cell0_24_p n2723 vss TN L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_11578 cla_cell1_26_ng cla_cell1_26_tsg vss vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11577 vss cla_cell0_26_p cla_cell1_26_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11576 vss cla_cell1_26_tsg n1893 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11575 n1893 cla_cell0_27_p cla_cell1_27_g vss TN L=0.18U W=1.62U 
+ AS=0.5832P AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11574 cla_cell1_27_g cla_cell0_27_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11573 vss cla_cell0_27_p n1892 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11572 n1892 cla_cell0_26_p n2260 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11571 n2260 cla_cell0_26_p n1892 vss TN L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_11570 vss cla_cell3_28_g1 n1128 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11569 n1128 cla_cell0_29_p cla_cell1_29_g vss TN L=0.18U W=1.62U 
+ AS=0.5832P AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11568 cla_cell1_29_g cla_cell0_29_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11567 vss cla_cell0_29_p n1377 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11566 n1377 cla_cell0_28_p cla_cell2_29_tsp vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11565 cla_cell2_29_tsp cla_cell0_28_p n1377 vss TN L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_11564 cla_cell1_30_ng cla_cell0_30_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11563 vss cla_cell0_30_p cla_cell1_30_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11562 vss cla_cell0_30_g n603 vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_11561 n603 cla_cell0_31_p cla_cell1_31_g vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11560 cla_cell1_31_g cla_cell0_31_g vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11559 n602 cla_cell0_30_p cla_cell2_31_pl vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11558 vss cla_cell0_31_p n602 vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_11557 cla_cell1_32_ng cla_cell0_32_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11556 vss cla_cell0_32_p cla_cell1_32_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11555 vss cla_cell0_32_g n3 vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_11554 n3 cla_cell0_33_p cla_cell1_33_g vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11553 cla_cell1_33_g cla_cell0_33_g vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11552 n2 cla_cell0_32_p n39 vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_11551 vss cla_cell0_33_p n2 vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_11550 n11476 cla_cell1_2_np vss vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11549 n11476 cla_cell1_2_ng cla_cell7_2_g vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11548 vss cla_cell1_1_co n11476 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11547 n10891 cla_cell1_3_g cla_cell3_4_g2 vss TN L=0.18U W=3.06U 
+ AS=1.1016P AD=1.1016P PS=6.84U PD=6.84U 
Mtr_11546 n10891 n11054 vss vss TN L=0.18U W=3.06U AS=1.1016P AD=1.1016P 
+ PS=6.84U PD=6.84U 
Mtr_11545 vss cla_cell1_1_co n10891 vss TN L=0.18U W=3.06U AS=1.1016P 
+ AD=1.1016P PS=6.84U PD=6.84U 
Mtr_11544 cla_cell2_5_ng cla_cell2_5_tsg vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11543 vss cla_cell2_5_tsp cla_cell2_5_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11542 vss cla_cell2_5_tsp cla_cell3_6_p1 vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11541 vss cla_cell1_6_np cla_cell3_6_p1 vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11540 n10068 cla_cell1_6_ng cla_cell2_6_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11539 vss cla_cell1_6_np n10068 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11538 n10068 cla_cell2_5_tsg vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11537 vss cla_cell2_5_tsp cla_cell3_7_p1 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11536 vss cla_cell2_7_pl cla_cell3_7_p1 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11535 n9534 cla_cell1_7_g cla_cell2_7_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11534 vss cla_cell2_7_pl n9534 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11533 n9534 cla_cell2_5_tsg vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11532 cla_cell2_10_g1 n8553 vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11531 n8551 n8549 vss vss TN L=0.18U W=0.72U AS=0.2592P AD=0.2592P 
+ PS=2.16U PD=2.16U 
Mtr_11530 cla_cell2_10_p_s n8546 cla_cell2_9_sp vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11529 cla_cell2_10_g_s n8546 cla_cell1_9_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11528 cla_cell1_11_g n8124 cla_cell2_10_g_s vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11527 vss n8124 n8546 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11526 cla_cell2_10_sg cla_cell2_10_g_s vss vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11525 n8121 cla_cell2_10_sp vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11524 vss cla_cell2_10_sg cla_cell2_10_g2 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11523 vss cla_cell2_10_p_s cla_cell2_10_sp vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11522 n8554 cla_cell1_10_ng n8553 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11521 n8554 cla_cell1_9_g vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_11520 vss cla_cell1_10_np n8554 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11519 vss cla_cell1_10_np n8549 vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11518 vss cla_cell2_9_sp n8549 vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11517 vdd n8124 cla_cell2_10_p_s vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_11516 cla_cell2_13_ng cla_cell1_13_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11515 vss cla_cell2_13_tsp cla_cell2_13_np vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11514 vss cla_cell2_13_tsp cla_cell3_14_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11513 vss cla_cell1_14_np cla_cell3_14_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11512 n7223 cla_cell1_14_ng cla_cell2_14_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11511 vss cla_cell1_14_np n7223 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11510 n7223 cla_cell1_13_g vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11509 vss cla_cell2_13_tsp cla_cell3_15_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11508 vss cla_cell2_15_pl cla_cell3_15_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11507 n6635 cla_cell2_15_gl cla_cell2_15_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11506 vss cla_cell2_15_pl n6635 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11505 n6635 cla_cell1_13_g vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11504 cla_cell2_17_ng cla_cell1_17_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11503 vss cla_cell2_17_tsp cla_cell2_17_np vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11502 vdd n5172 cla_cell2_18_p_s vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_11501 vss cla_cell2_17_tsp cla_cell5_18_p1 vss TN L=0.18U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11500 vss cla_cell1_18_np cla_cell5_18_p1 vss TN L=0.18U W=0.54U 
+ AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11499 vss cla_cell1_18_np n5615 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11498 n5615 cla_cell1_17_g vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11497 n5615 cla_cell1_18_ng cla_cell2_18_g1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11496 vss cla_cell2_18_p_s cla_cell2_18_sp vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11495 cla_cell2_18_sg cla_cell2_18_g_s vss vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11494 vss n5172 n5611 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11493 cla_cell1_19_g n5172 cla_cell2_18_g_s vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11492 cla_cell2_18_g_s n5611 cla_cell1_17_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11491 cla_cell2_18_p_s n5611 cla_cell2_17_tsp vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11490 cla_cell2_21_ng cla_cell1_21_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11489 vss cla_cell2_21_tsp cla_cell2_21_np vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11488 vss cla_cell2_21_tsp cla_cell3_22_p11 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11487 vss cla_cell1_22_np cla_cell3_22_p11 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11486 n4117 cla_cell1_22_ng cla_cell2_22_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11485 vss cla_cell1_22_np n4117 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11484 n4117 cla_cell1_21_g vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11483 vss cla_cell2_21_tsp cla_cell3_22_p21 vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11482 vss cla_cell2_23_pl cla_cell3_22_p21 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11481 n3528 cla_cell1_23_g cla_cell2_23_g vss TN L=0.18U W=1.62U 
+ AS=0.5832P AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11480 vss cla_cell2_23_pl n3528 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11479 n3528 cla_cell1_21_g vss vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11478 cla_cell2_26_g1 n2586 vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11477 cla_cell4_26_pl n2718 vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11476 cla_cell2_26_p_s n2717 cla_cell2_25_sp vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11475 cla_cell2_26_g_s n2717 cla_cell4_25_gl vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11474 cla_cell1_27_g n2260 cla_cell2_26_g_s vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11473 vss n2260 n2717 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11472 cla_cell2_26_sg cla_cell2_26_g_s vss vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11471 cla_cell4_27_pl cla_cell2_26_sp vss vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11470 vss cla_cell2_26_sg cla_cell4_27_gl vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11469 vss cla_cell2_26_p_s cla_cell2_26_sp vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11468 n2722 cla_cell1_26_ng n2586 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11467 n2722 cla_cell4_25_gl vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11466 vss cla_cell1_26_np n2722 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11465 vss cla_cell1_26_np n2718 vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11464 vss cla_cell2_25_sp n2718 vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11463 vdd n2260 cla_cell2_26_p_s vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_11462 cla_cell2_29_ng cla_cell1_29_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11461 vss cla_cell2_29_tsp cla_cell2_29_np vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11460 vss cla_cell2_29_tsp cla_cell3_30_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11459 vss cla_cell1_30_np cla_cell3_30_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11458 n1124 cla_cell1_30_ng cla_cell2_30_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11457 vss cla_cell1_30_np n1124 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11456 n1124 cla_cell1_29_g vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11455 vss cla_cell2_29_tsp cla_cell3_31_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11454 vss cla_cell2_31_pl cla_cell3_31_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11453 n601 cla_cell1_31_g cla_cell2_31_g vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11452 vss cla_cell2_31_pl n601 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11451 n601 cla_cell1_29_g vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_11450 vss cla_cell3_4_g2 n10890 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11449 n10890 cla_cell3_4_p1 cla_cell3_4_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11448 cla_cell3_4_co cla_cell0_4_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11447 vss cla_cell3_4_g2 n10065 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11446 n10065 cla_cell2_5_np cla_cell3_5_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11445 cla_cell3_5_co cla_cell2_5_ng vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11444 vss cla_cell3_4_g2 n10063 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11443 n10063 cla_cell3_6_p1 cla_cell3_6_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11442 cla_cell3_6_co cla_cell2_6_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11441 vss cla_cell3_7_p1 n9532 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11440 n9624 n9532 cla_cell2_7_g vss TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_11439 cla_cell3_4_g2 cla_cell3_7_p1 n9624 vss TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
Mtr_11438 vss n9624 cla_cell4_8_g2 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_11437 vss cla_cell2_10_sg n7812 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11436 n7812 cla_cell0_12_p cla_cell3_12_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11435 cla_cell3_12_g cla_cell0_12_g vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11434 n7811 cla_cell2_10_sp n7813 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11433 vss cla_cell0_12_p n7811 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11432 vss cla_cell2_10_sg n7220 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11431 n7220 cla_cell2_13_np cla_cell3_13_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11430 cla_cell3_13_g cla_cell2_13_ng vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11429 n7221 cla_cell2_10_sp n7384 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11428 vss cla_cell2_13_np n7221 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11427 vss cla_cell2_10_sg n7219 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11426 n7219 cla_cell3_14_p1 cla_cell3_14_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11425 cla_cell3_14_g cla_cell2_14_g vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11424 n7053 cla_cell2_10_sp n7052 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11423 vss cla_cell3_14_p1 n7053 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11422 vss cla_cell2_10_sg n6410 vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11421 n6410 cla_cell3_15_p1 cla_cell3_15_g vss TN L=0.18U W=1.62U 
+ AS=0.5832P AD=0.5832P PS=3.96U PD=3.96U 
Mtr_11420 cla_cell3_15_g cla_cell2_15_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11419 vss cla_cell3_15_p1 n6411 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11418 n6411 cla_cell2_10_sp cla_cell4_15_p1 vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11417 cla_cell4_15_p1 cla_cell2_10_sp n6411 vss TN L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_11416 vss cla_cell2_18_sg n4861 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11415 n4861 cla_cell0_20_p cla_cell3_20_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11414 cla_cell3_20_g cla_cell0_20_g vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11413 n4860 cla_cell2_18_sp cla_cell4_20_p vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11412 vss cla_cell0_20_p n4860 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11411 vss cla_cell2_18_sg n4352 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11410 n4352 cla_cell2_21_np cla_cell3_21_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11409 cla_cell3_21_g cla_cell2_21_ng vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11408 n4351 cla_cell2_18_sp cla_cell4_21_p vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11407 vss cla_cell2_21_np n4351 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11406 cla_cell5_22_p1 n4114 vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11405 cla_cell3_22_g1 n4112 vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11404 vss n4105 n4108 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P PS=3.6U 
+ PD=3.6U 
Mtr_11403 n4108 cla_cell3_22_p21 cla_cell2_18_sp vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11402 n3676 n4105 cla_cell2_23_g vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11401 cla_cell2_18_sg cla_cell3_22_p21 n3676 vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11400 vss cla_cell3_22_p21 n4105 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11399 cla_cell3_22_sg n3676 vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11398 cla_cell5_23_p1 cla_cell3_22_sp vss vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11397 vss cla_cell3_22_sg cla_cell3_22_g2 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11396 vss n4108 cla_cell3_22_sp vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11395 vss cla_cell3_22_p11 n4113 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11394 n4113 cla_cell2_18_sp n4114 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11393 n4112 cla_cell2_22_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11392 n4111 cla_cell3_22_p11 n4112 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11391 vss cla_cell2_18_sg n4111 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11390 vss cla_cell2_26_sg n1891 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11389 n1891 cla_cell0_28_p cla_cell3_28_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11388 cla_cell3_28_g cla_cell3_28_g1 vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11387 n1889 cla_cell2_26_sp cla_cell4_28_pl vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11386 vss cla_cell0_28_p n1889 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11385 vss cla_cell2_26_sg n1122 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11384 n1122 cla_cell2_29_np cla_cell3_29_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11383 cla_cell3_29_g cla_cell2_29_ng vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11382 n1376 cla_cell2_26_sp cla_cell4_29_pl vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11381 vss cla_cell2_29_np n1376 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11380 vss cla_cell2_26_sg n1120 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11379 n1120 cla_cell3_30_p1 cla_cell3_30_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11378 cla_cell3_30_g cla_cell2_30_g vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11377 n1119 cla_cell2_26_sp cla_cell4_30_pl vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11376 vss cla_cell3_30_p1 n1119 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11375 vss cla_cell2_26_sg n600 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11374 n600 cla_cell3_31_p1 cla_cell3_31_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11373 cla_cell3_31_g cla_cell2_31_g vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_11372 n599 cla_cell2_26_sp cla_cell4_31_pl vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11371 vss cla_cell3_31_p1 n599 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11370 n9281 cla_cell1_8_np vss vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11369 n9281 cla_cell1_8_ng cla_cell7_8_g vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11368 vss cla_cell4_8_g2 n9281 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11367 n8785 cla_cell2_9_sp vss vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11366 n8785 cla_cell1_9_g cla_cell7_10_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11365 vss cla_cell4_8_g2 n8785 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11364 n8545 n8551 vss vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P PS=3.6U 
+ PD=3.6U 
Mtr_11363 n8545 cla_cell2_10_g1 cla_cell7_10_g vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11362 vss cla_cell4_8_g2 n8545 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11361 n8028 n8121 vss vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P PS=3.6U 
+ PD=3.6U 
Mtr_11360 n8028 cla_cell2_10_g2 cla_cell7_12_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11359 vss cla_cell4_8_g2 n8028 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11358 n7810 n7813 vss vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P PS=3.6U 
+ PD=3.6U 
Mtr_11357 n7810 cla_cell3_12_g cla_cell7_12_g vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11356 vss cla_cell4_8_g2 n7810 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11355 n7218 n7384 vss vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P PS=3.6U 
+ PD=3.6U 
Mtr_11354 n7218 cla_cell3_13_g cla_cell7_14_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11353 vss cla_cell4_8_g2 n7218 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11352 n7217 n7052 vss vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P PS=3.6U 
+ PD=3.6U 
Mtr_11351 n7217 cla_cell3_14_g cla_cell7_14_g vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11350 vss cla_cell4_8_g2 n7217 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11349 vss n6783 cla_cell5_16_g2 vss TN L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_11348 cla_cell5_16_g2 n6783 vss vss TN L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_11347 vss cla_cell4_15_p1 n6632 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11346 cla_cell4_8_g2 n6632 n6783 vss TN L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_11345 n6783 cla_cell4_15_p1 cla_cell3_15_g vss TN L=0.18U W=2.16U 
+ AS=0.7776P AD=0.7776P PS=5.04U PD=5.04U 
Mtr_11344 cla_cell4_20_ng cla_cell3_20_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11343 vss cla_cell4_20_p cla_cell4_20_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11342 cla_cell4_21_ng cla_cell3_21_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11341 vss cla_cell4_21_p cla_cell4_21_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11340 vss cla_cell3_22_sp cla_cell5_24_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11339 vss cla_cell1_24_np cla_cell5_24_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11338 n3526 cla_cell1_24_ng cla_cell4_24_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11337 vss cla_cell1_24_np n3526 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11336 n3526 cla_cell3_22_sg vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11335 vss cla_cell3_22_sp cla_cell5_25_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11334 vss cla_cell2_25_sp cla_cell5_25_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11333 n2716 cla_cell4_25_gl cla_cell4_25_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11332 vss cla_cell2_25_sp n2716 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11331 n2716 cla_cell3_22_sg vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11330 vss cla_cell3_22_sp cla_cell5_26_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11329 vss cla_cell4_26_pl cla_cell5_26_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11328 n2714 cla_cell2_26_g1 cla_cell4_26_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11327 vss cla_cell4_26_pl n2714 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11326 n2714 cla_cell3_22_sg vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11325 vss cla_cell3_22_sp cla_cell5_27_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11324 vss cla_cell4_27_pl cla_cell5_27_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11323 n2131 cla_cell4_27_gl cla_cell4_27_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11322 vss cla_cell4_27_pl n2131 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11321 n2131 cla_cell3_22_sg vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11320 vss cla_cell3_22_sp cla_cell5_28_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11319 vss cla_cell4_28_pl cla_cell5_28_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11318 n1886 cla_cell3_28_g cla_cell4_28_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11317 vss cla_cell4_28_pl n1886 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11316 n1886 cla_cell3_22_sg vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11315 vss cla_cell3_22_sp cla_cell5_29_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11314 vss cla_cell4_29_pl cla_cell5_29_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11313 n1375 cla_cell3_29_g cla_cell4_29_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11312 vss cla_cell4_29_pl n1375 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11311 n1375 cla_cell3_22_sg vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11310 vss cla_cell3_22_sp cla_cell5_30_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11309 vss cla_cell4_30_pl cla_cell5_30_p1 vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11308 n1117 cla_cell3_30_g cla_cell4_30_g vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11307 vss cla_cell4_30_pl n1117 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11306 n1117 cla_cell3_22_sg vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11305 vss cla_cell3_22_sp n678 vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11304 vss cla_cell4_31_pl n678 vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11303 n598 cla_cell3_31_g cla_cell4_31_g vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11302 vss cla_cell4_31_pl n598 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11301 n598 cla_cell3_22_sg vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_11300 vss cla_cell5_16_g2 n6408 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11299 n6408 cla_cell5_16_p1 cla_cell5_16_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11298 cla_cell5_16_co cla_cell1_16_sg vss vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11297 vss cla_cell5_16_g2 n5610 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11296 n5610 cla_cell2_17_np cla_cell5_17_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11295 cla_cell5_17_co cla_cell2_17_ng vss vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11294 vss cla_cell5_16_g2 n5608 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11293 n5608 cla_cell5_18_p1 cla_cell5_18_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11292 cla_cell5_18_co cla_cell2_18_g1 vss vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11291 vss cla_cell5_16_g2 n4857 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11290 n4857 cla_cell2_18_sp cla_cell5_19_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11289 cla_cell5_19_co cla_cell2_18_sg vss vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11288 vss cla_cell5_16_g2 n4856 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11287 n4856 cla_cell4_20_np cla_cell5_20_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11286 cla_cell5_20_co cla_cell4_20_ng vss vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11285 vss cla_cell5_16_g2 n4350 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11284 n4350 cla_cell4_21_np cla_cell5_21_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11283 cla_cell5_21_co cla_cell4_21_ng vss vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11282 vss cla_cell5_16_g2 n4104 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11281 n4104 cla_cell5_22_p1 cla_cell5_22_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11280 cla_cell5_22_co cla_cell3_22_g1 vss vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11279 vss cla_cell5_16_g2 n3525 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11278 n3525 cla_cell5_23_p1 cla_cell5_23_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11277 cla_cell5_23_co cla_cell3_22_g2 vss vss TN L=0.18U W=0.72U 
+ AS=0.2592P AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11276 vss cla_cell5_16_g2 n3524 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11275 n3524 cla_cell5_24_p1 cla_cell5_24_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11274 cla_cell5_24_co cla_cell4_24_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11273 vss cla_cell5_16_g2 n2713 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11272 n2713 cla_cell5_25_p1 cla_cell5_25_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11271 cla_cell5_25_co cla_cell4_25_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11270 vss cla_cell5_16_g2 n2712 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11269 n2712 cla_cell5_26_p1 cla_cell5_26_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11268 cla_cell5_26_co cla_cell4_26_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11267 vss cla_cell5_16_g2 n1884 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11266 n1884 cla_cell5_27_p1 cla_cell5_27_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11265 cla_cell5_27_co cla_cell4_27_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11264 vss cla_cell5_16_g2 n1882 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11263 n1882 cla_cell5_28_p1 cla_cell5_28_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11262 cla_cell5_28_co cla_cell4_28_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11261 vss cla_cell5_16_g2 n1114 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11260 n1114 cla_cell5_29_p1 cla_cell5_29_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11259 cla_cell5_29_co cla_cell4_29_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11258 vss cla_cell5_16_g2 n1112 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11257 n1112 cla_cell5_30_p1 cla_cell5_30_co vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11256 cla_cell5_30_co cla_cell4_30_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_11255 vss cla_cell5_16_g2 n597 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_11254 n597 n678 cla_cell5_31_co vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_11253 cla_cell5_31_co cla_cell4_31_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11252 n389 cla_cell1_32_np vss vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11251 n389 cla_cell1_32_ng cla_cell7_32_g vss TN L=0.18U W=1.44U 
+ AS=0.5184P AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11250 vss cla_cell5_31_co n389 vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_11249 n1 n39 vss vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P PS=3.6U 
+ PD=3.6U 
Mtr_11248 n1 cla_cell1_33_g n38 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11247 vss cla_cell5_31_co n1 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_11246 n11779 cla_cell0_0_g cla_cell0_1_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11245 n11779 cla_cell0_1_p cla_cell0_0_g vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11244 p_31 n11779 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11243 n11473 cla_cell0_2_pn cla_cell1_1_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11242 n11473 cla_cell1_1_co cla_cell0_2_pn vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11241 p_32 n11473 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11240 n11265 cla_cell7_2_g cla_cell1_3_p1 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11239 n11265 cla_cell1_3_p1 cla_cell7_2_g vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11238 p_33 n11265 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11237 n10887 cla_cell3_4_p1 cla_cell3_4_g2 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11236 n10887 cla_cell3_4_g2 cla_cell3_4_p1 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11235 p_34 n10887 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11234 n10453 cla_cell3_4_co cla_cell7_5_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11233 n10453 cla_cell7_5_p cla_cell3_4_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11232 p_35 n10453 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11231 n10061 cla_cell7_6_p cla_cell3_5_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11230 n10061 cla_cell3_5_co cla_cell7_6_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11229 p_36 n10061 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11228 n9619 cla_cell3_6_co cla_cell0_7_pn vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11227 n9619 cla_cell0_7_pn cla_cell3_6_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11226 p_37 n9619 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11225 n9280 cla_cell7_8_p cla_cell4_8_g2 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11224 n9280 cla_cell4_8_g2 cla_cell7_8_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11223 p_38 n9280 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11222 n8857 cla_cell7_8_g cla_cell0_9_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11221 n8857 cla_cell0_9_p cla_cell7_8_g vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11220 p_39 n8857 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11219 n8543 cla_cell0_10_p cla_cell7_10_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11218 n8543 cla_cell7_10_co cla_cell0_10_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11217 p_40 n8543 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11216 n8117 cla_cell7_10_g cla_cell0_11_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11215 n8117 cla_cell0_11_p cla_cell7_10_g vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11214 p_41 n8117 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11213 n7808 cla_cell0_12_p cla_cell7_12_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11212 n7808 cla_cell7_12_co cla_cell0_12_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11211 p_42 n7808 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11210 n7600 cla_cell7_12_g cla_cell0_13_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11209 n7600 cla_cell0_13_p cla_cell7_12_g vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11208 p_43 n7600 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11207 n7216 cla_cell0_14_p cla_cell7_14_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11206 n7216 cla_cell7_14_co cla_cell0_14_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11205 p_44 n7216 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11204 n6779 cla_cell7_14_g cla_cell1_15_p1 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11203 n6779 cla_cell1_15_p1 cla_cell7_14_g vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11202 p_45 n6779 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11201 n6405 cla_cell5_16_p1 cla_cell5_16_g2 vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11200 n6405 cla_cell5_16_g2 cla_cell5_16_p1 vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11199 p_46 n6405 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11198 n5938 cla_cell5_16_co cla_cell0_17_pn vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11197 n5938 cla_cell0_17_pn cla_cell5_16_co vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11196 p_47 n5938 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11195 n5606 cla_cell7_18_p cla_cell5_17_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11194 n5606 cla_cell5_17_co cla_cell7_18_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11193 p_48 n5606 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11192 n5165 cla_cell5_18_co cla_cell0_19_pn vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11191 n5165 cla_cell0_19_pn cla_cell5_18_co vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11190 p_49 n5165 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11189 n4854 cla_cell0_20_pn cla_cell5_19_co vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11188 n4854 cla_cell5_19_co cla_cell0_20_pn vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11187 p_50 n4854 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11186 n4425 cla_cell5_20_co cla_cell0_21_pn vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11185 n4425 cla_cell0_21_pn cla_cell5_20_co vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11184 p_51 n4425 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11183 n4102 cla_cell0_22_pn cla_cell5_21_co vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11182 n4102 cla_cell5_21_co cla_cell0_22_pn vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11181 p_52 n4102 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11180 n3671 cla_cell5_22_co cla_cell0_23_pn vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11179 n3671 cla_cell0_23_pn cla_cell5_22_co vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11178 p_53 n3671 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11177 n3523 cla_cell0_24_pn cla_cell5_23_co vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11176 n3523 cla_cell5_23_co cla_cell0_24_pn vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11175 p_54 n3523 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11174 n3082 cla_cell5_24_co cla_cell0_25_pn vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11173 n3082 cla_cell0_25_pn cla_cell5_24_co vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11172 p_55 n3082 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11171 n2710 cla_cell7_26_p cla_cell5_25_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11170 n2710 cla_cell5_25_co cla_cell7_26_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11169 p_56 n2710 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11168 n2247 cla_cell5_26_co cla_cell7_27_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11167 n2247 cla_cell7_27_p cla_cell5_26_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11166 p_57 n2247 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11165 n1880 cla_cell7_28_p cla_cell5_27_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11164 n1880 cla_cell5_27_co cla_cell7_28_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11163 p_58 n1880 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11162 n1432 cla_cell5_28_co cla_cell0_29_pn vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11161 n1432 cla_cell0_29_pn cla_cell5_28_co vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11160 p_59 n1432 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11159 n1111 cla_cell0_30_pn cla_cell5_29_co vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11158 n1111 cla_cell5_29_co cla_cell0_30_pn vss TN L=0.18U W=0.9U 
+ AS=0.324P AD=0.324P PS=2.52U PD=2.52U 
Mtr_11157 p_60 n1111 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11156 n673 cla_cell5_30_co cla_cell0_31_pn vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11155 n673 cla_cell0_31_pn cla_cell5_30_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11154 p_61 n673 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11153 n387 cla_cell0_32_pn cla_cell5_31_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11152 n387 cla_cell5_31_co cla_cell0_32_pn vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11151 p_62 n387 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11150 n36 cla_cell7_32_g cla_cell0_33_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11149 n36 cla_cell0_33_p cla_cell7_32_g vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11148 p_63 n36 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_11147 vss n55 cla_cell0_33_a vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_11146 n6 p_18_33_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11145 vss c_18_31_a n6 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_11144 n55 c_18_32_cin n6 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11143 n5 p_18_33_pi2j n55 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11142 vss c_18_31_a n5 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_11141 n51 c_18_32_cin n54 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11140 n54 n51 c_18_32_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11139 c_18_31_a p_18_33_pi2j n50 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11138 n50 c_18_31_a p_18_33_pi2j vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11137 cla_cell0_32_a n54 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_11136 vss n50 n51 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P PS=6.48U 
+ PD=6.48U 
Mtr_11135 n59 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11134 n61 a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_11133 vss p_18_33_t_s p_18_33_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11132 p_18_33_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11131 n61 n59 p_18_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11130 p_18_33_t_s n61 n59 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11129 n412 p_18_2_d2j n411 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11128 n408 p_18_2_d2jbar n412 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11127 p_18_32_t_s n412 n409 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11126 n412 n409 p_18_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11125 p_18_32_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11124 vss p_18_32_t_s p_18_32_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11123 n409 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11122 vss a_31 n408 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_11121 n411 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_11120 vss n402 c_18_32_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_11119 n401 c_18_31_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11118 vss p_18_32_pi2j n401 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11117 n402 c_18_32_cin n401 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11116 n400 c_18_31_a n402 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11115 vss p_18_32_pi2j n400 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11114 n404 c_18_32_cin c_18_32_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11113 c_18_32_s2_s n404 c_18_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11112 p_18_32_pi2j c_18_31_a c_18_32_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11111 c_18_32_s1_s p_18_32_pi2j c_18_31_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11110 c_18_32_sum c_18_32_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_11109 vss c_18_32_s1_s n404 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_11108 vss n707 c_18_31_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_11107 n606 p_18_31_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11106 vss c_18_31_a n606 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11105 n707 c_18_31_cin n606 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11104 n605 p_18_31_pi2j n707 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11103 vss c_18_31_a n605 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11102 n704 c_18_31_cin c_18_31_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11101 c_18_31_s2_s n704 c_18_31_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11100 c_18_31_a p_18_31_pi2j c_18_31_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11099 c_18_31_s1_s c_18_31_a p_18_31_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11098 c_18_31_sum c_18_31_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_11097 vss c_18_31_s1_s n704 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_11096 n713 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11095 vss a_29 n607 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_11094 n607 p_18_2_d2j n715 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11093 n715 p_18_2_d2jbar n608 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11092 n608 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_11091 vss p_18_31_t_s p_18_31_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11090 p_18_31_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11089 n715 n713 p_18_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11088 p_18_31_t_s n715 n713 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11087 n1150 p_18_2_d2j n1151 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11086 n1147 p_18_2_d2jbar n1150 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11085 p_18_30_t_s n1150 n1148 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11084 n1150 n1148 p_18_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11083 p_18_30_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11082 vss p_18_30_t_s p_18_30_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11081 n1148 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11080 vss a_29 n1147 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_11079 n1151 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_11078 vss n1140 c_18_30_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_11077 n1139 c_18_30_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11076 vss p_18_30_pi2j n1139 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11075 n1140 c_18_30_cin n1139 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11074 n1138 c_18_30_a n1140 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11073 vss p_18_30_pi2j n1138 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11072 n1142 c_18_30_cin c_18_30_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11071 c_18_30_s2_s n1142 c_18_30_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11070 p_18_30_pi2j c_18_30_a c_18_30_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11069 c_18_30_s1_s p_18_30_pi2j c_18_30_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11068 c_18_30_sum c_18_30_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_11067 vss c_18_30_s1_s n1142 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_11066 vss n1467 c_18_29_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_11065 n1379 p_18_29_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11064 vss c_18_29_a n1379 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11063 n1467 c_18_29_cin n1379 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11062 n1378 p_18_29_pi2j n1467 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11061 vss c_18_29_a n1378 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11060 n1462 c_18_29_cin c_18_29_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11059 c_18_29_s2_s n1462 c_18_29_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11058 c_18_29_a p_18_29_pi2j c_18_29_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11057 c_18_29_s1_s c_18_29_a p_18_29_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11056 c_18_29_sum c_18_29_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_11055 vss c_18_29_s1_s n1462 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_11054 n1473 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11053 vss a_27 n1380 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_11052 n1380 p_18_2_d2j n1475 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11051 n1475 p_18_2_d2jbar n1381 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11050 n1381 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_11049 vss p_18_29_t_s p_18_29_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11048 p_18_29_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11047 n1475 n1473 p_18_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11046 p_18_29_t_s n1475 n1473 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11045 n1913 p_18_2_d2j n1914 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11044 n1910 p_18_2_d2jbar n1913 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11043 p_18_28_t_s n1913 n1911 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11042 n1913 n1911 p_18_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11041 p_18_28_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11040 vss p_18_28_t_s p_18_28_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11039 n1911 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11038 vss a_27 n1910 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_11037 n1914 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_11036 vss n1902 c_18_28_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_11035 n1904 c_18_28_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11034 vss p_18_28_pi2j n1904 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11033 n1902 c_18_28_cin n1904 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11032 n1903 c_18_28_a n1902 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11031 vss p_18_28_pi2j n1903 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11030 n1774 c_18_28_cin c_18_28_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11029 c_18_28_s2_s n1774 c_18_28_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11028 p_18_28_pi2j c_18_28_a c_18_28_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11027 c_18_28_s1_s p_18_28_pi2j c_18_28_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11026 c_18_28_sum c_18_28_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_11025 vss c_18_28_s1_s n1774 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_11024 vss n2279 c_18_27_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_11023 n2134 c_18_27_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11022 vss c_18_27_a n2134 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11021 n2279 c_18_27_cin n2134 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11020 n1901 c_18_27_b n2279 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11019 vss c_18_27_a n1901 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_11018 n2272 c_18_27_cin c_18_27_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11017 c_18_27_s2_s n2272 c_18_27_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11016 c_18_27_a c_18_27_b c_18_27_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11015 c_18_27_s1_s c_18_27_a c_18_27_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_11014 c_18_27_sum c_18_27_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_11013 vss c_18_27_s1_s n2272 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_11012 n2283 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11011 vss a_25 n2138 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_11010 n2138 p_18_2_d2j n2280 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11009 n2280 p_18_2_d2jbar n2140 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11008 n2140 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_11007 vss p_18_27_t_s c_18_27_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11006 c_18_27_b p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_11005 n2280 n2283 p_18_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11004 p_18_27_t_s n2280 n2283 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11003 n2595 p_18_2_d2j n2594 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11002 n2592 p_18_2_d2jbar n2595 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_11001 p_18_26_t_s n2595 n2593 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_11000 n2595 n2593 p_18_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10999 p_18_26_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10998 vss p_18_26_t_s p_18_26_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10997 n2593 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10996 vss a_25 n2592 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10995 n2594 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10994 vss n2736 c_18_26_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10993 n2738 c_18_26_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10992 vss p_18_26_pi2j n2738 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10991 n2736 c_18_26_cin n2738 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10990 n2737 c_18_26_a n2736 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10989 vss p_18_26_pi2j n2737 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10988 n2591 c_18_26_cin c_18_26_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10987 c_18_26_s2_s n2591 c_18_26_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10986 p_18_26_pi2j c_18_26_a c_18_26_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10985 c_18_26_s1_s p_18_26_pi2j c_18_26_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10984 c_18_26_sum c_18_26_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10983 vss c_18_26_s1_s n2591 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10982 vss n3107 c_18_25_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10981 n2735 c_18_25_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10980 vss c_18_25_a n2735 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10979 n3107 c_18_25_cin n2735 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10978 n2734 c_18_25_b n3107 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10977 vss c_18_25_a n2734 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10976 n2939 c_18_25_cin c_18_25_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10975 c_18_25_s2_s n2939 c_18_25_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10974 c_18_25_a c_18_25_b c_18_25_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10973 c_18_25_s1_s c_18_25_a c_18_25_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10972 c_18_25_sum c_18_25_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10971 vss c_18_25_s1_s n2939 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10970 n3112 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10969 vss a_23 n2744 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10968 n2744 p_18_2_d2j n2944 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10967 n2944 p_18_2_d2jbar n2745 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10966 n2745 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10965 vss p_18_25_t_s c_18_25_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10964 c_18_25_b p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10963 n2944 n3112 p_18_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10962 p_18_25_t_s n2944 n3112 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10961 n3362 p_18_2_d2j n3363 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10960 n3360 p_18_2_d2jbar n3362 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10959 p_18_24_t_s n3362 n3361 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10958 n3362 n3361 p_18_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10957 c_18_24_b p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10956 vss p_18_24_t_s c_18_24_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10955 n3361 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10954 vss a_23 n3360 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10953 n3363 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10952 vss n3353 c_18_24_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10951 n3538 c_18_24_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10950 vss c_18_24_b n3538 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10949 n3353 c_18_24_cin n3538 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10948 n3539 c_18_24_a n3353 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10947 vss c_18_24_b n3539 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10946 n3356 c_18_24_cin c_18_24_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10945 c_18_24_s2_s n3356 c_18_24_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10944 c_18_24_b c_18_24_a c_18_24_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10943 c_18_24_s1_s c_18_24_b c_18_24_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10942 c_18_24_sum c_18_24_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10941 vss c_18_24_s1_s n3356 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10940 vss n3697 c_18_23_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10939 n3537 c_18_23_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10938 vss c_18_23_a n3537 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10937 n3697 c_18_23_cin n3537 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10936 n3536 c_18_23_b n3697 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10935 vss c_18_23_a n3536 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10934 n3699 c_18_23_cin c_18_23_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10933 c_18_23_s2_s n3699 c_18_23_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10932 c_18_23_a c_18_23_b c_18_23_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10931 c_18_23_s1_s c_18_23_a c_18_23_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10930 c_18_23_sum c_18_23_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10929 vss c_18_23_s1_s n3699 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10928 n3703 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10927 vss a_21 n3542 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10926 n3542 p_18_2_d2j n3705 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10925 n3705 p_18_2_d2jbar n3544 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10924 n3544 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10923 vss p_18_23_t_s c_18_23_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10922 c_18_23_b p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10921 n3705 n3703 p_18_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10920 p_18_23_t_s n3705 n3703 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10919 n4141 p_18_2_d2j n4140 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10918 n4138 p_18_2_d2jbar n4141 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10917 p_18_22_t_s n4141 n4139 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10916 n4141 n4139 p_18_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10915 p_18_22_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10914 vss p_18_22_t_s p_18_22_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10913 n4139 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10912 vss a_21 n4138 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10911 n4140 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10910 vss n4130 c_18_22_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10909 n4129 c_18_22_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10908 vss p_18_22_pi2j n4129 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10907 n4130 c_18_22_cin n4129 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10906 n4128 c_18_22_a n4130 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10905 vss p_18_22_pi2j n4128 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10904 n4132 c_18_22_cin c_18_22_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10903 c_18_22_s2_s n4132 c_18_22_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10902 p_18_22_pi2j c_18_22_a c_18_22_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10901 c_18_22_s1_s p_18_22_pi2j c_18_22_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10900 c_18_22_sum c_18_22_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10899 vss c_18_22_s1_s n4132 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10898 vss n4453 c_18_21_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10897 n4357 p_18_21_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10896 vss c_18_21_a n4357 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10895 n4453 c_18_21_cin n4357 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10894 n4356 p_18_21_pi2j n4453 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10893 vss c_18_21_a n4356 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10892 n4449 c_18_21_cin c_18_21_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10891 c_18_21_s2_s n4449 c_18_21_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10890 c_18_21_a p_18_21_pi2j c_18_21_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10889 c_18_21_s1_s c_18_21_a p_18_21_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10888 c_18_21_sum c_18_21_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10887 vss c_18_21_s1_s n4449 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10886 n4460 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10885 vss a_19 n4358 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10884 n4358 p_18_2_d2j n4462 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10883 n4462 p_18_2_d2jbar n4359 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10882 n4359 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10881 vss p_18_21_t_s p_18_21_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10880 p_18_21_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10879 n4462 n4460 p_18_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10878 p_18_21_t_s n4462 n4460 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10877 n4886 p_18_2_d2j n4887 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10876 n4884 p_18_2_d2jbar n4886 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10875 p_18_20_t_s n4886 n4885 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10874 n4886 n4885 p_18_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10873 p_18_20_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10872 vss p_18_20_t_s p_18_20_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10871 n4885 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10870 vss a_19 n4884 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10869 n4887 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10868 vss n4876 c_18_20_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10867 n4875 c_18_20_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10866 vss p_18_20_pi2j n4875 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10865 n4876 c_18_20_cin n4875 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10864 n4874 c_18_20_a n4876 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10863 vss p_18_20_pi2j n4874 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10862 n4878 c_18_20_cin c_18_20_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10861 c_18_20_s2_s n4878 c_18_20_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10860 p_18_20_pi2j c_18_20_a c_18_20_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10859 c_18_20_s1_s p_18_20_pi2j c_18_20_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10858 c_18_20_sum c_18_20_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10857 vss c_18_20_s1_s n4878 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10856 vss n5193 c_18_19_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10855 n5097 p_18_19_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10854 vss c_18_19_a n5097 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10853 n5193 c_18_19_cin n5097 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10852 n5098 p_18_19_pi2j n5193 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10851 vss c_18_19_a n5098 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10850 n5189 c_18_19_cin c_18_19_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10849 c_18_19_s2_s n5189 c_18_19_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10848 c_18_19_a p_18_19_pi2j c_18_19_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10847 c_18_19_s1_s c_18_19_a p_18_19_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10846 c_18_19_sum c_18_19_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10845 vss c_18_19_s1_s n5189 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10844 n5200 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10843 vss a_17 n5099 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10842 n5099 p_18_2_d2j n5203 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10841 n5203 p_18_2_d2jbar n5100 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10840 n5100 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10839 vss p_18_19_t_s p_18_19_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10838 p_18_19_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10837 n5203 n5200 p_18_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10836 p_18_19_t_s n5203 n5200 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10835 n5640 p_18_2_d2j n5639 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10834 n5636 p_18_2_d2jbar n5640 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10833 p_18_18_t_s n5640 n5637 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10832 n5640 n5637 p_18_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10831 p_18_18_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10830 vss p_18_18_t_s p_18_18_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10829 n5637 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10828 vss a_17 n5636 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10827 n5639 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10826 vss n5628 c_18_18_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10825 n5630 c_18_18_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10824 vss p_18_18_pi2j n5630 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10823 n5628 c_18_18_cin n5630 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10822 n5629 c_18_18_a n5628 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10821 vss p_18_18_pi2j n5629 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10820 n5500 c_18_18_cin c_18_18_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10819 c_18_18_s2_s n5500 c_18_18_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10818 p_18_18_pi2j c_18_18_a c_18_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10817 c_18_18_s1_s p_18_18_pi2j c_18_18_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10816 c_18_18_sum c_18_18_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10815 vss c_18_18_s1_s n5500 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10814 vss n5964 c_18_17_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10813 n5857 p_18_17_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10812 vss c_18_17_a n5857 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10811 n5964 c_18_17_cin n5857 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10810 n5627 p_18_17_pi2j n5964 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10809 vss c_18_17_a n5627 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10808 n5958 c_18_17_cin c_18_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10807 c_18_17_s2_s n5958 c_18_17_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10806 c_18_17_a p_18_17_pi2j c_18_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10805 c_18_17_s1_s c_18_17_a p_18_17_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10804 c_18_17_sum c_18_17_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10803 vss c_18_17_s1_s n5958 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10802 n5972 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10801 vss a_15 n5859 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10800 n5859 p_18_2_d2j n5968 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10799 n5968 p_18_2_d2jbar n5861 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10798 n5861 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10797 vss p_18_17_t_s p_18_17_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10796 p_18_17_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10795 n5968 n5972 p_18_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10794 p_18_17_t_s n5968 n5972 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10793 n6305 p_18_2_d2j n6304 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10792 n6303 p_18_2_d2jbar n6305 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10791 p_18_16_t_s n6305 n6429 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10790 n6305 n6429 p_18_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10789 p_18_16_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10788 vss p_18_16_t_s p_18_16_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10787 n6429 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10786 vss a_15 n6303 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10785 n6304 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10784 vss n6423 c_18_16_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10783 n6422 c_18_16_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10782 vss p_18_16_pi2j n6422 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10781 n6423 c_18_16_cin n6422 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10780 n6421 c_18_16_a n6423 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10779 vss p_18_16_pi2j n6421 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10778 n6302 c_18_16_cin c_18_16_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10777 c_18_16_s2_s n6302 c_18_16_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10776 p_18_16_pi2j c_18_16_a c_18_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10775 c_18_16_s1_s p_18_16_pi2j c_18_16_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10774 c_18_16_sum c_18_16_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10773 vss c_18_16_s1_s n6302 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10772 vss n6810 c_18_15_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10771 n6637 c_18_15_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10770 vss c_18_15_a n6637 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10769 n6810 c_18_15_cin n6637 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10768 n6420 c_18_15_b n6810 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10767 vss c_18_15_a n6420 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10766 n6640 c_18_15_cin c_18_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10765 c_18_15_s2_s n6640 c_18_15_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10764 c_18_15_a c_18_15_b c_18_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10763 c_18_15_s1_s c_18_15_a c_18_15_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10762 c_18_15_sum c_18_15_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10761 vss c_18_15_s1_s n6640 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10760 n6814 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10759 vss a_13 n6430 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10758 n6430 p_18_2_d2j n6645 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10757 n6645 p_18_2_d2jbar n6431 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10756 n6431 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10755 vss p_18_15_t_s c_18_15_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10754 c_18_15_b p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10753 n6645 n6814 p_18_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10752 p_18_15_t_s n6645 n6814 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10751 n7069 p_18_2_d2j n7070 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10750 n7067 p_18_2_d2jbar n7069 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10749 p_18_14_t_s n7069 n7068 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10748 n7069 n7068 p_18_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10747 p_18_14_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10746 vss p_18_14_t_s p_18_14_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10745 n7068 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10744 vss a_13 n7067 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10743 n7070 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10742 vss n7061 c_18_14_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10741 n7234 c_18_14_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10740 vss p_18_14_pi2j n7234 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10739 n7061 c_18_14_cin n7234 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10738 n7235 c_18_14_a n7061 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10737 vss p_18_14_pi2j n7235 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10736 n7064 c_18_14_cin c_18_14_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10735 c_18_14_s2_s n7064 c_18_14_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10734 p_18_14_pi2j c_18_14_a c_18_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10733 c_18_14_s1_s p_18_14_pi2j c_18_14_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10732 c_18_14_sum c_18_14_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10731 vss c_18_14_s1_s n7064 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10730 vss n7397 c_18_13_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10729 n7233 c_18_13_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10728 vss c_18_13_a n7233 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10727 n7397 c_18_13_cin n7233 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10726 n7232 c_18_13_b n7397 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10725 vss c_18_13_a n7232 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10724 n7400 c_18_13_cin c_18_13_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10723 c_18_13_s2_s n7400 c_18_13_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10722 c_18_13_a c_18_13_b c_18_13_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10721 c_18_13_s1_s c_18_13_a c_18_13_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10720 c_18_13_sum c_18_13_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10719 vss c_18_13_s1_s n7400 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10718 n7404 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10717 vss a_11 n7239 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10716 n7239 p_18_2_d2j n7406 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10715 n7406 p_18_2_d2jbar n7240 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10714 n7240 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10713 vss p_18_13_t_s c_18_13_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10712 c_18_13_b p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10711 n7406 n7404 p_18_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10710 p_18_13_t_s n7406 n7404 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10709 n7834 p_18_2_d2j n7833 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10708 n7831 p_18_2_d2jbar n7834 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10707 p_18_12_t_s n7834 n7832 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10706 n7834 n7832 p_18_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10705 c_18_12_b p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10704 vss p_18_12_t_s c_18_12_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10703 n7832 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10702 vss a_11 n7831 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10701 n7833 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10700 vss n7824 c_18_12_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10699 n7823 c_18_12_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10698 vss c_18_12_b n7823 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10697 n7824 c_18_12_cin n7823 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10696 n7822 c_18_12_a n7824 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10695 vss c_18_12_b n7822 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10694 n7826 c_18_12_cin c_18_12_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10693 c_18_12_s2_s n7826 c_18_12_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10692 c_18_12_b c_18_12_a c_18_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10691 c_18_12_s1_s c_18_12_b c_18_12_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10690 c_18_12_sum c_18_12_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10689 vss c_18_12_s1_s n7826 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10688 vss n8142 c_18_11_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10687 n8033 p_18_11_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10686 vss c_18_11_a n8033 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10685 n8142 c_18_11_cin n8033 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10684 n8032 p_18_11_pi2j n8142 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10683 vss c_18_11_a n8032 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10682 n8137 c_18_11_cin c_18_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10681 c_18_11_s2_s n8137 c_18_11_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10680 c_18_11_a p_18_11_pi2j c_18_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10679 c_18_11_s1_s c_18_11_a p_18_11_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10678 c_18_11_sum c_18_11_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10677 vss c_18_11_s1_s n8137 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10676 n8148 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10675 vss a_9 n8035 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10674 n8035 p_18_2_d2j n8150 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10673 n8150 p_18_2_d2jbar n8036 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10672 n8036 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10671 vss p_18_11_t_s p_18_11_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10670 p_18_11_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10669 n8150 n8148 p_18_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10668 p_18_11_t_s n8150 n8148 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10667 n8575 p_18_2_d2j n8576 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10666 n8573 p_18_2_d2jbar n8575 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10665 p_18_10_t_s n8575 n8574 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10664 n8575 n8574 p_18_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10663 p_18_10_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10662 vss p_18_10_t_s p_18_10_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10661 n8574 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10660 vss a_9 n8573 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10659 n8576 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10658 vss n8562 c_18_10_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10657 n8565 c_18_10_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10656 vss p_18_10_pi2j n8565 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10655 n8562 c_18_10_cin n8565 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10654 n8564 c_18_10_a n8562 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10653 vss p_18_10_pi2j n8564 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10652 n8567 c_18_10_cin c_18_10_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10651 c_18_10_s2_s n8567 c_18_10_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10650 p_18_10_pi2j c_18_10_a c_18_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10649 c_18_10_s1_s p_18_10_pi2j c_18_10_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10648 c_18_10_sum c_18_10_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_10647 vss c_18_10_s1_s n8567 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10646 vss n8882 c_18_9_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10645 n8790 p_18_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10644 vss c_18_9_a n8790 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10643 n8882 c_18_9_cin n8790 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10642 n8789 p_18_9_pi2j n8882 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10641 vss c_18_9_a n8789 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10640 n8877 c_18_9_cin c_18_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10639 c_18_9_s2_s n8877 c_18_9_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10638 c_18_9_a p_18_9_pi2j c_18_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10637 c_18_9_s1_s c_18_9_a p_18_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10636 c_18_9_sum c_18_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10635 vss c_18_9_s1_s n8877 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10634 n8888 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10633 vss a_7 n8791 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10632 n8791 p_18_2_d2j n8891 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10631 n8891 p_18_2_d2jbar n8792 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10630 n8792 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10629 vss p_18_9_t_s p_18_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10628 p_18_9_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10627 n8891 n8888 p_18_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10626 p_18_9_t_s n8891 n8888 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10625 n9308 p_18_2_d2j n9307 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10624 n9304 p_18_2_d2jbar n9308 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10623 p_18_8_t_s n9308 n9305 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10622 n9308 n9305 p_18_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10621 p_18_8_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10620 vss p_18_8_t_s p_18_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10619 n9305 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10618 vss a_7 n9304 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10617 n9307 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10616 vss n9296 c_18_8_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10615 n9297 c_18_8_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10614 vss p_18_8_pi2j n9297 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10613 n9296 c_18_8_cin n9297 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10612 n9298 c_18_8_a n9296 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10611 vss p_18_8_pi2j n9298 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10610 n9294 c_18_8_cin c_18_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10609 c_18_8_s2_s n9294 c_18_8_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10608 p_18_8_pi2j c_18_8_a c_18_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10607 c_18_8_s1_s p_18_8_pi2j c_18_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10606 c_18_8_sum c_18_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10605 vss c_18_8_s1_s n9294 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10604 vss n9651 c_18_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10603 n9535 p_18_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10602 vss c_18_7_a n9535 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10601 n9651 c_18_7_cin n9535 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10600 n9295 p_18_7_pi2j n9651 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10599 vss c_18_7_a n9295 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10598 n9646 c_18_7_cin c_18_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10597 c_18_7_s2_s n9646 c_18_7_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10596 c_18_7_a p_18_7_pi2j c_18_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10595 c_18_7_s1_s c_18_7_a p_18_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10594 c_18_7_sum c_18_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10593 vss c_18_7_s1_s n9646 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10592 n9656 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10591 vss a_5 n9537 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10590 n9537 p_18_2_d2j n9652 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10589 n9652 p_18_2_d2jbar n9539 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10588 n9539 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10587 vss p_18_7_t_s p_18_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10586 p_18_7_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10585 n9652 n9656 p_18_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10584 p_18_7_t_s n9652 n9656 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10583 n10090 p_18_2_d2j n9989 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10582 n9988 p_18_2_d2jbar n10090 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10581 p_18_6_t_s n10090 n10091 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10580 n10090 n10091 p_18_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10579 p_18_6_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10578 vss p_18_6_t_s p_18_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10577 n10091 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10576 vss a_5 n9988 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10575 n9989 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10574 vss n10084 c_18_6_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10573 n10083 c_18_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10572 vss p_18_6_pi2j n10083 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10571 n10084 c_18_6_cin n10083 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10570 n10082 c_18_6_a n10084 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10569 vss p_18_6_pi2j n10082 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10568 n9987 c_18_6_cin c_18_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10567 c_18_6_s2_s n9987 c_18_6_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10566 p_18_6_pi2j c_18_6_a c_18_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10565 c_18_6_s1_s p_18_6_pi2j c_18_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10564 c_18_6_sum c_18_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10563 vss c_18_6_s1_s n9987 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10562 vss n10475 c_18_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10561 n10312 c_18_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10560 vss c_18_5_a n10312 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10559 n10475 c_18_5_cin n10312 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10558 n10081 c_18_5_b n10475 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10557 vss c_18_5_a n10081 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10556 n10315 c_18_5_cin c_18_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10555 c_18_5_s2_s n10315 c_18_5_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10554 c_18_5_a c_18_5_b c_18_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10553 c_18_5_s1_s c_18_5_a c_18_5_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10552 c_18_5_sum c_18_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10551 vss c_18_5_s1_s n10315 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10550 n10481 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10549 vss a_3 n10092 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10548 n10092 p_18_2_d2j n10477 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10547 n10477 p_18_2_d2jbar n10093 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10546 n10093 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10545 vss p_18_5_t_s c_18_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_10544 c_18_5_b p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_10543 n10477 n10481 p_18_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10542 p_18_5_t_s n10477 n10481 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10541 n10744 p_18_2_d2j n10743 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10540 n10741 p_18_2_d2jbar n10744 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10539 p_18_4_t_s n10744 n10742 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10538 n10744 n10742 p_18_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10537 p_18_4_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10536 vss p_18_4_t_s p_18_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10535 n10742 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10534 vss a_3 n10741 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10533 n10743 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10532 vss n10735 c_18_4_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10531 n10902 c_18_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10530 vss p_18_4_pi2j n10902 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10529 n10735 c_18_4_cin n10902 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10528 n10903 c_18_4_a n10735 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10527 vss p_18_4_pi2j n10903 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10526 n10738 c_18_4_cin c_18_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10525 c_18_4_s2_s n10738 c_18_4_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10524 p_18_4_pi2j c_18_4_a c_18_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10523 c_18_4_s1_s p_18_4_pi2j c_18_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10522 c_18_4_sum c_18_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10521 vss c_18_4_s1_s n10738 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10520 vss n11062 c_18_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10519 n10901 c_18_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10518 vss c_18_3_a n10901 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10517 n11062 c_18_3_cin n10901 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10516 n10900 c_18_3_b n11062 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10515 vss c_18_3_a n10900 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10514 n11064 c_18_3_cin c_18_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10513 c_18_3_s2_s n11064 c_18_3_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10512 c_18_3_a c_18_3_b c_18_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10511 c_18_3_s1_s c_18_3_a c_18_3_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10510 c_18_3_sum c_18_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10509 vss c_18_3_s1_s n11064 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10508 n11069 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10507 vss a_1 n10907 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10506 n10907 p_18_2_d2j n11071 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10505 n11071 p_18_2_d2jbar n10908 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10504 n10908 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10503 vss p_18_3_t_s c_18_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_10502 c_18_3_b p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_10501 n11071 n11069 p_18_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10500 p_18_3_t_s n11071 n11069 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10499 n11496 p_18_2_d2j n11497 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10498 n11494 p_18_2_d2jbar n11496 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10497 p_18_2_t_s n11496 n11495 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10496 n11496 n11495 p_18_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10495 c_18_2_b p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_10494 vss p_18_2_t_s c_18_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_10493 n11495 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10492 vss a_1 n11494 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10491 n11497 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10490 vss n11487 c_18_2_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10489 n11486 c_18_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10488 vss c_18_2_b n11486 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10487 n11487 c_18_2_cin n11486 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10486 n11485 c_18_2_a n11487 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10485 vss c_18_2_b n11485 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10484 n11489 c_18_2_cin c_18_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10483 c_18_2_s2_s n11489 c_18_2_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10482 c_18_2_b c_18_2_a c_18_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10481 c_18_2_s1_s c_18_2_b c_18_2_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10480 c_18_2_sum c_18_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10479 vss c_18_2_s1_s n11489 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10478 vss n11796 c_18_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10477 n11695 p_18_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10476 vss c_18_1_a n11695 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10475 n11796 c_18_1_cin n11695 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10474 n11694 p_18_1_pi2j n11796 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10473 vss c_18_1_a n11694 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10472 n11792 c_18_1_cin c_18_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10471 c_18_1_s2_s n11792 c_18_1_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10470 c_18_1_a p_18_1_pi2j c_18_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10469 c_18_1_s1_s c_18_1_a p_18_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10468 c_18_1_sum c_18_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10467 vss c_18_1_s1_s n11792 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10466 n11805 p_18_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10465 n11806 p_18_2_d2jbar n11698 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10464 n11698 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10463 vss p_18_1_t_s p_18_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10462 p_18_1_pi2j p_18_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10461 n11806 n11805 p_18_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10460 p_18_1_t_s n11806 n11805 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10459 cl4_18_s1_s n12187 c_17_1_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10458 n12187 c_17_1_sum cl4_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10457 vss cl4_18_s1_s p_28 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_10456 vss c_17_1_sum n12177 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10455 n12177 n12187 n12176 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10454 n12175 n12176 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_10453 n12173 c_17_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_10452 vss c_17_2_sum n12173 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_10451 n12170 c_17_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10450 n12172 c_17_1_cout n12170 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10449 n12171 c_17_1_sum n12172 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10448 n12173 n12187 n12171 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10447 cla_cell0_0_a n12172 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10446 cl4_18_s2_s c_17_1_cout c_17_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10445 c_17_1_cout c_17_2_sum cl4_18_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10444 vss cl4_18_s2_s n12167 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10443 cl4_18_s3_s n12167 n12175 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10442 n12167 n12175 cl4_18_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10441 vss cl4_18_s3_s p_29 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_10440 vss c_17_33_s1_s n65 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10439 c_18_31_a c_17_33_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10438 c_17_33_s1_s c_17_31_a p_17_33_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10437 c_17_31_a p_17_33_pi2j c_17_33_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10436 c_17_33_s2_s n65 c_17_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10435 n65 c_17_32_cin c_17_33_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10434 vss c_17_31_a n8 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_10433 n8 p_17_33_pi2j n64 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10432 n64 c_17_32_cin n7 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10431 vss c_17_31_a n7 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_10430 n7 p_17_33_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10429 vss n64 c_18_32_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10428 n74 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10427 n75 a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10426 vss p_17_33_t_s p_17_33_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10425 p_17_33_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10424 n75 n74 p_17_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10423 p_17_33_t_s n75 n74 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10422 n424 p_17_2_d2j n427 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10421 n423 p_17_2_d2jbar n424 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10420 p_17_32_t_s n424 n422 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10419 n424 n422 p_17_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10418 p_17_32_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10417 vss p_17_32_t_s p_17_32_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10416 n422 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10415 vss a_31 n423 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10414 n427 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10413 vss c_17_32_s1_s n418 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10412 c_18_30_a c_17_32_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10411 c_17_32_s1_s p_17_32_pi2j c_17_31_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10410 c_17_32_s2_s n418 c_17_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10409 n418 c_17_32_cin c_17_32_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10408 vss p_17_32_pi2j n415 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10407 n415 c_17_31_a n414 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10406 n414 c_17_32_cin n413 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10405 vss p_17_32_pi2j n413 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10404 n413 c_17_31_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10403 vss n414 c_18_31_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10402 p_17_32_pi2j c_17_31_a c_17_32_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10401 vss n726 c_18_30_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10400 n610 p_17_31_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10399 vss c_17_31_a n610 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10398 n726 c_17_31_cin n610 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10397 n609 p_17_31_pi2j n726 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10396 vss c_17_31_a n609 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10395 n722 c_17_31_cin c_17_31_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10394 c_17_31_s2_s n722 c_17_31_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10393 c_17_31_a p_17_31_pi2j c_17_31_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10392 c_17_31_s1_s c_17_31_a p_17_31_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10391 c_18_29_a c_17_31_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10390 vss c_17_31_s1_s n722 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10389 n732 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10388 vss a_29 n611 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10387 n611 p_17_2_d2j n731 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10386 n731 p_17_2_d2jbar n613 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10385 n613 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10384 vss p_17_31_t_s p_17_31_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10383 p_17_31_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10382 n731 n732 p_17_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10381 p_17_31_t_s n731 n732 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10380 n1165 p_17_2_d2j n1169 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10379 n1164 p_17_2_d2jbar n1165 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10378 p_17_30_t_s n1165 n1163 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10377 n1165 n1163 p_17_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10376 p_17_30_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10375 vss p_17_30_t_s p_17_30_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10374 n1163 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10373 vss a_29 n1164 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10372 n1169 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10371 vss c_17_30_s1_s n1160 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10370 c_18_28_a c_17_30_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10369 c_17_30_s1_s p_17_30_pi2j c_17_30_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10368 c_17_30_s2_s n1160 c_16_31_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10367 n1160 c_16_31_cout c_17_30_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10366 vss p_17_30_pi2j n1153 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10365 n1153 c_17_30_a n1155 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10364 n1155 c_16_31_cout n1154 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10363 vss p_17_30_pi2j n1154 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10362 n1154 c_17_30_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10361 vss n1155 c_18_29_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10360 p_17_30_pi2j c_17_30_a c_17_30_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10359 vss n1488 c_18_28_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10358 n1382 p_17_29_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10357 vss c_17_29_a n1382 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10356 n1488 c_17_29_cin n1382 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10355 n1152 p_17_29_pi2j n1488 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10354 vss c_17_29_a n1152 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10353 n1484 c_17_29_cin c_17_29_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10352 c_17_29_s2_s n1484 c_17_29_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10351 c_17_29_a p_17_29_pi2j c_17_29_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10350 c_17_29_s1_s c_17_29_a p_17_29_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10349 c_18_27_a c_17_29_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10348 vss c_17_29_s1_s n1484 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10347 n1495 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10346 vss a_27 n1383 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10345 n1383 p_17_2_d2j n1493 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10344 n1493 p_17_2_d2jbar n1384 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10343 n1384 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10342 vss p_17_29_t_s p_17_29_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10341 p_17_29_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10340 n1493 n1495 p_17_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10339 p_17_29_t_s n1493 n1495 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10338 n1927 p_17_2_d2j n1931 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10337 n1926 p_17_2_d2jbar n1927 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10336 p_17_28_t_s n1927 n1925 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10335 n1927 n1925 p_17_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10334 p_17_28_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10333 vss p_17_28_t_s p_17_28_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10332 n1925 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10331 vss a_27 n1926 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10330 n1931 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10329 vss c_17_28_s1_s n1781 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10328 c_18_26_a c_17_28_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10327 c_17_28_s1_s p_17_28_pi2j c_17_28_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10326 c_17_28_s2_s n1781 c_16_29_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10325 n1781 c_16_29_cout c_17_28_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10324 vss p_17_28_pi2j n1917 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10323 n1917 c_17_28_a n1918 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10322 n1918 c_16_29_cout n1916 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10321 vss p_17_28_pi2j n1916 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10320 n1916 c_17_28_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10319 vss n1918 c_18_27_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10318 p_17_28_pi2j c_17_28_a c_17_28_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10317 vss n2300 c_18_26_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10316 n2141 c_17_27_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10315 vss c_17_27_a n2141 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10314 n2300 c_17_27_cin n2141 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10313 n1915 c_17_27_b n2300 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10312 vss c_17_27_a n1915 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10311 n2291 c_17_27_cin c_17_27_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10310 c_17_27_s2_s n2291 c_17_27_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10309 c_17_27_a c_17_27_b c_17_27_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10308 c_17_27_s1_s c_17_27_a c_17_27_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10307 c_18_25_a c_17_27_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10306 vss c_17_27_s1_s n2291 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10305 n2305 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10304 vss a_25 n2145 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10303 n2145 p_17_2_d2j n2301 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10302 n2301 p_17_2_d2jbar n2147 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10301 n2147 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10300 vss p_17_27_t_s c_17_27_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10299 c_17_27_b p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10298 n2301 n2305 p_17_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10297 p_17_27_t_s n2301 n2305 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10296 n2601 p_17_2_d2j n2603 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10295 n2602 p_17_2_d2jbar n2601 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10294 p_17_26_t_s n2601 n2600 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10293 n2601 n2600 p_17_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10292 p_17_26_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10291 vss p_17_26_t_s p_17_26_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10290 n2600 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10289 vss a_25 n2602 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10288 n2603 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10287 vss c_17_26_s1_s n2599 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10286 c_18_24_a c_17_26_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10285 c_17_26_s1_s p_17_26_pi2j c_17_26_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10284 c_17_26_s2_s n2599 c_16_27_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10283 n2599 c_16_27_cout c_17_26_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10282 vss p_17_26_pi2j n2750 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10281 n2750 c_17_26_a n2749 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10280 n2749 c_16_27_cout n2746 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10279 vss p_17_26_pi2j n2746 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10278 n2746 c_17_26_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10277 vss n2749 c_18_25_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10276 p_17_26_pi2j c_17_26_a c_17_26_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10275 vss n3123 c_18_24_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10274 n2748 c_17_25_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10273 vss c_17_25_a n2748 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10272 n3123 c_17_25_cin n2748 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10271 n2747 c_17_25_b n3123 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10270 vss c_17_25_a n2747 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10269 n2949 c_17_25_cin c_17_25_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10268 c_17_25_s2_s n2949 c_17_25_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10267 c_17_25_a c_17_25_b c_17_25_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10266 c_17_25_s1_s c_17_25_a c_17_25_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10265 c_18_23_a c_17_25_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10264 vss c_17_25_s1_s n2949 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10263 n3128 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10262 vss a_23 n2756 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10261 n2756 p_17_2_d2j n2952 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10260 n2952 p_17_2_d2jbar n2761 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10259 n2761 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10258 vss p_17_25_t_s c_17_25_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10257 c_17_25_b p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10256 n2952 n3128 p_17_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10255 p_17_25_t_s n2952 n3128 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10254 n3372 p_17_2_d2j n3374 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10253 n3373 p_17_2_d2jbar n3372 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10252 p_17_24_t_s n3372 n3371 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10251 n3372 n3371 p_17_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10250 c_17_24_b p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10249 vss p_17_24_t_s c_17_24_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10248 n3371 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10247 vss a_23 n3373 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10246 n3374 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10245 vss c_17_24_s1_s n3368 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10244 c_18_22_a c_17_24_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10243 c_17_24_s1_s c_17_24_b c_17_24_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10242 c_17_24_s2_s n3368 c_16_25_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10241 n3368 c_16_25_cout c_17_24_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10240 vss c_17_24_b n3547 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10239 n3547 c_17_24_a n3364 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10238 n3364 c_16_25_cout n3543 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10237 vss c_17_24_b n3543 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10236 n3543 c_17_24_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10235 vss n3364 c_18_23_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10234 c_17_24_b c_17_24_a c_17_24_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10233 vss n3713 c_18_22_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10232 n3546 c_17_23_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10231 vss c_17_23_a n3546 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10230 n3713 c_17_23_cin n3546 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10229 n3545 c_17_23_b n3713 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10228 vss c_17_23_a n3545 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10227 n3715 c_17_23_cin c_17_23_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10226 c_17_23_s2_s n3715 c_17_23_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10225 c_17_23_a c_17_23_b c_17_23_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10224 c_17_23_s1_s c_17_23_a c_17_23_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10223 c_18_21_a c_17_23_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10222 vss c_17_23_s1_s n3715 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10221 n3720 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10220 vss a_21 n3550 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10219 n3550 p_17_2_d2j n3719 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10218 n3719 p_17_2_d2jbar n3554 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10217 n3554 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10216 vss p_17_23_t_s c_17_23_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10215 c_17_23_b p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10214 n3719 n3720 p_17_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10213 p_17_23_t_s n3719 n3720 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10212 n4153 p_17_2_d2j n4157 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10211 n4154 p_17_2_d2jbar n4153 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10210 p_17_22_t_s n4153 n4151 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10209 n4153 n4151 p_17_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10208 p_17_22_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10207 vss p_17_22_t_s p_17_22_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10206 n4151 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10205 vss a_21 n4154 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10204 n4157 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10203 vss c_17_22_s1_s n4147 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10202 c_18_20_a c_17_22_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10201 c_17_22_s1_s p_17_22_pi2j c_17_22_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10200 c_17_22_s2_s n4147 c_16_23_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10199 n4147 c_16_23_cout c_17_22_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10198 vss p_17_22_pi2j n4144 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10197 n4144 c_17_22_a n4143 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10196 n4143 c_16_23_cout n4142 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10195 vss p_17_22_pi2j n4142 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10194 n4142 c_17_22_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10193 vss n4143 c_18_21_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10192 p_17_22_pi2j c_17_22_a c_17_22_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10191 vss n4472 c_18_20_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10190 n4361 p_17_21_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10189 vss c_17_21_a n4361 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10188 n4472 c_17_21_cin n4361 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10187 n4360 p_17_21_pi2j n4472 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10186 vss c_17_21_a n4360 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10185 n4469 c_17_21_cin c_17_21_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10184 c_17_21_s2_s n4469 c_17_21_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10183 c_17_21_a p_17_21_pi2j c_17_21_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10182 c_17_21_s1_s c_17_21_a p_17_21_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10181 c_18_19_a c_17_21_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10180 vss c_17_21_s1_s n4469 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10179 n4479 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10178 vss a_19 n4362 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10177 n4362 p_17_2_d2j n4478 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10176 n4478 p_17_2_d2jbar n4364 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10175 n4364 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10174 vss p_17_21_t_s p_17_21_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10173 p_17_21_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10172 n4478 n4479 p_17_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10171 p_17_21_t_s n4478 n4479 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10170 n4899 p_17_2_d2j n4902 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10169 n4900 p_17_2_d2jbar n4899 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10168 p_17_20_t_s n4899 n4897 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10167 n4899 n4897 p_17_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10166 p_17_20_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10165 vss p_17_20_t_s p_17_20_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10164 n4897 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10163 vss a_19 n4900 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10162 n4902 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10161 vss c_17_20_s1_s n4895 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10160 c_18_18_a c_17_20_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10159 c_17_20_s1_s p_17_20_pi2j c_17_20_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10158 c_17_20_s2_s n4895 c_16_21_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10157 n4895 c_16_21_cout c_17_20_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10156 vss p_17_20_pi2j n4888 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10155 n4888 c_17_20_a n4890 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10154 n4890 c_16_21_cout n4889 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10153 vss p_17_20_pi2j n4889 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10152 n4889 c_17_20_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10151 vss n4890 c_18_19_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10150 p_17_20_pi2j c_17_20_a c_17_20_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10149 vss n5214 c_18_18_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10148 n5102 p_17_19_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10147 vss c_17_19_a n5102 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10146 n5214 c_17_19_cin n5102 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10145 n5101 p_17_19_pi2j n5214 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10144 vss c_17_19_a n5101 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10143 n5209 c_17_19_cin c_17_19_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10142 c_17_19_s2_s n5209 c_17_19_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10141 c_17_19_a p_17_19_pi2j c_17_19_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10140 c_17_19_s1_s c_17_19_a p_17_19_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10139 c_18_17_a c_17_19_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10138 vss c_17_19_s1_s n5209 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10137 n5222 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10136 vss a_17 n5103 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10135 n5103 p_17_2_d2j n5220 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10134 n5220 p_17_2_d2jbar n5105 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10133 n5105 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10132 vss p_17_19_t_s p_17_19_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10131 p_17_19_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10130 n5220 n5222 p_17_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10129 p_17_19_t_s n5220 n5222 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10128 n5651 p_17_2_d2j n5657 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10127 n5650 p_17_2_d2jbar n5651 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10126 p_17_18_t_s n5651 n5653 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10125 n5651 n5653 p_17_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10124 p_17_18_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10123 vss p_17_18_t_s p_17_18_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10122 n5653 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10121 vss a_17 n5650 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10120 n5657 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10119 vss c_17_18_s1_s n5507 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10118 c_18_16_a c_17_18_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10117 c_17_18_s1_s p_17_18_pi2j c_17_18_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10116 c_17_18_s2_s n5507 c_16_19_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10115 n5507 c_16_19_cout c_17_18_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10114 vss p_17_18_pi2j n5644 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10113 n5644 c_17_18_a n5642 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10112 n5642 c_16_19_cout n5643 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10111 vss p_17_18_pi2j n5643 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10110 n5643 c_17_18_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10109 vss n5642 c_18_17_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10108 p_17_18_pi2j c_17_18_a c_17_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10107 vss n5989 c_18_16_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10106 n5862 p_17_17_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10105 vss c_17_17_a n5862 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10104 n5989 c_17_17_cin n5862 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10103 n5641 p_17_17_pi2j n5989 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10102 vss c_17_17_a n5641 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10101 n5979 c_17_17_cin c_17_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10100 c_17_17_s2_s n5979 c_17_17_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10099 c_17_17_a p_17_17_pi2j c_17_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10098 c_17_17_s1_s c_17_17_a p_17_17_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10097 c_18_15_a c_17_17_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10096 vss c_17_17_s1_s n5979 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10095 n5996 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10094 vss a_15 n5864 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10093 n5864 p_17_2_d2j n5990 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10092 n5990 p_17_2_d2jbar n5866 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10091 n5866 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10090 vss p_17_17_t_s p_17_17_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10089 p_17_17_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10088 n5990 n5996 p_17_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10087 p_17_17_t_s n5990 n5996 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10086 n6310 p_17_2_d2j n6312 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10085 n6311 p_17_2_d2jbar n6310 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10084 p_17_16_t_s n6310 n6442 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10083 n6310 n6442 p_17_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10082 p_17_16_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10081 vss p_17_16_t_s p_17_16_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10080 n6442 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10079 vss a_15 n6311 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10078 n6312 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10077 vss c_17_16_s1_s n6309 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10076 c_18_14_a c_17_16_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10075 c_17_16_s1_s p_17_16_pi2j c_17_16_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10074 c_17_16_s2_s n6309 c_16_17_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10073 n6309 c_16_17_cout c_17_16_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10072 vss p_17_16_pi2j n6435 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10071 n6435 c_17_16_a n6436 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10070 n6436 c_16_17_cout n6432 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10069 vss p_17_16_pi2j n6432 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10068 n6432 c_17_16_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10067 vss n6436 c_18_15_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10066 p_17_16_pi2j c_17_16_a c_17_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10065 vss n6826 c_18_14_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10064 n6434 c_17_15_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10063 vss c_17_15_a n6434 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10062 n6826 c_17_15_cin n6434 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10061 n6433 c_17_15_b n6826 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10060 vss c_17_15_a n6433 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10059 n6650 c_17_15_cin c_17_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10058 c_17_15_s2_s n6650 c_17_15_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10057 c_17_15_a c_17_15_b c_17_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10056 c_17_15_s1_s c_17_15_a c_17_15_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10055 c_18_13_a c_17_15_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10054 vss c_17_15_s1_s n6650 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10053 n6830 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10052 vss a_13 n6443 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10051 n6443 p_17_2_d2j n6653 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10050 n6653 p_17_2_d2jbar n6448 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10049 n6448 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10048 vss p_17_15_t_s c_17_15_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10047 c_17_15_b p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10046 n6653 n6830 p_17_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10045 p_17_15_t_s n6653 n6830 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10044 n7078 p_17_2_d2j n7080 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10043 n7079 p_17_2_d2jbar n7078 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10042 p_17_14_t_s n7078 n7077 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10041 n7078 n7077 p_17_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10040 p_17_14_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10039 vss p_17_14_t_s p_17_14_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10038 n7077 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10037 vss a_13 n7079 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10036 n7080 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10035 vss c_17_14_s1_s n7074 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10034 c_18_12_a c_17_14_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10033 c_17_14_s1_s p_17_14_pi2j c_17_14_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10032 c_17_14_s2_s n7074 c_16_15_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10031 n7074 c_16_15_cout c_17_14_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10030 vss p_17_14_pi2j n7244 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10029 n7244 c_17_14_a n7071 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10028 n7071 c_16_15_cout n7241 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10027 vss p_17_14_pi2j n7241 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10026 n7241 c_17_14_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10025 vss n7071 c_18_13_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10024 p_17_14_pi2j c_17_14_a c_17_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10023 vss n7411 c_18_12_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_10022 n7243 c_17_13_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10021 vss c_17_13_a n7243 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10020 n7411 c_17_13_cin n7243 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10019 n7242 c_17_13_b n7411 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10018 vss c_17_13_a n7242 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_10017 n7414 c_17_13_cin c_17_13_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10016 c_17_13_s2_s n7414 c_17_13_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10015 c_17_13_a c_17_13_b c_17_13_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10014 c_17_13_s1_s c_17_13_a c_17_13_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_10013 c_18_11_a c_17_13_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_10012 vss c_17_13_s1_s n7414 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_10011 n7418 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10010 vss a_11 n7248 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10009 n7248 p_17_2_d2j n7417 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10008 n7417 p_17_2_d2jbar n7251 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10007 n7251 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_10006 vss p_17_13_t_s c_17_13_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10005 c_17_13_b p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_10004 n7417 n7418 p_17_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10003 p_17_13_t_s n7417 n7418 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10002 n7845 p_17_2_d2j n7848 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_10001 n7846 p_17_2_d2jbar n7845 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_10000 p_17_12_t_s n7845 n7843 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09999 n7845 n7843 p_17_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09998 c_17_12_b p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09997 vss p_17_12_t_s c_17_12_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09996 n7843 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09995 vss a_11 n7846 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09994 n7848 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09993 vss c_17_12_s1_s n7840 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09992 c_18_10_a c_17_12_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09991 c_17_12_s1_s c_17_12_b c_17_12_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09990 c_17_12_s2_s n7840 c_16_13_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09989 n7840 c_16_13_cout c_17_12_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09988 vss c_17_12_b n7836 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09987 n7836 c_17_12_a n7837 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09986 n7837 c_16_13_cout n7835 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09985 vss c_17_12_b n7835 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09984 n7835 c_17_12_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09983 vss n7837 c_18_11_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09982 c_17_12_b c_17_12_a c_17_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09981 vss n8159 c_18_10_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09980 n8038 p_17_11_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09979 vss c_17_11_a n8038 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09978 n8159 c_17_11_cin n8038 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09977 n8037 p_17_11_pi2j n8159 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09976 vss c_17_11_a n8037 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09975 n8155 c_17_11_cin c_17_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09974 c_17_11_s2_s n8155 c_17_11_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09973 c_17_11_a p_17_11_pi2j c_17_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09972 c_17_11_s1_s c_17_11_a p_17_11_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09971 c_18_9_a c_17_11_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09970 vss c_17_11_s1_s n8155 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09969 n8167 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09968 vss a_9 n8040 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09967 n8040 p_17_2_d2j n8166 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09966 n8166 p_17_2_d2jbar n8042 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09965 n8042 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09964 vss p_17_11_t_s p_17_11_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09963 p_17_11_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09962 n8166 n8167 p_17_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09961 p_17_11_t_s n8166 n8167 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09960 n8588 p_17_2_d2j n8591 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09959 n8589 p_17_2_d2jbar n8588 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09958 p_17_10_t_s n8588 n8586 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09957 n8588 n8586 p_17_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09956 p_17_10_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09955 vss p_17_10_t_s p_17_10_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09954 n8586 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09953 vss a_9 n8589 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09952 n8591 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09951 vss c_17_10_s1_s n8584 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09950 c_18_8_a c_17_10_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09949 c_17_10_s1_s p_17_10_pi2j c_17_10_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09948 c_17_10_s2_s n8584 c_16_11_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09947 n8584 c_16_11_cout c_17_10_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09946 vss p_17_10_pi2j n8577 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09945 n8577 c_17_10_a n8579 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09944 n8579 c_16_11_cout n8578 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09943 vss p_17_10_pi2j n8578 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09942 n8578 c_17_10_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09941 vss n8579 c_18_9_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09940 p_17_10_pi2j c_17_10_a c_17_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09939 vss n8902 c_18_8_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09938 n8794 p_17_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09937 vss c_17_9_a n8794 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09936 n8902 c_17_9_cin n8794 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09935 n8793 p_17_9_pi2j n8902 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09934 vss c_17_9_a n8793 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09933 n8897 c_17_9_cin c_17_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09932 c_17_9_s2_s n8897 c_17_9_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09931 c_17_9_a p_17_9_pi2j c_17_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09930 c_17_9_s1_s c_17_9_a p_17_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09929 c_18_7_a c_17_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09928 vss c_17_9_s1_s n8897 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09927 n8910 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09926 vss a_7 n8795 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09925 n8795 p_17_2_d2j n8908 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09924 n8908 p_17_2_d2jbar n8797 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09923 n8797 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09922 vss p_17_9_t_s p_17_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09921 p_17_9_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09920 n8908 n8910 p_17_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09919 p_17_9_t_s n8908 n8910 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09918 n9320 p_17_2_d2j n9326 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09917 n9319 p_17_2_d2jbar n9320 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09916 p_17_8_t_s n9320 n9322 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09915 n9320 n9322 p_17_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09914 p_17_8_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09913 vss p_17_8_t_s p_17_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09912 n9322 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09911 vss a_7 n9319 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09910 n9326 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09909 vss c_17_8_s1_s n9309 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09908 c_18_6_a c_17_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09907 c_17_8_s1_s p_17_8_pi2j c_17_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09906 c_17_8_s2_s n9309 c_16_9_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09905 n9309 c_16_9_cout c_17_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09904 vss p_17_8_pi2j n9313 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09903 n9313 c_17_8_a n9311 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09902 n9311 c_16_9_cout n9312 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09901 vss p_17_8_pi2j n9312 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09900 n9312 c_17_8_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09899 vss n9311 c_18_7_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09898 p_17_8_pi2j c_17_8_a c_17_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09897 vss n9670 c_18_6_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09896 n9540 p_17_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09895 vss c_17_7_a n9540 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09894 n9670 c_17_7_cin n9540 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09893 n9310 p_17_7_pi2j n9670 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09892 vss c_17_7_a n9310 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09891 n9667 c_17_7_cin c_17_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09890 c_17_7_s2_s n9667 c_17_7_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09889 c_17_7_a p_17_7_pi2j c_17_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09888 c_17_7_s1_s c_17_7_a p_17_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09887 c_18_5_a c_17_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09886 vss c_17_7_s1_s n9667 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09885 n9680 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09884 vss a_5 n9542 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09883 n9542 p_17_2_d2j n9674 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09882 n9674 p_17_2_d2jbar n9544 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09881 n9544 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09880 vss p_17_7_t_s p_17_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09879 p_17_7_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09878 n9674 n9680 p_17_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09877 p_17_7_t_s n9674 n9680 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09876 n10105 p_17_2_d2j n9994 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09875 n9993 p_17_2_d2jbar n10105 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09874 p_17_6_t_s n10105 n10104 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09873 n10105 n10104 p_17_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09872 p_17_6_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09871 vss p_17_6_t_s p_17_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09870 n10104 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09869 vss a_5 n9993 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09868 n9994 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09867 vss c_17_6_s1_s n9992 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09866 c_18_4_a c_17_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09865 c_17_6_s1_s p_17_6_pi2j c_17_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09864 c_17_6_s2_s n9992 c_16_7_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09863 n9992 c_16_7_cout c_17_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09862 vss p_17_6_pi2j n10098 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09861 n10098 c_17_6_a n10097 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09860 n10097 c_16_7_cout n10094 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09859 vss p_17_6_pi2j n10094 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09858 n10094 c_17_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09857 vss n10097 c_18_5_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09856 p_17_6_pi2j c_17_6_a c_17_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09855 vss n10494 c_18_4_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09854 n10321 c_17_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09853 vss c_17_5_a n10321 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09852 n10494 c_17_5_cin n10321 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09851 n10096 c_17_5_b n10494 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09850 vss c_17_5_a n10096 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09849 n10325 c_17_5_cin c_17_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09848 c_17_5_s2_s n10325 c_17_5_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09847 c_17_5_a c_17_5_b c_17_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09846 c_17_5_s1_s c_17_5_a c_17_5_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09845 c_18_3_a c_17_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09844 vss c_17_5_s1_s n10325 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09843 n10498 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09842 vss a_3 n10106 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09841 n10106 p_17_2_d2j n10495 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09840 n10495 p_17_2_d2jbar n10111 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09839 n10111 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09838 vss p_17_5_t_s c_17_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09837 c_17_5_b p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09836 n10495 n10498 p_17_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09835 p_17_5_t_s n10495 n10498 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09834 n10752 p_17_2_d2j n10754 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09833 n10753 p_17_2_d2jbar n10752 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09832 p_17_4_t_s n10752 n10751 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09831 n10752 n10751 p_17_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09830 p_17_4_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09829 vss p_17_4_t_s p_17_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09828 n10751 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09827 vss a_3 n10753 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09826 n10754 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09825 vss c_17_4_s1_s n10750 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09824 c_18_2_a c_17_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09823 c_17_4_s1_s p_17_4_pi2j c_17_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09822 c_17_4_s2_s n10750 c_16_5_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09821 n10750 c_16_5_cout c_17_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09820 vss p_17_4_pi2j n10912 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09819 n10912 c_17_4_a n10745 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09818 n10745 c_16_5_cout n10909 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09817 vss p_17_4_pi2j n10909 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09816 n10909 c_17_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09815 vss n10745 c_18_3_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09814 p_17_4_pi2j c_17_4_a c_17_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09813 vss n11076 c_18_2_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09812 n10911 c_17_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09811 vss c_17_3_a n10911 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09810 n11076 c_17_3_cin n10911 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09809 n10910 c_17_3_b n11076 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09808 vss c_17_3_a n10910 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09807 n11079 c_17_3_cin c_17_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09806 c_17_3_s2_s n11079 c_17_3_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09805 c_17_3_a c_17_3_b c_17_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09804 c_17_3_s1_s c_17_3_a c_17_3_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09803 c_18_1_a c_17_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09802 vss c_17_3_s1_s n11079 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09801 n11083 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09800 vss a_1 n10916 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09799 n10916 p_17_2_d2j n11082 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09798 n11082 p_17_2_d2jbar n10919 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09797 n10919 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09796 vss p_17_3_t_s c_17_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09795 c_17_3_b p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09794 n11082 n11083 p_17_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09793 p_17_3_t_s n11082 n11083 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09792 n11508 p_17_2_d2j n11511 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09791 n11509 p_17_2_d2jbar n11508 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09790 p_17_2_t_s n11508 n11506 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09789 n11508 n11506 p_17_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09788 c_17_2_b p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09787 vss p_17_2_t_s c_17_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09786 n11506 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09785 vss a_1 n11509 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09784 n11511 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09783 vss c_17_2_s1_s n11503 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09782 c_17_2_sum c_17_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09781 c_17_2_s1_s c_17_2_b c_17_2_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09780 c_17_2_s2_s n11503 c_16_3_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09779 n11503 c_16_3_cout c_17_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09778 vss c_17_2_b n11498 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09777 n11498 c_17_2_a n11500 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09776 n11500 c_16_3_cout n11499 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09775 vss c_17_2_b n11499 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09774 n11499 c_17_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09773 vss n11500 c_18_1_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09772 c_17_2_b c_17_2_a c_17_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09771 vss n11816 c_17_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09770 n11700 p_17_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09769 vss c_17_1_a n11700 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09768 n11816 c_17_1_cin n11700 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09767 n11699 p_17_1_pi2j n11816 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09766 vss c_17_1_a n11699 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09765 n11813 c_17_1_cin c_17_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09764 c_17_1_s2_s n11813 c_17_1_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09763 c_17_1_a p_17_1_pi2j c_17_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09762 c_17_1_s1_s c_17_1_a p_17_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09761 c_17_1_sum c_17_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09760 vss c_17_1_s1_s n11813 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09759 n11824 p_17_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09758 n11825 p_17_2_d2jbar n11704 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09757 n11704 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09756 vss p_17_1_t_s p_17_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09755 p_17_1_pi2j p_17_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09754 n11825 n11824 p_17_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09753 p_17_1_t_s n11825 n11824 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09752 cl4_17_s1_s n12204 c_16_1_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09751 n12204 c_16_1_sum cl4_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09750 vss cl4_17_s1_s p_26 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09749 vss c_16_1_sum n12194 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09748 n12194 n12204 n12193 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09747 n12192 n12193 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_09746 n12189 c_16_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_09745 vss c_16_2_sum n12189 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_09744 n12190 c_16_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09743 n12191 c_16_1_cout n12190 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09742 n12186 c_16_1_sum n12191 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09741 n12189 n12204 n12186 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09740 n12187 n12191 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_09739 cl4_17_s2_s c_16_1_cout c_16_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09738 c_16_1_cout c_16_2_sum cl4_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09737 vss cl4_17_s2_s n12185 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09736 cl4_17_s3_s n12185 n12192 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09735 n12185 n12192 cl4_17_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09734 vss cl4_17_s3_s p_27 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09733 vss c_16_33_s1_s n81 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09732 c_17_31_a c_16_33_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09731 c_16_33_s1_s c_16_31_a p_16_33_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09730 c_16_31_a p_16_33_pi2j c_16_33_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09729 c_16_33_s2_s n81 c_16_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09728 n81 c_16_32_cin c_16_33_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09727 vss c_16_31_a n9 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_09726 n9 p_16_33_pi2j n80 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09725 n80 c_16_32_cin n10 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09724 vss c_16_31_a n10 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_09723 n10 p_16_33_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09722 vss n80 c_17_32_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09721 n88 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09720 n89 a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09719 vss p_16_33_t_s p_16_33_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09718 p_16_33_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09717 n89 n88 p_16_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09716 p_16_33_t_s n89 n88 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09715 n437 p_16_2_d2j n436 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09714 n438 p_16_2_d2jbar n437 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09713 p_16_32_t_s n437 n435 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09712 n437 n435 p_16_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09711 p_16_32_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09710 vss p_16_32_t_s p_16_32_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09709 n435 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09708 vss a_31 n438 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09707 n436 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09706 vss c_16_32_s1_s n431 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09705 c_17_30_a c_16_32_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09704 c_16_32_s1_s p_16_32_pi2j c_16_31_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09703 c_16_32_s2_s n431 c_16_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09702 n431 c_16_32_cin c_16_32_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09701 vss p_16_32_pi2j n426 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09700 n426 c_16_31_a n425 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09699 n425 c_16_32_cin n428 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09698 vss p_16_32_pi2j n428 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09697 n428 c_16_31_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09696 vss n425 c_17_31_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09695 p_16_32_pi2j c_16_31_a c_16_32_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09694 vss n745 c_16_31_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09693 n614 p_16_31_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09692 vss c_16_31_a n614 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09691 n745 c_16_31_cin n614 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09690 n612 p_16_31_pi2j n745 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09689 vss c_16_31_a n612 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09688 n740 c_16_31_cin c_16_31_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09687 c_16_31_s2_s n740 c_16_31_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09686 c_16_31_a p_16_31_pi2j c_16_31_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09685 c_16_31_s1_s c_16_31_a p_16_31_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09684 c_17_29_a c_16_31_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09683 vss c_16_31_s1_s n740 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09682 n749 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09681 vss a_29 n615 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09680 n615 p_16_2_d2j n751 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09679 n751 p_16_2_d2jbar n616 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09678 n616 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09677 vss p_16_31_t_s p_16_31_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09676 p_16_31_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09675 n751 n749 p_16_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09674 p_16_31_t_s n751 n749 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09673 n1181 p_16_2_d2j n1179 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09672 n1180 p_16_2_d2jbar n1181 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09671 p_16_30_t_s n1181 n1178 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09670 n1181 n1178 p_16_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09669 p_16_30_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09668 vss p_16_30_t_s p_16_30_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09667 n1178 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09666 vss a_29 n1180 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09665 n1179 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09664 vss c_16_30_s1_s n1173 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09663 c_17_28_a c_16_30_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09662 c_16_30_s1_s p_16_30_pi2j c_16_30_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09661 c_16_30_s2_s n1173 c_15_31_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09660 n1173 c_15_31_cout c_16_30_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09659 vss p_16_30_pi2j n1168 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09658 n1168 c_16_30_a n1167 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09657 n1167 c_15_31_cout n1170 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09656 vss p_16_30_pi2j n1170 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09655 n1170 c_16_30_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09654 vss n1167 c_17_29_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09653 p_16_30_pi2j c_16_30_a c_16_30_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09652 vss n1509 c_16_29_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09651 n1385 p_16_29_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09650 vss c_16_29_a n1385 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09649 n1509 c_16_29_cin n1385 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09648 n1166 p_16_29_pi2j n1509 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09647 vss c_16_29_a n1166 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09646 n1506 c_16_29_cin c_16_29_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09645 c_16_29_s2_s n1506 c_16_29_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09644 c_16_29_a p_16_29_pi2j c_16_29_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09643 c_16_29_s1_s c_16_29_a p_16_29_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09642 c_17_27_a c_16_29_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09641 vss c_16_29_s1_s n1506 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09640 n1513 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09639 vss a_27 n1386 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09638 n1386 p_16_2_d2j n1516 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09637 n1516 p_16_2_d2jbar n1387 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09636 n1387 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09635 vss p_16_29_t_s p_16_29_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09634 p_16_29_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09633 n1516 n1513 p_16_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09632 p_16_29_t_s n1516 n1513 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09631 n1942 p_16_2_d2j n1940 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09630 n1941 p_16_2_d2jbar n1942 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09629 p_16_28_t_s n1942 n1939 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09628 n1942 n1939 p_16_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09627 p_16_28_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09626 vss p_16_28_t_s p_16_28_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09625 n1939 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09624 vss a_27 n1941 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09623 n1940 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09622 vss c_16_28_s1_s n1789 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09621 c_17_26_a c_16_28_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09620 c_16_28_s1_s p_16_28_pi2j c_16_28_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09619 c_16_28_s2_s n1789 c_15_29_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09618 n1789 c_15_29_cout c_16_28_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09617 vss p_16_28_pi2j n1930 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09616 n1930 c_16_28_a n1929 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09615 n1929 c_15_29_cout n1933 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09614 vss p_16_28_pi2j n1933 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09613 n1933 c_16_28_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09612 vss n1929 c_17_27_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09611 p_16_28_pi2j c_16_28_a c_16_28_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09610 vss n2320 c_16_27_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09609 n2148 c_16_27_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09608 vss c_16_27_a n2148 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09607 n2320 c_16_27_cin n2148 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09606 n1928 c_16_27_b n2320 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09605 vss c_16_27_a n1928 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09604 n2312 c_16_27_cin c_16_27_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09603 c_16_27_s2_s n2312 c_16_27_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09602 c_16_27_a c_16_27_b c_16_27_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09601 c_16_27_s1_s c_16_27_a c_16_27_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09600 c_17_25_a c_16_27_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09599 vss c_16_27_s1_s n2312 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09598 n2323 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09597 vss a_25 n2154 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09596 n2154 p_16_2_d2j n2322 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09595 n2322 p_16_2_d2jbar n2153 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09594 n2153 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09593 vss p_16_27_t_s c_16_27_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09592 c_16_27_b p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09591 n2322 n2323 p_16_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09590 p_16_27_t_s n2322 n2323 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09589 n2610 p_16_2_d2j n2609 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09588 n2611 p_16_2_d2jbar n2610 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09587 p_16_26_t_s n2610 n2608 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09586 n2610 n2608 p_16_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09585 p_16_26_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09584 vss p_16_26_t_s p_16_26_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09583 n2608 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09582 vss a_25 n2611 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09581 n2609 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09580 vss c_16_26_s1_s n2607 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09579 c_17_24_a c_16_26_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09578 c_16_26_s1_s p_16_26_pi2j c_16_26_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09577 c_16_26_s2_s n2607 c_15_27_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09576 n2607 c_15_27_cout c_16_26_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09575 vss p_16_26_pi2j n2759 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09574 n2759 c_16_26_a n2758 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09573 n2758 c_15_27_cout n2760 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09572 vss p_16_26_pi2j n2760 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09571 n2760 c_16_26_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09570 vss n2758 c_17_25_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09569 p_16_26_pi2j c_16_26_a c_16_26_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09568 vss n3141 c_16_25_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09567 n2763 c_16_25_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09566 vss c_16_25_a n2763 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09565 n3141 c_16_25_cin n2763 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09564 n2757 c_16_25_b n3141 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09563 vss c_16_25_a n2757 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09562 n2959 c_16_25_cin c_16_25_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09561 c_16_25_s2_s n2959 c_16_25_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09560 c_16_25_a c_16_25_b c_16_25_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09559 c_16_25_s1_s c_16_25_a c_16_25_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09558 c_17_23_a c_16_25_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09557 vss c_16_25_s1_s n2959 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09556 n3143 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09555 vss a_23 n2768 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09554 n2768 p_16_2_d2j n2962 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09553 n2962 p_16_2_d2jbar n2769 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09552 n2769 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09551 vss p_16_25_t_s c_16_25_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09550 c_16_25_b p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09549 n2962 n3143 p_16_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09548 p_16_25_t_s n2962 n3143 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09547 n3384 p_16_2_d2j n3383 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09546 n3385 p_16_2_d2jbar n3384 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09545 p_16_24_t_s n3384 n3382 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09544 n3384 n3382 p_16_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09543 c_16_24_b p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09542 vss p_16_24_t_s c_16_24_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09541 n3382 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09540 vss a_23 n3385 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09539 n3383 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09538 vss c_16_24_s1_s n3379 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09537 c_17_22_a c_16_24_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09536 c_16_24_s1_s c_16_24_b c_16_24_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09535 c_16_24_s2_s n3379 c_15_25_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09534 n3379 c_15_25_cout c_16_24_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09533 vss c_16_24_b n3553 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09532 n3553 c_16_24_a n3375 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09531 n3375 c_15_25_cout n3552 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09530 vss c_16_24_b n3552 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09529 n3552 c_16_24_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09528 vss n3375 c_17_23_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09527 c_16_24_b c_16_24_a c_16_24_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09526 vss n3731 c_16_23_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09525 n3555 c_16_23_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09524 vss c_16_23_a n3555 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09523 n3731 c_16_23_cin n3555 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09522 n3551 c_16_23_b n3731 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09521 vss c_16_23_a n3551 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09520 n3732 c_16_23_cin c_16_23_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09519 c_16_23_s2_s n3732 c_16_23_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09518 c_16_23_a c_16_23_b c_16_23_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09517 c_16_23_s1_s c_16_23_a c_16_23_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09516 c_17_21_a c_16_23_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09515 vss c_16_23_s1_s n3732 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09514 n3735 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09513 vss a_21 n3558 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09512 n3558 p_16_2_d2j n3737 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09511 n3737 p_16_2_d2jbar n3559 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09510 n3559 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09509 vss p_16_23_t_s c_16_23_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09508 c_16_23_b p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09507 n3737 n3735 p_16_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09506 p_16_23_t_s n3737 n3735 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09505 n4168 p_16_2_d2j n4167 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09504 n4169 p_16_2_d2jbar n4168 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09503 p_16_22_t_s n4168 n4166 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09502 n4168 n4166 p_16_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09501 p_16_22_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09500 vss p_16_22_t_s p_16_22_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09499 n4166 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09498 vss a_21 n4169 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09497 n4167 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09496 vss c_16_22_s1_s n4161 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09495 c_17_20_a c_16_22_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09494 c_16_22_s1_s p_16_22_pi2j c_16_22_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09493 c_16_22_s2_s n4161 c_15_23_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09492 n4161 c_15_23_cout c_16_22_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09491 vss p_16_22_pi2j n4156 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09490 n4156 c_16_22_a n4155 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09489 n4155 c_15_23_cout n4158 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09488 vss p_16_22_pi2j n4158 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09487 n4158 c_16_22_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09486 vss n4155 c_17_21_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09485 p_16_22_pi2j c_16_22_a c_16_22_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09484 vss n4492 c_16_21_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09483 n4365 p_16_21_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09482 vss c_16_21_a n4365 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09481 n4492 c_16_21_cin n4365 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09480 n4363 p_16_21_pi2j n4492 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09479 vss c_16_21_a n4363 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09478 n4489 c_16_21_cin c_16_21_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09477 c_16_21_s2_s n4489 c_16_21_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09476 c_16_21_a p_16_21_pi2j c_16_21_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09475 c_16_21_s1_s c_16_21_a p_16_21_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09474 c_17_19_a c_16_21_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09473 vss c_16_21_s1_s n4489 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09472 n4496 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09471 vss a_19 n4366 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09470 n4366 p_16_2_d2j n4498 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09469 n4498 p_16_2_d2jbar n4367 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09468 n4367 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09467 vss p_16_21_t_s p_16_21_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09466 p_16_21_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09465 n4498 n4496 p_16_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09464 p_16_21_t_s n4498 n4496 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09463 n4914 p_16_2_d2j n4913 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09462 n4915 p_16_2_d2jbar n4914 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09461 p_16_20_t_s n4914 n4912 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09460 n4914 n4912 p_16_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09459 p_16_20_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09458 vss p_16_20_t_s p_16_20_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09457 n4912 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09456 vss a_19 n4915 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09455 n4913 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09454 vss c_16_20_s1_s n4909 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09453 c_17_18_a c_16_20_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09452 c_16_20_s1_s p_16_20_pi2j c_16_20_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09451 c_16_20_s2_s n4909 c_15_21_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09450 n4909 c_15_21_cout c_16_20_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09449 vss p_16_20_pi2j n4903 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09448 n4903 c_16_20_a n4901 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09447 n4901 c_15_21_cout n4904 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09446 vss p_16_20_pi2j n4904 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09445 n4904 c_16_20_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09444 vss n4901 c_17_19_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09443 p_16_20_pi2j c_16_20_a c_16_20_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09442 vss n5236 c_16_19_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09441 n5106 p_16_19_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09440 vss c_16_19_a n5106 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09439 n5236 c_16_19_cin n5106 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09438 n5104 p_16_19_pi2j n5236 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09437 vss c_16_19_a n5104 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09436 n5232 c_16_19_cin c_16_19_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09435 c_16_19_s2_s n5232 c_16_19_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09434 c_16_19_a p_16_19_pi2j c_16_19_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09433 c_16_19_s1_s c_16_19_a p_16_19_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09432 c_17_17_a c_16_19_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09431 vss c_16_19_s1_s n5232 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09430 n5240 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09429 vss a_17 n5107 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09428 n5107 p_16_2_d2j n5243 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09427 n5243 p_16_2_d2jbar n5108 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09426 n5108 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09425 vss p_16_19_t_s p_16_19_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09424 p_16_19_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09423 n5243 n5240 p_16_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09422 p_16_19_t_s n5243 n5240 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09421 n5666 p_16_2_d2j n5668 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09420 n5665 p_16_2_d2jbar n5666 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09419 p_16_18_t_s n5666 n5667 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09418 n5666 n5667 p_16_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09417 p_16_18_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09416 vss p_16_18_t_s p_16_18_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09415 n5667 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09414 vss a_17 n5665 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09413 n5668 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09412 vss c_16_18_s1_s n5515 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09411 c_17_16_a c_16_18_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09410 c_16_18_s1_s p_16_18_pi2j c_16_18_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09409 c_16_18_s2_s n5515 c_15_19_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09408 n5515 c_15_19_cout c_16_18_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09407 vss p_16_18_pi2j n5655 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09406 n5655 c_16_18_a n5656 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09405 n5656 c_15_19_cout n5659 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09404 vss p_16_18_pi2j n5659 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09403 n5659 c_16_18_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09402 vss n5656 c_17_17_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09401 p_16_18_pi2j c_16_18_a c_16_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09400 vss n6013 c_16_17_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09399 n5867 p_16_17_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09398 vss c_16_17_a n5867 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09397 n6013 c_16_17_cin n5867 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09396 n5654 p_16_17_pi2j n6013 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09395 vss c_16_17_a n5654 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09394 n6003 c_16_17_cin c_16_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09393 c_16_17_s2_s n6003 c_16_17_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09392 c_16_17_a p_16_17_pi2j c_16_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09391 c_16_17_s1_s c_16_17_a p_16_17_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09390 c_17_15_a c_16_17_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09389 vss c_16_17_s1_s n6003 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09388 n6015 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09387 vss a_15 n5870 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09386 n5870 p_16_2_d2j n6014 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09385 n6014 p_16_2_d2jbar n5871 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09384 n5871 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09383 vss p_16_17_t_s p_16_17_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09382 p_16_17_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09381 n6014 n6015 p_16_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09380 p_16_17_t_s n6014 n6015 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09379 n6318 p_16_2_d2j n6317 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09378 n6319 p_16_2_d2jbar n6318 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09377 p_16_16_t_s n6318 n6454 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09376 n6318 n6454 p_16_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09375 p_16_16_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09374 vss p_16_16_t_s p_16_16_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09373 n6454 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09372 vss a_15 n6319 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09371 n6317 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09370 vss c_16_16_s1_s n6316 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09369 c_17_14_a c_16_16_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09368 c_16_16_s1_s p_16_16_pi2j c_16_16_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09367 c_16_16_s2_s n6316 c_15_17_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09366 n6316 c_15_17_cout c_16_16_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09365 vss p_16_16_pi2j n6446 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09364 n6446 c_16_16_a n6447 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09363 n6447 c_15_17_cout n6445 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09362 vss p_16_16_pi2j n6445 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09361 n6445 c_16_16_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09360 vss n6447 c_17_15_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09359 p_16_16_pi2j c_16_16_a c_16_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09358 vss n6842 c_16_15_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09357 n6450 c_16_15_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09356 vss c_16_15_a n6450 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09355 n6842 c_16_15_cin n6450 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09354 n6444 c_16_15_b n6842 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09353 vss c_16_15_a n6444 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09352 n6660 c_16_15_cin c_16_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09351 c_16_15_s2_s n6660 c_16_15_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09350 c_16_15_a c_16_15_b c_16_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09349 c_16_15_s1_s c_16_15_a c_16_15_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09348 c_17_13_a c_16_15_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09347 vss c_16_15_s1_s n6660 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09346 n6845 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09345 vss a_13 n6456 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09344 n6456 p_16_2_d2j n6663 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09343 n6663 p_16_2_d2jbar n6457 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09342 n6457 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09341 vss p_16_15_t_s c_16_15_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09340 c_16_15_b p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09339 n6663 n6845 p_16_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09338 p_16_15_t_s n6663 n6845 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09337 n7089 p_16_2_d2j n7088 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09336 n7090 p_16_2_d2jbar n7089 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09335 p_16_14_t_s n7089 n7087 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09334 n7089 n7087 p_16_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09333 p_16_14_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09332 vss p_16_14_t_s p_16_14_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09331 n7087 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09330 vss a_13 n7090 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09329 n7088 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09328 vss c_16_14_s1_s n7084 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09327 c_17_12_a c_16_14_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09326 c_16_14_s1_s p_16_14_pi2j c_16_14_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09325 c_16_14_s2_s n7084 c_15_15_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09324 n7084 c_15_15_cout c_16_14_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09323 vss p_16_14_pi2j n7252 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09322 n7252 c_16_14_a n7081 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09321 n7081 c_15_15_cout n7250 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09320 vss p_16_14_pi2j n7250 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09319 n7250 c_16_14_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09318 vss n7081 c_17_13_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09317 p_16_14_pi2j c_16_14_a c_16_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09316 vss n7425 c_16_13_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09315 n7254 c_16_13_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09314 vss c_16_13_a n7254 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09313 n7425 c_16_13_cin n7254 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09312 n7249 c_16_13_b n7425 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09311 vss c_16_13_a n7249 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09310 n7428 c_16_13_cin c_16_13_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09309 c_16_13_s2_s n7428 c_16_13_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09308 c_16_13_a c_16_13_b c_16_13_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09307 c_16_13_s1_s c_16_13_a c_16_13_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09306 c_17_11_a c_16_13_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09305 vss c_16_13_s1_s n7428 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09304 n7430 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09303 vss a_11 n7257 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09302 n7257 p_16_2_d2j n7432 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09301 n7432 p_16_2_d2jbar n7258 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09300 n7258 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09299 vss p_16_13_t_s c_16_13_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09298 c_16_13_b p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09297 n7432 n7430 p_16_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09296 p_16_13_t_s n7432 n7430 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09295 n7859 p_16_2_d2j n7858 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09294 n7860 p_16_2_d2jbar n7859 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09293 p_16_12_t_s n7859 n7857 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09292 n7859 n7857 p_16_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09291 c_16_12_b p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09290 vss p_16_12_t_s c_16_12_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09289 n7857 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09288 vss a_11 n7860 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09287 n7858 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09286 vss c_16_12_s1_s n7853 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09285 c_17_10_a c_16_12_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09284 c_16_12_s1_s c_16_12_b c_16_12_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09283 c_16_12_s2_s n7853 c_15_13_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09282 n7853 c_15_13_cout c_16_12_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09281 vss c_16_12_b n7849 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09280 n7849 c_16_12_a n7847 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09279 n7847 c_15_13_cout n7850 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09278 vss c_16_12_b n7850 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09277 n7850 c_16_12_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09276 vss n7847 c_17_11_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09275 c_16_12_b c_16_12_a c_16_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09274 vss n8178 c_16_11_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09273 n8043 p_16_11_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09272 vss c_16_11_a n8043 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09271 n8178 c_16_11_cin n8043 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09270 n8041 p_16_11_pi2j n8178 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09269 vss c_16_11_a n8041 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09268 n8177 c_16_11_cin c_16_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09267 c_16_11_s2_s n8177 c_16_11_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09266 c_16_11_a p_16_11_pi2j c_16_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09265 c_16_11_s1_s c_16_11_a p_16_11_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09264 c_17_9_a c_16_11_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09263 vss c_16_11_s1_s n8177 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09262 n8184 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09261 vss a_9 n8045 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09260 n8045 p_16_2_d2j n8186 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09259 n8186 p_16_2_d2jbar n8046 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09258 n8046 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09257 vss p_16_11_t_s p_16_11_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09256 p_16_11_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09255 n8186 n8184 p_16_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09254 p_16_11_t_s n8186 n8184 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09253 n8603 p_16_2_d2j n8602 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09252 n8604 p_16_2_d2jbar n8603 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09251 p_16_10_t_s n8603 n8601 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09250 n8603 n8601 p_16_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09249 p_16_10_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09248 vss p_16_10_t_s p_16_10_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09247 n8601 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09246 vss a_9 n8604 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09245 n8602 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09244 vss c_16_10_s1_s n8596 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09243 c_17_8_a c_16_10_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09242 c_16_10_s1_s p_16_10_pi2j c_16_10_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09241 c_16_10_s2_s n8596 c_15_11_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09240 n8596 c_15_11_cout c_16_10_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09239 vss p_16_10_pi2j n8592 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09238 n8592 c_16_10_a n8590 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09237 n8590 c_15_11_cout n8593 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09236 vss p_16_10_pi2j n8593 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09235 n8593 c_16_10_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09234 vss n8590 c_17_9_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09233 p_16_10_pi2j c_16_10_a c_16_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09232 vss n8924 c_16_9_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09231 n8798 p_16_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09230 vss c_16_9_a n8798 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09229 n8924 c_16_9_cin n8798 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09228 n8796 p_16_9_pi2j n8924 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09227 vss c_16_9_a n8796 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09226 n8920 c_16_9_cin c_16_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09225 c_16_9_s2_s n8920 c_16_9_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09224 c_16_9_a p_16_9_pi2j c_16_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09223 c_16_9_s1_s c_16_9_a p_16_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09222 c_17_7_a c_16_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09221 vss c_16_9_s1_s n8920 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09220 n8928 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09219 vss a_7 n8799 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09218 n8799 p_16_2_d2j n8931 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09217 n8931 p_16_2_d2jbar n8800 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09216 n8800 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09215 vss p_16_9_t_s p_16_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09214 p_16_9_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09213 n8931 n8928 p_16_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09212 p_16_9_t_s n8931 n8928 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09211 n9336 p_16_2_d2j n9338 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09210 n9335 p_16_2_d2jbar n9336 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09209 p_16_8_t_s n9336 n9337 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09208 n9336 n9337 p_16_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09207 p_16_8_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09206 vss p_16_8_t_s p_16_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09205 n9337 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09204 vss a_7 n9335 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09203 n9338 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09202 vss c_16_8_s1_s n9327 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09201 c_17_6_a c_16_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09200 c_16_8_s1_s p_16_8_pi2j c_16_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09199 c_16_8_s2_s n9327 c_15_9_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09198 n9327 c_15_9_cout c_16_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09197 vss p_16_8_pi2j n9324 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09196 n9324 c_16_8_a n9325 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09195 n9325 c_15_9_cout n9329 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09194 vss p_16_8_pi2j n9329 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09193 n9329 c_16_8_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09192 vss n9325 c_17_7_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09191 p_16_8_pi2j c_16_8_a c_16_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09190 vss n9697 c_16_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09189 n9545 p_16_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09188 vss c_16_7_a n9545 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09187 n9697 c_16_7_cin n9545 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09186 n9323 p_16_7_pi2j n9697 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09185 vss c_16_7_a n9323 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09184 n9693 c_16_7_cin c_16_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09183 c_16_7_s2_s n9693 c_16_7_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09182 c_16_7_a p_16_7_pi2j c_16_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09181 c_16_7_s1_s c_16_7_a p_16_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09180 c_17_5_a c_16_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09179 vss c_16_7_s1_s n9693 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09178 n9699 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09177 vss a_5 n9548 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09176 n9548 p_16_2_d2j n9698 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09175 n9698 p_16_2_d2jbar n9549 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09174 n9549 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09173 vss p_16_7_t_s p_16_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09172 p_16_7_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09171 n9698 n9699 p_16_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09170 p_16_7_t_s n9698 n9699 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09169 n10118 p_16_2_d2j n9998 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09168 n9999 p_16_2_d2jbar n10118 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09167 p_16_6_t_s n10118 n10117 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09166 n10118 n10117 p_16_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09165 p_16_6_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09164 vss p_16_6_t_s p_16_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09163 n10117 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09162 vss a_5 n9999 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09161 n9998 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09160 vss c_16_6_s1_s n9997 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09159 c_17_4_a c_16_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09158 c_16_6_s1_s p_16_6_pi2j c_16_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09157 c_16_6_s2_s n9997 c_15_7_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09156 n9997 c_15_7_cout c_16_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09155 vss p_16_6_pi2j n10109 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09154 n10109 c_16_6_a n10110 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09153 n10110 c_15_7_cout n10108 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09152 vss p_16_6_pi2j n10108 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09151 n10108 c_16_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09150 vss n10110 c_17_5_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09149 p_16_6_pi2j c_16_6_a c_16_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09148 vss n10511 c_16_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09147 n10330 c_16_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09146 vss c_16_5_a n10330 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09145 n10511 c_16_5_cin n10330 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09144 n10107 c_16_5_b n10511 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09143 vss c_16_5_a n10107 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09142 n10335 c_16_5_cin c_16_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09141 c_16_5_s2_s n10335 c_16_5_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09140 c_16_5_a c_16_5_b c_16_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09139 c_16_5_s1_s c_16_5_a c_16_5_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09138 c_17_3_a c_16_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09137 vss c_16_5_s1_s n10335 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09136 n10515 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09135 vss a_3 n10120 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09134 n10120 p_16_2_d2j n10513 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09133 n10513 p_16_2_d2jbar n10121 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09132 n10121 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09131 vss p_16_5_t_s c_16_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09130 c_16_5_b p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09129 n10513 n10515 p_16_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09128 p_16_5_t_s n10513 n10515 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09127 n10763 p_16_2_d2j n10762 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09126 n10764 p_16_2_d2jbar n10763 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09125 p_16_4_t_s n10763 n10761 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09124 n10763 n10761 p_16_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09123 p_16_4_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09122 vss p_16_4_t_s p_16_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09121 n10761 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09120 vss a_3 n10764 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09119 n10762 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09118 vss c_16_4_s1_s n10759 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09117 c_17_2_a c_16_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09116 c_16_4_s1_s p_16_4_pi2j c_16_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09115 c_16_4_s2_s n10759 c_15_5_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09114 n10759 c_15_5_cout c_16_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09113 vss p_16_4_pi2j n10920 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09112 n10920 c_16_4_a n10755 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09111 n10755 c_15_5_cout n10918 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09110 vss p_16_4_pi2j n10918 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09109 n10918 c_16_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09108 vss n10755 c_17_3_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09107 p_16_4_pi2j c_16_4_a c_16_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09106 vss n11090 c_16_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09105 n10922 c_16_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09104 vss c_16_3_a n10922 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09103 n11090 c_16_3_cin n10922 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09102 n10917 c_16_3_b n11090 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09101 vss c_16_3_a n10917 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09100 n11093 c_16_3_cin c_16_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09099 c_16_3_s2_s n11093 c_16_3_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09098 c_16_3_a c_16_3_b c_16_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09097 c_16_3_s1_s c_16_3_a c_16_3_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09096 c_17_1_a c_16_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09095 vss c_16_3_s1_s n11093 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09094 n11095 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09093 vss a_1 n10925 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09092 n10925 p_16_2_d2j n11097 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09091 n11097 p_16_2_d2jbar n10926 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09090 n10926 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09089 vss p_16_3_t_s c_16_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09088 c_16_3_b p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09087 n11097 n11095 p_16_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09086 p_16_3_t_s n11097 n11095 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09085 n11522 p_16_2_d2j n11521 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09084 n11523 p_16_2_d2jbar n11522 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09083 p_16_2_t_s n11522 n11520 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09082 n11522 n11520 p_16_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09081 c_16_2_b p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09080 vss p_16_2_t_s c_16_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09079 n11520 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09078 vss a_1 n11523 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09077 n11521 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09076 vss c_16_2_s1_s n11516 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09075 c_16_2_sum c_16_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09074 c_16_2_s1_s c_16_2_b c_16_2_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09073 c_16_2_s2_s n11516 c_15_3_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09072 n11516 c_15_3_cout c_16_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09071 vss c_16_2_b n11512 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09070 n11512 c_16_2_a n11510 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09069 n11510 c_15_3_cout n11513 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09068 vss c_16_2_b n11513 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09067 n11513 c_16_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09066 vss n11510 c_17_1_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09065 c_16_2_b c_16_2_a c_16_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09064 vss n11837 c_16_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09063 n11705 p_16_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09062 vss c_16_1_a n11705 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09061 n11837 c_16_1_cin n11705 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09060 n11703 p_16_1_pi2j n11837 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09059 vss c_16_1_a n11703 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09058 n11833 c_16_1_cin c_16_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09057 c_16_1_s2_s n11833 c_16_1_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09056 c_16_1_a p_16_1_pi2j c_16_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09055 c_16_1_s1_s c_16_1_a p_16_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09054 c_16_1_sum c_16_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09053 vss c_16_1_s1_s n11833 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09052 n11844 p_16_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09051 n11845 p_16_2_d2jbar n11708 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09050 n11708 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09049 vss p_16_1_t_s p_16_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09048 p_16_1_pi2j p_16_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09047 n11845 n11844 p_16_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09046 p_16_1_t_s n11845 n11844 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_09045 cl4_16_s1_s n12221 c_15_1_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09044 n12221 c_15_1_sum cl4_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09043 vss cl4_16_s1_s p_24 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09042 vss c_15_1_sum n12211 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09041 n12211 n12221 n12210 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09040 n12209 n12210 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_09039 n12208 c_15_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_09038 vss c_15_2_sum n12208 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_09037 n12207 c_15_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09036 n12205 c_15_1_cout n12207 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09035 n12203 c_15_1_sum n12205 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09034 n12208 n12221 n12203 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09033 n12204 n12205 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_09032 cl4_16_s2_s c_15_1_cout c_15_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09031 c_15_1_cout c_15_2_sum cl4_16_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09030 vss cl4_16_s2_s n12200 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09029 cl4_16_s3_s n12200 n12209 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09028 n12200 n12209 cl4_16_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09027 vss cl4_16_s3_s p_25 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_09026 vss c_15_33_s1_s n98 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_09025 c_16_31_a c_15_33_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_09024 c_15_33_s1_s c_15_31_a p_15_33_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09023 c_15_31_a p_15_33_pi2j c_15_33_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09022 c_15_33_s2_s n98 c_15_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09021 n98 c_15_32_cin c_15_33_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_09020 vss c_15_31_a n11 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_09019 n11 p_15_33_pi2j n91 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09018 n91 c_15_32_cin n12 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09017 vss c_15_31_a n12 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_09016 n12 p_15_33_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_09015 vss n91 c_16_32_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_09014 n100 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09013 n103 a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09012 vss p_15_33_t_s p_15_33_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09011 p_15_33_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09010 n103 n100 p_15_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09009 p_15_33_t_s n103 n100 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09008 n450 p_15_2_d2j n451 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09007 n449 p_15_2_d2jbar n450 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09006 p_15_32_t_s n450 n447 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09005 n450 n447 p_15_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09004 p_15_32_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09003 vss p_15_32_t_s p_15_32_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_09002 n447 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_09001 vss a_31 n449 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_09000 n451 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08999 vss c_15_32_s1_s n444 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08998 c_16_30_a c_15_32_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08997 c_15_32_s1_s p_15_32_pi2j c_15_31_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08996 c_15_32_s2_s n444 c_15_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08995 n444 c_15_32_cin c_15_32_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08994 vss p_15_32_pi2j n440 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08993 n440 c_15_31_a n439 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08992 n439 c_15_32_cin n441 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08991 vss p_15_32_pi2j n441 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08990 n441 c_15_31_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08989 vss n439 c_16_31_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08988 p_15_32_pi2j c_15_31_a c_15_32_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08987 vss n756 c_15_31_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08986 n618 p_15_31_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08985 vss c_15_31_a n618 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08984 n756 c_15_31_cin n618 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08983 n617 p_15_31_pi2j n756 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08982 vss c_15_31_a n617 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08981 n764 c_15_31_cin c_15_31_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08980 c_15_31_s2_s n764 c_15_31_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08979 c_15_31_a p_15_31_pi2j c_15_31_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08978 c_15_31_s1_s c_15_31_a p_15_31_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08977 c_16_29_a c_15_31_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08976 vss c_15_31_s1_s n764 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08975 n767 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08974 vss a_29 n620 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08973 n620 p_15_2_d2j n769 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08972 n769 p_15_2_d2jbar n619 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08971 n619 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08970 vss p_15_31_t_s p_15_31_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08969 p_15_31_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08968 n769 n767 p_15_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08967 p_15_31_t_s n769 n767 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08966 n1196 p_15_2_d2j n1194 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08965 n1195 p_15_2_d2jbar n1196 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08964 p_15_30_t_s n1196 n1192 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08963 n1196 n1192 p_15_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08962 p_15_30_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08961 vss p_15_30_t_s p_15_30_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08960 n1192 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08959 vss a_29 n1195 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08958 n1194 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08957 vss c_15_30_s1_s n1188 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08956 c_16_28_a c_15_30_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08955 c_15_30_s1_s p_15_30_pi2j c_15_30_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08954 c_15_30_s2_s n1188 c_14_31_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08953 n1188 c_14_31_cout c_15_30_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08952 vss p_15_30_pi2j n1185 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08951 n1185 c_15_30_a n1183 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08950 n1183 c_14_31_cout n1184 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08949 vss p_15_30_pi2j n1184 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08948 n1184 c_15_30_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08947 vss n1183 c_16_29_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08946 p_15_30_pi2j c_15_30_a c_15_30_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08945 vss n1523 c_15_29_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08944 n1388 p_15_29_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08943 vss c_15_29_a n1388 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08942 n1523 c_15_29_cin n1388 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08941 n1182 p_15_29_pi2j n1523 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08940 vss c_15_29_a n1182 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08939 n1527 c_15_29_cin c_15_29_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08938 c_15_29_s2_s n1527 c_15_29_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08937 c_15_29_a p_15_29_pi2j c_15_29_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08936 c_15_29_s1_s c_15_29_a p_15_29_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08935 c_16_27_a c_15_29_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08934 vss c_15_29_s1_s n1527 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08933 n1533 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08932 vss a_27 n1390 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08931 n1390 p_15_2_d2j n1534 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08930 n1534 p_15_2_d2jbar n1389 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08929 n1389 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08928 vss p_15_29_t_s p_15_29_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08927 p_15_29_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08926 n1534 n1533 p_15_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08925 p_15_29_t_s n1534 n1533 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08924 n1956 p_15_2_d2j n1954 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08923 n1955 p_15_2_d2jbar n1956 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08922 p_15_28_t_s n1956 n1952 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08921 n1956 n1952 p_15_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08920 p_15_28_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08919 vss p_15_28_t_s p_15_28_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08918 n1952 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08917 vss a_27 n1955 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08916 n1954 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08915 vss c_15_28_s1_s n1795 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08914 c_16_26_a c_15_28_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08913 c_15_28_s1_s p_15_28_pi2j c_15_28_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08912 c_15_28_s2_s n1795 c_14_29_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08911 n1795 c_14_29_cout c_15_28_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08910 vss p_15_28_pi2j n1946 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08909 n1946 c_15_28_a n1945 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08908 n1945 c_14_29_cout n1944 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08907 vss p_15_28_pi2j n1944 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08906 n1944 c_15_28_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08905 vss n1945 c_16_27_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08904 p_15_28_pi2j c_15_28_a c_15_28_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08903 vss n2335 c_15_27_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08902 n2155 c_15_27_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08901 vss c_15_27_a n2155 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08900 n2335 c_15_27_cin n2155 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08899 n1943 c_15_27_b n2335 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08898 vss c_15_27_a n1943 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08897 n2331 c_15_27_cin c_15_27_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08896 c_15_27_s2_s n2331 c_15_27_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08895 c_15_27_a c_15_27_b c_15_27_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08894 c_15_27_s1_s c_15_27_a c_15_27_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08893 c_16_25_a c_15_27_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08892 vss c_15_27_s1_s n2331 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08891 n2343 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08890 vss a_25 n2160 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08889 n2160 p_15_2_d2j n2342 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08888 n2342 p_15_2_d2jbar n2161 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08887 n2161 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08886 vss p_15_27_t_s c_15_27_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08885 c_15_27_b p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08884 n2342 n2343 p_15_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08883 p_15_27_t_s n2342 n2343 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08882 n2618 p_15_2_d2j n2619 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08881 n2617 p_15_2_d2jbar n2618 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08880 p_15_26_t_s n2618 n2616 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08879 n2618 n2616 p_15_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08878 p_15_26_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08877 vss p_15_26_t_s p_15_26_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08876 n2616 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08875 vss a_25 n2617 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08874 n2619 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08873 vss c_15_26_s1_s n2615 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08872 c_16_24_a c_15_26_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08871 c_15_26_s1_s p_15_26_pi2j c_15_26_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08870 c_15_26_s2_s n2615 c_14_27_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08869 n2615 c_14_27_cout c_15_26_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08868 vss p_15_26_pi2j n2773 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08867 n2773 c_15_26_a n2772 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08866 n2772 c_14_27_cout n2774 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08865 vss p_15_26_pi2j n2774 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08864 n2774 c_15_26_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08863 vss n2772 c_16_25_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08862 p_15_26_pi2j c_15_26_a c_15_26_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08861 vss n3151 c_15_25_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08860 n2771 c_15_25_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08859 vss c_15_25_a n2771 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08858 n3151 c_15_25_cin n2771 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08857 n2770 c_15_25_b n3151 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08856 vss c_15_25_a n2770 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08855 n2968 c_15_25_cin c_15_25_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08854 c_15_25_s2_s n2968 c_15_25_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08853 c_15_25_a c_15_25_b c_15_25_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08852 c_15_25_s1_s c_15_25_a c_15_25_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08851 c_16_23_a c_15_25_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08850 vss c_15_25_s1_s n2968 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08849 n3159 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08848 vss a_23 n2780 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08847 n2780 p_15_2_d2j n2971 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08846 n2971 p_15_2_d2jbar n2781 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08845 n2781 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08844 vss p_15_25_t_s c_15_25_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08843 c_15_25_b p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08842 n2971 n3159 p_15_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08841 p_15_25_t_s n2971 n3159 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08840 n3395 p_15_2_d2j n3396 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08839 n3394 p_15_2_d2jbar n3395 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08838 p_15_24_t_s n3395 n3393 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08837 n3395 n3393 p_15_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08836 c_15_24_b p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08835 vss p_15_24_t_s c_15_24_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08834 n3393 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08833 vss a_23 n3394 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08832 n3396 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08831 vss c_15_24_s1_s n3390 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08830 c_16_22_a c_15_24_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08829 c_15_24_s1_s c_15_24_b c_15_24_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08828 c_15_24_s2_s n3390 c_14_25_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08827 n3390 c_14_25_cout c_15_24_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08826 vss c_15_24_b n3562 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08825 n3562 c_15_24_a n3386 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08824 n3386 c_14_25_cout n3563 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08823 vss c_15_24_b n3563 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08822 n3563 c_15_24_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08821 vss n3386 c_16_23_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08820 c_15_24_b c_15_24_a c_15_24_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08819 vss n3741 c_15_23_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08818 n3561 c_15_23_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08817 vss c_15_23_a n3561 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08816 n3741 c_15_23_cin n3561 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08815 n3560 c_15_23_b n3741 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08814 vss c_15_23_a n3560 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08813 n3747 c_15_23_cin c_15_23_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08812 c_15_23_s2_s n3747 c_15_23_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08811 c_15_23_a c_15_23_b c_15_23_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08810 c_15_23_s1_s c_15_23_a c_15_23_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08809 c_16_21_a c_15_23_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08808 vss c_15_23_s1_s n3747 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08807 n3751 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08806 vss a_21 n3567 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08805 n3567 p_15_2_d2j n3753 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08804 n3753 p_15_2_d2jbar n3566 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08803 n3566 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08802 vss p_15_23_t_s c_15_23_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08801 c_15_23_b p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08800 n3753 n3751 p_15_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08799 p_15_23_t_s n3753 n3751 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08798 n4182 p_15_2_d2j n4183 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08797 n4181 p_15_2_d2jbar n4182 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08796 p_15_22_t_s n4182 n4179 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08795 n4182 n4179 p_15_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08794 p_15_22_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08793 vss p_15_22_t_s p_15_22_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08792 n4179 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08791 vss a_21 n4181 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08790 n4183 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08789 vss c_15_22_s1_s n4175 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08788 c_16_20_a c_15_22_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08787 c_15_22_s1_s p_15_22_pi2j c_15_22_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08786 c_15_22_s2_s n4175 c_14_23_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08785 n4175 c_14_23_cout c_15_22_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08784 vss p_15_22_pi2j n4171 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08783 n4171 c_15_22_a n4170 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08782 n4170 c_14_23_cout n4172 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08781 vss p_15_22_pi2j n4172 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08780 n4172 c_15_22_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08779 vss n4170 c_16_21_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08778 p_15_22_pi2j c_15_22_a c_15_22_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08777 vss n4504 c_15_21_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08776 n4369 p_15_21_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08775 vss c_15_21_a n4369 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08774 n4504 c_15_21_cin n4369 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08773 n4368 p_15_21_pi2j n4504 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08772 vss c_15_21_a n4368 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08771 n4511 c_15_21_cin c_15_21_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08770 c_15_21_s2_s n4511 c_15_21_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08769 c_15_21_a p_15_21_pi2j c_15_21_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08768 c_15_21_s1_s c_15_21_a p_15_21_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08767 c_16_19_a c_15_21_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08766 vss c_15_21_s1_s n4511 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08765 n4514 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08764 vss a_19 n4371 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08763 n4371 p_15_2_d2j n4516 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08762 n4516 p_15_2_d2jbar n4370 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08761 n4370 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08760 vss p_15_21_t_s p_15_21_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08759 p_15_21_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08758 n4516 n4514 p_15_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08757 p_15_21_t_s n4516 n4514 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08756 n4928 p_15_2_d2j n4929 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08755 n4927 p_15_2_d2jbar n4928 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08754 p_15_20_t_s n4928 n4925 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08753 n4928 n4925 p_15_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08752 p_15_20_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08751 vss p_15_20_t_s p_15_20_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08750 n4925 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08749 vss a_19 n4927 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08748 n4929 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08747 vss c_15_20_s1_s n4921 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08746 c_16_18_a c_15_20_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08745 c_15_20_s1_s p_15_20_pi2j c_15_20_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08744 c_15_20_s2_s n4921 c_14_21_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08743 n4921 c_14_21_cout c_15_20_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08742 vss p_15_20_pi2j n4917 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08741 n4917 c_15_20_a n4918 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08740 n4918 c_14_21_cout n4916 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08739 vss p_15_20_pi2j n4916 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08738 n4916 c_15_20_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08737 vss n4918 c_16_19_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08736 p_15_20_pi2j c_15_20_a c_15_20_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08735 vss n5249 c_15_19_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08734 n5110 p_15_19_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08733 vss c_15_19_a n5110 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08732 n5249 c_15_19_cin n5110 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08731 n5109 p_15_19_pi2j n5249 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08730 vss c_15_19_a n5109 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08729 n5257 c_15_19_cin c_15_19_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08728 c_15_19_s2_s n5257 c_15_19_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08727 c_15_19_a p_15_19_pi2j c_15_19_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08726 c_15_19_s1_s c_15_19_a p_15_19_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08725 c_16_17_a c_15_19_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08724 vss c_15_19_s1_s n5257 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08723 n5260 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08722 vss a_17 n5112 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08721 n5112 p_15_2_d2j n5261 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08720 n5261 p_15_2_d2jbar n5111 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08719 n5111 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08718 vss p_15_19_t_s p_15_19_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08717 p_15_19_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08716 n5261 n5260 p_15_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08715 p_15_19_t_s n5261 n5260 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08714 n5681 p_15_2_d2j n5682 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08713 n5680 p_15_2_d2jbar n5681 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08712 p_15_18_t_s n5681 n5678 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08711 n5681 n5678 p_15_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08710 p_15_18_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08709 vss p_15_18_t_s p_15_18_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08708 n5678 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08707 vss a_17 n5680 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08706 n5682 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08705 vss c_15_18_s1_s n5521 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08704 c_16_16_a c_15_18_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08703 c_15_18_s1_s p_15_18_pi2j c_15_18_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08702 c_15_18_s2_s n5521 c_14_19_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08701 n5521 c_14_19_cout c_15_18_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08700 vss p_15_18_pi2j n5670 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08699 n5670 c_15_18_a n5672 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08698 n5672 c_14_19_cout n5671 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08697 vss p_15_18_pi2j n5671 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08696 n5671 c_15_18_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08695 vss n5672 c_16_17_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08694 p_15_18_pi2j c_15_18_a c_15_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08693 vss n6029 c_15_17_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08692 n5872 p_15_17_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08691 vss c_15_17_a n5872 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08690 n6029 c_15_17_cin n5872 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08689 n5669 p_15_17_pi2j n6029 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08688 vss c_15_17_a n5669 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08687 n6023 c_15_17_cin c_15_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08686 c_15_17_s2_s n6023 c_15_17_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08685 c_15_17_a p_15_17_pi2j c_15_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08684 c_15_17_s1_s c_15_17_a p_15_17_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08683 c_16_15_a c_15_17_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08682 vss c_15_17_s1_s n6023 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08681 n6038 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08680 vss a_15 n5875 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08679 n5875 p_15_2_d2j n6037 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08678 n6037 p_15_2_d2jbar n5876 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08677 n5876 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08676 vss p_15_17_t_s p_15_17_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08675 p_15_17_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08674 n6037 n6038 p_15_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08673 p_15_17_t_s n6037 n6038 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08672 n6325 p_15_2_d2j n6326 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08671 n6324 p_15_2_d2jbar n6325 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08670 p_15_16_t_s n6325 n6468 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08669 n6325 n6468 p_15_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08668 c_15_16_b p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08667 vss p_15_16_t_s c_15_16_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08666 n6468 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08665 vss a_15 n6324 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08664 n6326 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08663 vss c_15_16_s1_s n6323 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08662 c_16_14_a c_15_16_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08661 c_15_16_s1_s c_15_16_b c_15_16_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08660 c_15_16_s2_s n6323 c_14_17_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08659 n6323 c_14_17_cout c_15_16_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08658 vss c_15_16_b n6461 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08657 n6461 c_15_16_a n6462 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08656 n6462 c_14_17_cout n6460 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08655 vss c_15_16_b n6460 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08654 n6460 c_15_16_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08653 vss n6462 c_16_15_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08652 c_15_16_b c_15_16_a c_15_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08651 vss n6854 c_15_15_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08650 n6459 c_15_15_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08649 vss c_15_15_a n6459 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08648 n6854 c_15_15_cin n6459 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08647 n6458 c_15_15_b n6854 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08646 vss c_15_15_a n6458 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08645 n6669 c_15_15_cin c_15_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08644 c_15_15_s2_s n6669 c_15_15_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08643 c_15_15_a c_15_15_b c_15_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08642 c_15_15_s1_s c_15_15_a c_15_15_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08641 c_16_13_a c_15_15_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08640 vss c_15_15_s1_s n6669 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08639 n6861 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08638 vss a_13 n6469 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08637 n6469 p_15_2_d2j n6672 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08636 n6672 p_15_2_d2jbar n6470 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08635 n6470 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08634 vss p_15_15_t_s c_15_15_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08633 c_15_15_b p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08632 n6672 n6861 p_15_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08631 p_15_15_t_s n6672 n6861 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08630 n7099 p_15_2_d2j n7100 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08629 n7098 p_15_2_d2jbar n7099 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08628 p_15_14_t_s n7099 n7097 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08627 n7099 n7097 p_15_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08626 p_15_14_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08625 vss p_15_14_t_s p_15_14_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08624 n7097 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08623 vss a_13 n7098 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08622 n7100 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08621 vss c_15_14_s1_s n7094 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08620 c_16_12_a c_15_14_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08619 c_15_14_s1_s p_15_14_pi2j c_15_14_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08618 c_15_14_s2_s n7094 c_14_15_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08617 n7094 c_14_15_cout c_15_14_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08616 vss p_15_14_pi2j n7261 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08615 n7261 c_15_14_a n7091 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08614 n7091 c_14_15_cout n7262 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08613 vss p_15_14_pi2j n7262 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08612 n7262 c_15_14_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08611 vss n7091 c_16_13_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08610 p_15_14_pi2j c_15_14_a c_15_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08609 vss n7434 c_15_13_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08608 n7260 c_15_13_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08607 vss c_15_13_a n7260 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08606 n7434 c_15_13_cin n7260 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08605 n7259 c_15_13_b n7434 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08604 vss c_15_13_a n7259 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08603 n7440 c_15_13_cin c_15_13_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08602 c_15_13_s2_s n7440 c_15_13_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08601 c_15_13_a c_15_13_b c_15_13_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08600 c_15_13_s1_s c_15_13_a c_15_13_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08599 c_16_11_a c_15_13_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08598 vss c_15_13_s1_s n7440 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08597 n7443 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08596 vss a_11 n7267 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08595 n7267 p_15_2_d2j n7445 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08594 n7445 p_15_2_d2jbar n7266 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08593 n7266 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08592 vss p_15_13_t_s c_15_13_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08591 c_15_13_b p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08590 n7445 n7443 p_15_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08589 p_15_13_t_s n7445 n7443 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08588 n7872 p_15_2_d2j n7873 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08587 n7871 p_15_2_d2jbar n7872 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08586 p_15_12_t_s n7872 n7869 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08585 n7872 n7869 p_15_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08584 c_15_12_b p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08583 vss p_15_12_t_s c_15_12_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08582 n7869 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08581 vss a_11 n7871 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08580 n7873 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08579 vss c_15_12_s1_s n7866 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08578 c_16_10_a c_15_12_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08577 c_15_12_s1_s c_15_12_b c_15_12_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08576 c_15_12_s2_s n7866 c_14_13_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08575 n7866 c_14_13_cout c_15_12_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08574 vss c_15_12_b n7862 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08573 n7862 c_15_12_a n7863 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08572 n7863 c_14_13_cout n7861 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08571 vss c_15_12_b n7861 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08570 n7861 c_15_12_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08569 vss n7863 c_16_11_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08568 c_15_12_b c_15_12_a c_15_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08567 vss n8193 c_15_11_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08566 n8048 p_15_11_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08565 vss c_15_11_a n8048 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08564 n8193 c_15_11_cin n8048 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08563 n8047 p_15_11_pi2j n8193 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08562 vss c_15_11_a n8047 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08561 n8196 c_15_11_cin c_15_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08560 c_15_11_s2_s n8196 c_15_11_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08559 c_15_11_a p_15_11_pi2j c_15_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08558 c_15_11_s1_s c_15_11_a p_15_11_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08557 c_16_9_a c_15_11_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08556 vss c_15_11_s1_s n8196 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08555 n8202 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08554 vss a_9 n8051 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08553 n8051 p_15_2_d2j n8204 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08552 n8204 p_15_2_d2jbar n8050 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08551 n8050 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08550 vss p_15_11_t_s p_15_11_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08549 p_15_11_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08548 n8204 n8202 p_15_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08547 p_15_11_t_s n8204 n8202 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08546 n8617 p_15_2_d2j n8618 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08545 n8616 p_15_2_d2jbar n8617 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08544 p_15_10_t_s n8617 n8615 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08543 n8617 n8615 p_15_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08542 p_15_10_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08541 vss p_15_10_t_s p_15_10_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08540 n8615 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08539 vss a_9 n8616 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08538 n8618 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08537 vss c_15_10_s1_s n8610 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08536 c_16_8_a c_15_10_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08535 c_15_10_s1_s p_15_10_pi2j c_15_10_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08534 c_15_10_s2_s n8610 c_14_11_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08533 n8610 c_14_11_cout c_15_10_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08532 vss p_15_10_pi2j n8607 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08531 n8607 c_15_10_a n8605 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08530 n8605 c_14_11_cout n8606 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08529 vss p_15_10_pi2j n8606 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08528 n8606 c_15_10_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08527 vss n8605 c_16_9_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08526 p_15_10_pi2j c_15_10_a c_15_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08525 vss n8937 c_15_9_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08524 n8802 p_15_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08523 vss c_15_9_a n8802 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08522 n8937 c_15_9_cin n8802 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08521 n8801 p_15_9_pi2j n8937 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08520 vss c_15_9_a n8801 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08519 n8945 c_15_9_cin c_15_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08518 c_15_9_s2_s n8945 c_15_9_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08517 c_15_9_a p_15_9_pi2j c_15_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08516 c_15_9_s1_s c_15_9_a p_15_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08515 c_16_7_a c_15_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08514 vss c_15_9_s1_s n8945 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08513 n8948 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08512 vss a_7 n8804 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08511 n8804 p_15_2_d2j n8950 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08510 n8950 p_15_2_d2jbar n8803 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08509 n8803 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08508 vss p_15_9_t_s p_15_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08507 p_15_9_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08506 n8950 n8948 p_15_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08505 p_15_9_t_s n8950 n8948 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08504 n9352 p_15_2_d2j n9353 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08503 n9351 p_15_2_d2jbar n9352 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08502 p_15_8_t_s n9352 n9349 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08501 n9352 n9349 p_15_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08500 p_15_8_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08499 vss p_15_8_t_s p_15_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08498 n9349 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08497 vss a_7 n9351 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08496 n9353 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08495 vss c_15_8_s1_s n9343 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08494 c_16_6_a c_15_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08493 c_15_8_s1_s p_15_8_pi2j c_15_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08492 c_15_8_s2_s n9343 c_14_9_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08491 n9343 c_14_9_cout c_15_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08490 vss p_15_8_pi2j n9340 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08489 n9340 c_15_8_a n9341 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08488 n9341 c_14_9_cout n9342 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08487 vss p_15_8_pi2j n9342 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08486 n9342 c_15_8_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08485 vss n9341 c_16_7_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08484 p_15_8_pi2j c_15_8_a c_15_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08483 vss n9711 c_15_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08482 n9550 p_15_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08481 vss c_15_7_a n9550 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08480 n9711 c_15_7_cin n9550 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08479 n9339 p_15_7_pi2j n9711 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08478 vss c_15_7_a n9339 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08477 n9717 c_15_7_cin c_15_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08476 c_15_7_s2_s n9717 c_15_7_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08475 c_15_7_a p_15_7_pi2j c_15_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08474 c_15_7_s1_s c_15_7_a p_15_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08473 c_16_5_a c_15_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08472 vss c_15_7_s1_s n9717 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08471 n9722 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08470 vss a_5 n9554 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08469 n9554 p_15_2_d2j n9721 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08468 n9721 p_15_2_d2jbar n9553 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08467 n9553 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08466 vss p_15_7_t_s p_15_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08465 p_15_7_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08464 n9721 n9722 p_15_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08463 p_15_7_t_s n9721 n9722 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08462 n10132 p_15_2_d2j n10004 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08461 n10003 p_15_2_d2jbar n10132 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08460 p_15_6_t_s n10132 n10133 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08459 n10132 n10133 p_15_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08458 c_15_6_b p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_08457 vss p_15_6_t_s c_15_6_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_08456 n10133 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08455 vss a_5 n10003 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08454 n10004 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08453 vss c_15_6_s1_s n10002 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08452 c_16_4_a c_15_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08451 c_15_6_s1_s c_15_6_b c_15_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08450 c_15_6_s2_s n10002 c_14_7_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08449 n10002 c_14_7_cout c_15_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08448 vss c_15_6_b n10124 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08447 n10124 c_15_6_a n10125 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08446 n10125 c_14_7_cout n10123 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08445 vss c_15_6_b n10123 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08444 n10123 c_15_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08443 vss n10125 c_16_5_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08442 c_15_6_b c_15_6_a c_15_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08441 vss n10523 c_15_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08440 n10339 c_15_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08439 vss c_15_5_a n10339 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08438 n10523 c_15_5_cin n10339 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08437 n10122 c_15_5_b n10523 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08436 vss c_15_5_a n10122 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08435 n10343 c_15_5_cin c_15_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08434 c_15_5_s2_s n10343 c_15_5_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08433 c_15_5_a c_15_5_b c_15_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08432 c_15_5_s1_s c_15_5_a c_15_5_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08431 c_16_3_a c_15_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08430 vss c_15_5_s1_s n10343 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08429 n10532 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08428 vss a_3 n10134 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08427 n10134 p_15_2_d2j n10530 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08426 n10530 p_15_2_d2jbar n10135 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08425 n10135 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08424 vss p_15_5_t_s c_15_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_08423 c_15_5_b p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_08422 n10530 n10532 p_15_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08421 p_15_5_t_s n10530 n10532 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08420 n10773 p_15_2_d2j n10774 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08419 n10772 p_15_2_d2jbar n10773 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08418 p_15_4_t_s n10773 n10771 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08417 n10773 n10771 p_15_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08416 p_15_4_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08415 vss p_15_4_t_s p_15_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08414 n10771 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08413 vss a_3 n10772 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08412 n10774 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08411 vss c_15_4_s1_s n10768 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08410 c_16_2_a c_15_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08409 c_15_4_s1_s p_15_4_pi2j c_15_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08408 c_15_4_s2_s n10768 c_14_5_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08407 n10768 c_14_5_cout c_15_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08406 vss p_15_4_pi2j n10929 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08405 n10929 c_15_4_a n10765 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08404 n10765 c_14_5_cout n10930 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08403 vss p_15_4_pi2j n10930 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08402 n10930 c_15_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08401 vss n10765 c_16_3_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08400 p_15_4_pi2j c_15_4_a c_15_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08399 vss n11099 c_15_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08398 n10928 c_15_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08397 vss c_15_3_a n10928 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08396 n11099 c_15_3_cin n10928 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08395 n10927 c_15_3_b n11099 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08394 vss c_15_3_a n10927 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08393 n11105 c_15_3_cin c_15_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08392 c_15_3_s2_s n11105 c_15_3_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08391 c_15_3_a c_15_3_b c_15_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08390 c_15_3_s1_s c_15_3_a c_15_3_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08389 c_16_1_a c_15_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08388 vss c_15_3_s1_s n11105 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08387 n11108 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08386 vss a_1 n10935 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08385 n10935 p_15_2_d2j n11110 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08384 n11110 p_15_2_d2jbar n10934 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08383 n10934 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08382 vss p_15_3_t_s c_15_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_08381 c_15_3_b p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_08380 n11110 n11108 p_15_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08379 p_15_3_t_s n11110 n11108 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08378 n11535 p_15_2_d2j n11536 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08377 n11534 p_15_2_d2jbar n11535 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08376 p_15_2_t_s n11535 n11532 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08375 n11535 n11532 p_15_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08374 c_15_2_b p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_08373 vss p_15_2_t_s c_15_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_08372 n11532 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08371 vss a_1 n11534 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08370 n11536 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08369 vss c_15_2_s1_s n11529 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08368 c_15_2_sum c_15_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08367 c_15_2_s1_s c_15_2_b c_15_2_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08366 c_15_2_s2_s n11529 c_14_3_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08365 n11529 c_14_3_cout c_15_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08364 vss c_15_2_b n11525 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08363 n11525 c_15_2_a n11526 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08362 n11526 c_14_3_cout n11524 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08361 vss c_15_2_b n11524 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08360 n11524 c_15_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08359 vss n11526 c_16_1_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08358 c_15_2_b c_15_2_a c_15_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08357 vss n11850 c_15_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08356 n11710 p_15_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08355 vss c_15_1_a n11710 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08354 n11850 c_15_1_cin n11710 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08353 n11709 p_15_1_pi2j n11850 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08352 vss c_15_1_a n11709 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08351 n11856 c_15_1_cin c_15_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08350 c_15_1_s2_s n11856 c_15_1_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08349 c_15_1_a p_15_1_pi2j c_15_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08348 c_15_1_s1_s c_15_1_a p_15_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08347 c_15_1_sum c_15_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08346 vss c_15_1_s1_s n11856 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08345 n11860 p_15_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08344 n11864 p_15_2_d2jbar n11713 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08343 n11713 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08342 vss p_15_1_t_s p_15_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08341 p_15_1_pi2j p_15_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08340 n11864 n11860 p_15_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08339 p_15_1_t_s n11864 n11860 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08338 cl4_15_s1_s n12236 c_14_1_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08337 n12236 c_14_1_sum cl4_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08336 vss cl4_15_s1_s p_22 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_08335 vss c_14_1_sum n12226 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08334 n12226 n12236 n12227 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08333 n12228 n12227 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_08332 n12225 c_14_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_08331 vss c_14_2_sum n12225 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_08330 n12222 c_14_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08329 n12223 c_14_1_cout n12222 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08328 n12220 c_14_1_sum n12223 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08327 n12225 n12236 n12220 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08326 n12221 n12223 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_08325 cl4_15_s2_s c_14_1_cout c_14_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08324 c_14_1_cout c_14_2_sum cl4_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08323 vss cl4_15_s2_s n12219 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08322 cl4_15_s3_s n12219 n12228 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08321 n12219 n12228 cl4_15_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08320 vss cl4_15_s3_s p_23 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_08319 vss c_14_33_s1_s n107 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08318 c_15_31_a c_14_33_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08317 c_14_33_s1_s c_14_31_a p_14_33_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08316 c_14_31_a p_14_33_pi2j c_14_33_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08315 c_14_33_s2_s n107 c_14_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08314 n107 c_14_32_cin c_14_33_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08313 vss c_14_31_a n13 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_08312 n13 p_14_33_pi2j n106 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08311 n106 c_14_32_cin n14 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08310 vss c_14_31_a n14 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_08309 n14 p_14_33_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08308 vss n106 c_15_32_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08307 n115 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08306 n117 a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08305 vss p_14_33_t_s p_14_33_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08304 p_14_33_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08303 n117 n115 p_14_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08302 p_14_33_t_s n117 n115 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08301 n464 p_14_2_d2j n463 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08300 n462 p_14_2_d2jbar n464 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08299 p_14_32_t_s n464 n460 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08298 n464 n460 p_14_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08297 p_14_32_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08296 vss p_14_32_t_s p_14_32_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08295 n460 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08294 vss a_31 n462 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08293 n463 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08292 vss c_14_32_s1_s n457 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08291 c_15_30_a c_14_32_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08290 c_14_32_s1_s p_14_32_pi2j c_14_31_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08289 c_14_32_s2_s n457 c_14_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08288 n457 c_14_32_cin c_14_32_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08287 vss p_14_32_pi2j n453 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08286 n453 c_14_31_a n452 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08285 n452 c_14_32_cin n454 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08284 vss p_14_32_pi2j n454 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08283 n454 c_14_31_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08282 vss n452 c_15_31_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08281 p_14_32_pi2j c_14_31_a c_14_32_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08280 vss n779 c_14_31_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08279 n622 p_14_31_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08278 vss c_14_31_a n622 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08277 n779 c_14_31_cin n622 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08276 n621 p_14_31_pi2j n779 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08275 vss c_14_31_a n621 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08274 n775 c_14_31_cin c_14_31_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08273 c_14_31_s2_s n775 c_14_31_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08272 c_14_31_a p_14_31_pi2j c_14_31_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08271 c_14_31_s1_s c_14_31_a p_14_31_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08270 c_15_29_a c_14_31_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08269 vss c_14_31_s1_s n775 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08268 n785 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08267 vss a_29 n623 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08266 n623 p_14_2_d2j n788 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08265 n788 p_14_2_d2jbar n624 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08264 n624 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08263 vss p_14_31_t_s p_14_31_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08262 p_14_31_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08261 n788 n785 p_14_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08260 p_14_31_t_s n788 n785 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08259 n1210 p_14_2_d2j n1209 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08258 n1211 p_14_2_d2jbar n1210 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08257 p_14_30_t_s n1210 n1208 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08256 n1210 n1208 p_14_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08255 p_14_30_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08254 vss p_14_30_t_s p_14_30_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08253 n1208 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08252 vss a_29 n1211 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08251 n1209 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08250 vss c_14_30_s1_s n1204 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08249 c_15_28_a c_14_30_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08248 c_14_30_s1_s p_14_30_pi2j c_14_30_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08247 c_14_30_s2_s n1204 c_12_31_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08246 n1204 c_12_31_cout c_14_30_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08245 vss p_14_30_pi2j n1200 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08244 n1200 c_14_30_a n1198 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08243 n1198 c_12_31_cout n1199 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08242 vss p_14_30_pi2j n1199 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08241 n1199 c_14_30_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08240 vss n1198 c_15_29_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08239 p_14_30_pi2j c_14_30_a c_14_30_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08238 vss n1546 c_14_29_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08237 n1391 p_14_29_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08236 vss c_14_29_a n1391 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08235 n1546 c_14_29_cin n1391 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08234 n1197 p_14_29_pi2j n1546 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08233 vss c_14_29_a n1197 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08232 n1541 c_14_29_cin c_14_29_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08231 c_14_29_s2_s n1541 c_14_29_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08230 c_14_29_a p_14_29_pi2j c_14_29_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08229 c_14_29_s1_s c_14_29_a p_14_29_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08228 c_15_27_a c_14_29_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08227 vss c_14_29_s1_s n1541 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08226 n1553 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08225 vss a_27 n1392 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08224 n1392 p_14_2_d2j n1554 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08223 n1554 p_14_2_d2jbar n1393 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08222 n1393 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08221 vss p_14_29_t_s p_14_29_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08220 p_14_29_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08219 n1554 n1553 p_14_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08218 p_14_29_t_s n1554 n1553 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08217 n1970 p_14_2_d2j n1968 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08216 n1969 p_14_2_d2jbar n1970 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08215 p_14_28_t_s n1970 n1967 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08214 n1970 n1967 p_14_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08213 p_14_28_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08212 vss p_14_28_t_s p_14_28_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08211 n1967 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08210 vss a_27 n1969 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08209 n1968 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08208 vss c_14_28_s1_s n1802 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08207 c_15_26_a c_14_28_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08206 c_14_28_s1_s p_14_28_pi2j c_14_28_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08205 c_14_28_s2_s n1802 c_12_29_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08204 n1802 c_12_29_cout c_14_28_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08203 vss p_14_28_pi2j n1959 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08202 n1959 c_14_28_a n1958 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08201 n1958 c_12_29_cout n1960 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08200 vss p_14_28_pi2j n1960 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08199 n1960 c_14_28_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08198 vss n1958 c_15_27_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08197 p_14_28_pi2j c_14_28_a c_14_28_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08196 vss n2358 c_14_27_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08195 n2162 c_14_27_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08194 vss c_14_27_a n2162 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08193 n2358 c_14_27_cin n2162 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08192 n1957 c_14_27_b n2358 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08191 vss c_14_27_a n1957 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08190 n2351 c_14_27_cin c_14_27_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08189 c_14_27_s2_s n2351 c_14_27_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08188 c_14_27_a c_14_27_b c_14_27_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08187 c_14_27_s1_s c_14_27_a c_14_27_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08186 c_15_25_a c_14_27_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08185 vss c_14_27_s1_s n2351 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08184 n2363 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08183 vss a_25 n2167 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08182 n2167 p_14_2_d2j n2359 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08181 n2359 p_14_2_d2jbar n2168 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08180 n2168 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08179 vss p_14_27_t_s c_14_27_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08178 c_14_27_b p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08177 n2359 n2363 p_14_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08176 p_14_27_t_s n2359 n2363 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08175 n2627 p_14_2_d2j n2626 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08174 n2625 p_14_2_d2jbar n2627 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08173 p_14_26_t_s n2627 n2624 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08172 n2627 n2624 p_14_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08171 p_14_26_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08170 vss p_14_26_t_s p_14_26_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08169 n2624 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08168 vss a_25 n2625 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08167 n2626 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08166 vss c_14_26_s1_s n2623 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08165 c_15_24_a c_14_26_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08164 c_14_26_s1_s p_14_26_pi2j c_14_26_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08163 c_14_26_s2_s n2623 c_12_27_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08162 n2623 c_12_27_cout c_14_26_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08161 vss p_14_26_pi2j n2785 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08160 n2785 c_14_26_a n2784 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08159 n2784 c_12_27_cout n2786 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08158 vss p_14_26_pi2j n2786 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08157 n2786 c_14_26_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08156 vss n2784 c_15_25_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08155 p_14_26_pi2j c_14_26_a c_14_26_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08154 vss n3170 c_14_25_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08153 n2783 c_14_25_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08152 vss c_14_25_a n2783 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08151 n3170 c_14_25_cin n2783 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08150 n2782 c_14_25_b n3170 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08149 vss c_14_25_a n2782 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08148 n2975 c_14_25_cin c_14_25_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08147 c_14_25_s2_s n2975 c_14_25_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08146 c_14_25_a c_14_25_b c_14_25_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08145 c_14_25_s1_s c_14_25_a c_14_25_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08144 c_15_23_a c_14_25_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08143 vss c_14_25_s1_s n2975 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08142 n3176 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08141 vss a_23 n2792 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08140 n2792 p_14_2_d2j n2981 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08139 n2981 p_14_2_d2jbar n2793 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08138 n2793 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08137 vss p_14_25_t_s c_14_25_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08136 c_14_25_b p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08135 n2981 n3176 p_14_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08134 p_14_25_t_s n2981 n3176 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08133 n3407 p_14_2_d2j n3406 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08132 n3405 p_14_2_d2jbar n3407 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08131 p_14_24_t_s n3407 n3404 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08130 n3407 n3404 p_14_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08129 c_14_24_b p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08128 vss p_14_24_t_s c_14_24_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08127 n3404 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08126 vss a_23 n3405 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08125 n3406 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08124 vss c_14_24_s1_s n3401 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08123 c_15_22_a c_14_24_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08122 c_14_24_s1_s c_14_24_b c_14_24_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08121 c_14_24_s2_s n3401 c_12_25_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08120 n3401 c_12_25_cout c_14_24_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08119 vss c_14_24_b n3571 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08118 n3571 c_14_24_a n3397 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08117 n3397 c_12_25_cout n3570 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08116 vss c_14_24_b n3570 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08115 n3570 c_14_24_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08114 vss n3397 c_15_23_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08113 c_14_24_b c_14_24_a c_14_24_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08112 vss n3759 c_14_23_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08111 n3569 c_14_23_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08110 vss c_14_23_a n3569 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08109 n3759 c_14_23_cin n3569 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08108 n3568 c_14_23_b n3759 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08107 vss c_14_23_a n3568 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08106 n3762 c_14_23_cin c_14_23_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08105 c_14_23_s2_s n3762 c_14_23_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08104 c_14_23_a c_14_23_b c_14_23_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08103 c_14_23_s1_s c_14_23_a c_14_23_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08102 c_15_21_a c_14_23_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08101 vss c_14_23_s1_s n3762 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08100 n3767 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08099 vss a_21 n3574 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08098 n3574 p_14_2_d2j n3770 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08097 n3770 p_14_2_d2jbar n3575 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08096 n3575 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08095 vss p_14_23_t_s c_14_23_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08094 c_14_23_b p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08093 n3770 n3767 p_14_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08092 p_14_23_t_s n3770 n3767 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08091 n4197 p_14_2_d2j n4196 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08090 n4195 p_14_2_d2jbar n4197 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08089 p_14_22_t_s n4197 n4194 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08088 n4197 n4194 p_14_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08087 p_14_22_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08086 vss p_14_22_t_s p_14_22_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08085 n4194 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08084 vss a_21 n4195 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08083 n4196 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08082 vss c_14_22_s1_s n4189 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08081 c_15_20_a c_14_22_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08080 c_14_22_s1_s p_14_22_pi2j c_14_22_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08079 c_14_22_s2_s n4189 c_12_23_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08078 n4189 c_12_23_cout c_14_22_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08077 vss p_14_22_pi2j n4185 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08076 n4185 c_14_22_a n4184 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08075 n4184 c_12_23_cout n4186 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08074 vss p_14_22_pi2j n4186 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08073 n4186 c_14_22_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08072 vss n4184 c_15_21_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08071 p_14_22_pi2j c_14_22_a c_14_22_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08070 vss n4524 c_14_21_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08069 n4373 p_14_21_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08068 vss c_14_21_a n4373 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08067 n4524 c_14_21_cin n4373 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08066 n4372 p_14_21_pi2j n4524 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08065 vss c_14_21_a n4372 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08064 n4520 c_14_21_cin c_14_21_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08063 c_14_21_s2_s n4520 c_14_21_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08062 c_14_21_a p_14_21_pi2j c_14_21_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08061 c_14_21_s1_s c_14_21_a p_14_21_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08060 c_15_19_a c_14_21_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08059 vss c_14_21_s1_s n4520 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08058 n4532 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08057 vss a_19 n4374 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08056 n4374 p_14_2_d2j n4535 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08055 n4535 p_14_2_d2jbar n4375 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08054 n4375 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08053 vss p_14_21_t_s p_14_21_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08052 p_14_21_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08051 n4535 n4532 p_14_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08050 p_14_21_t_s n4535 n4532 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08049 n4943 p_14_2_d2j n4942 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08048 n4941 p_14_2_d2jbar n4943 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08047 p_14_20_t_s n4943 n4940 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08046 n4943 n4940 p_14_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08045 p_14_20_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08044 vss p_14_20_t_s p_14_20_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08043 n4940 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08042 vss a_19 n4941 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08041 n4942 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08040 vss c_14_20_s1_s n4936 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08039 c_15_18_a c_14_20_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08038 c_14_20_s1_s p_14_20_pi2j c_14_20_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08037 c_14_20_s2_s n4936 c_12_21_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08036 n4936 c_12_21_cout c_14_20_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08035 vss p_14_20_pi2j n4931 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08034 n4931 c_14_20_a n4932 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08033 n4932 c_12_21_cout n4930 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08032 vss p_14_20_pi2j n4930 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08031 n4930 c_14_20_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08030 vss n4932 c_15_19_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08029 p_14_20_pi2j c_14_20_a c_14_20_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08028 vss n5272 c_14_19_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_08027 n5114 p_14_19_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08026 vss c_14_19_a n5114 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08025 n5272 c_14_19_cin n5114 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08024 n5113 p_14_19_pi2j n5272 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08023 vss c_14_19_a n5113 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_08022 n5268 c_14_19_cin c_14_19_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08021 c_14_19_s2_s n5268 c_14_19_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08020 c_14_19_a p_14_19_pi2j c_14_19_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08019 c_14_19_s1_s c_14_19_a p_14_19_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_08018 c_15_17_a c_14_19_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_08017 vss c_14_19_s1_s n5268 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_08016 n5280 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08015 vss a_17 n5115 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08014 n5115 p_14_2_d2j n5281 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08013 n5281 p_14_2_d2jbar n5116 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08012 n5116 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_08011 vss p_14_19_t_s p_14_19_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08010 p_14_19_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08009 n5281 n5280 p_14_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08008 p_14_19_t_s n5281 n5280 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08007 n5696 p_14_2_d2j n5694 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08006 n5695 p_14_2_d2jbar n5696 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_08005 p_14_18_t_s n5696 n5693 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08004 n5696 n5693 p_14_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08003 p_14_18_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08002 vss p_14_18_t_s p_14_18_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_08001 n5693 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_08000 vss a_17 n5695 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07999 n5694 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07998 vss c_14_18_s1_s n5528 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07997 c_15_16_a c_14_18_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07996 c_14_18_s1_s p_14_18_pi2j c_14_18_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07995 c_14_18_s2_s n5528 c_12_19_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07994 n5528 c_12_19_cout c_14_18_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07993 vss p_14_18_pi2j n5684 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07992 n5684 c_14_18_a n5686 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07991 n5686 c_12_19_cout n5685 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07990 vss p_14_18_pi2j n5685 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07989 n5685 c_14_18_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07988 vss n5686 c_15_17_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07987 p_14_18_pi2j c_14_18_a c_14_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07986 vss n6053 c_14_17_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07985 n5877 p_14_17_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07984 vss c_14_17_a n5877 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07983 n6053 c_14_17_cin n5877 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07982 n5683 p_14_17_pi2j n6053 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07981 vss c_14_17_a n5683 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07980 n6045 c_14_17_cin c_14_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07979 c_14_17_s2_s n6045 c_14_17_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07978 c_14_17_a p_14_17_pi2j c_14_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07977 c_14_17_s1_s c_14_17_a p_14_17_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07976 c_15_15_a c_14_17_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07975 vss c_14_17_s1_s n6045 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07974 n6060 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07973 vss a_15 n5881 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07972 n5881 p_14_2_d2j n6055 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07971 n6055 p_14_2_d2jbar n5880 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07970 n5880 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07969 vss p_14_17_t_s p_14_17_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07968 p_14_17_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07967 n6055 n6060 p_14_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07966 p_14_17_t_s n6055 n6060 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07965 n6333 p_14_2_d2j n6332 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07964 n6331 p_14_2_d2jbar n6333 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07963 p_14_16_t_s n6333 n6481 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07962 n6333 n6481 p_14_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07961 p_14_16_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07960 vss p_14_16_t_s p_14_16_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07959 n6481 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07958 vss a_15 n6331 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07957 n6332 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07956 vss c_14_16_s1_s n6330 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07955 c_15_14_a c_14_16_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07954 c_14_16_s1_s p_14_16_pi2j c_14_16_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07953 c_14_16_s2_s n6330 c_12_17_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07952 n6330 c_12_17_cout c_14_16_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07951 vss p_14_16_pi2j n6473 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07950 n6473 c_14_16_a n6474 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07949 n6474 c_12_17_cout n6475 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07948 vss p_14_16_pi2j n6475 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07947 n6475 c_14_16_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07946 vss n6474 c_15_15_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07945 p_14_16_pi2j c_14_16_a c_14_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07944 vss n6873 c_14_15_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07943 n6472 c_14_15_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07942 vss c_14_15_a n6472 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07941 n6873 c_14_15_cin n6472 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07940 n6471 c_14_15_b n6873 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07939 vss c_14_15_a n6471 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07938 n6676 c_14_15_cin c_14_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07937 c_14_15_s2_s n6676 c_14_15_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07936 c_14_15_a c_14_15_b c_14_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07935 c_14_15_s1_s c_14_15_a c_14_15_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07934 c_15_13_a c_14_15_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07933 vss c_14_15_s1_s n6676 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07932 n6878 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07931 vss a_13 n6482 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07930 n6482 p_14_2_d2j n6682 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07929 n6682 p_14_2_d2jbar n6483 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07928 n6483 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07927 vss p_14_15_t_s c_14_15_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07926 c_14_15_b p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07925 n6682 n6878 p_14_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07924 p_14_15_t_s n6682 n6878 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07923 n7110 p_14_2_d2j n7109 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07922 n7108 p_14_2_d2jbar n7110 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07921 p_14_14_t_s n7110 n7107 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07920 n7110 n7107 p_14_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07919 p_14_14_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07918 vss p_14_14_t_s p_14_14_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07917 n7107 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07916 vss a_13 n7108 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07915 n7109 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07914 vss c_14_14_s1_s n7104 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07913 c_15_12_a c_14_14_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07912 c_14_14_s1_s p_14_14_pi2j c_14_14_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07911 c_14_14_s2_s n7104 c_12_15_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07910 n7104 c_12_15_cout c_14_14_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07909 vss p_14_14_pi2j n7270 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07908 n7270 c_14_14_a n7101 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07907 n7101 c_12_15_cout n7271 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07906 vss p_14_14_pi2j n7271 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07905 n7271 c_14_14_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07904 vss n7101 c_15_13_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07903 p_14_14_pi2j c_14_14_a c_14_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07902 vss n7449 c_14_13_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07901 n7269 c_14_13_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07900 vss c_14_13_a n7269 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07899 n7449 c_14_13_cin n7269 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07898 n7268 c_14_13_b n7449 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07897 vss c_14_13_a n7268 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07896 n7452 c_14_13_cin c_14_13_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07895 c_14_13_s2_s n7452 c_14_13_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07894 c_14_13_a c_14_13_b c_14_13_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07893 c_14_13_s1_s c_14_13_a c_14_13_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07892 c_15_11_a c_14_13_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07891 vss c_14_13_s1_s n7452 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07890 n7456 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07889 vss a_11 n7275 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07888 n7275 p_14_2_d2j n7459 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07887 n7459 p_14_2_d2jbar n7276 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07886 n7276 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07885 vss p_14_13_t_s c_14_13_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07884 c_14_13_b p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07883 n7459 n7456 p_14_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07882 p_14_13_t_s n7459 n7456 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07881 n7886 p_14_2_d2j n7885 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07880 n7884 p_14_2_d2jbar n7886 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07879 p_14_12_t_s n7886 n7883 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07878 n7886 n7883 p_14_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07877 c_14_12_b p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07876 vss p_14_12_t_s c_14_12_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07875 n7883 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07874 vss a_11 n7884 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07873 n7885 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07872 vss c_14_12_s1_s n7879 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07871 c_15_10_a c_14_12_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07870 c_14_12_s1_s c_14_12_b c_14_12_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07869 c_14_12_s2_s n7879 c_12_13_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07868 n7879 c_12_13_cout c_14_12_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07867 vss c_14_12_b n7875 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07866 n7875 c_14_12_a n7876 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07865 n7876 c_12_13_cout n7874 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07864 vss c_14_12_b n7874 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07863 n7874 c_14_12_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07862 vss n7876 c_15_11_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07861 c_14_12_b c_14_12_a c_14_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07860 vss n8213 c_14_11_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07859 n8053 p_14_11_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07858 vss c_14_11_a n8053 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07857 n8213 c_14_11_cin n8053 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07856 n8052 p_14_11_pi2j n8213 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07855 vss c_14_11_a n8052 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07854 n8208 c_14_11_cin c_14_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07853 c_14_11_s2_s n8208 c_14_11_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07852 c_14_11_a p_14_11_pi2j c_14_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07851 c_14_11_s1_s c_14_11_a p_14_11_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07850 c_15_9_a c_14_11_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07849 vss c_14_11_s1_s n8208 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07848 n8220 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07847 vss a_9 n8055 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07846 n8055 p_14_2_d2j n8223 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07845 n8223 p_14_2_d2jbar n8056 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07844 n8056 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07843 vss p_14_11_t_s p_14_11_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07842 p_14_11_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07841 n8223 n8220 p_14_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07840 p_14_11_t_s n8223 n8220 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07839 n8632 p_14_2_d2j n8631 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07838 n8630 p_14_2_d2jbar n8632 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07837 p_14_10_t_s n8632 n8629 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07836 n8632 n8629 p_14_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07835 p_14_10_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07834 vss p_14_10_t_s p_14_10_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07833 n8629 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07832 vss a_9 n8630 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07831 n8631 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07830 vss c_14_10_s1_s n8625 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07829 c_15_8_a c_14_10_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07828 c_14_10_s1_s p_14_10_pi2j c_14_10_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07827 c_14_10_s2_s n8625 c_12_11_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07826 n8625 c_12_11_cout c_14_10_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07825 vss p_14_10_pi2j n8621 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07824 n8621 c_14_10_a n8619 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07823 n8619 c_12_11_cout n8620 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07822 vss p_14_10_pi2j n8620 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07821 n8620 c_14_10_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07820 vss n8619 c_15_9_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07819 p_14_10_pi2j c_14_10_a c_14_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07818 vss n8960 c_14_9_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07817 n8806 p_14_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07816 vss c_14_9_a n8806 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07815 n8960 c_14_9_cin n8806 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07814 n8805 p_14_9_pi2j n8960 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07813 vss c_14_9_a n8805 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07812 n8956 c_14_9_cin c_14_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07811 c_14_9_s2_s n8956 c_14_9_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07810 c_14_9_a p_14_9_pi2j c_14_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07809 c_14_9_s1_s c_14_9_a p_14_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07808 c_15_7_a c_14_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07807 vss c_14_9_s1_s n8956 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07806 n8968 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07805 vss a_7 n8807 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07804 n8807 p_14_2_d2j n8969 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07803 n8969 p_14_2_d2jbar n8808 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07802 n8808 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07801 vss p_14_9_t_s p_14_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07800 p_14_9_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07799 n8969 n8968 p_14_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07798 p_14_9_t_s n8969 n8968 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07797 n9368 p_14_2_d2j n9366 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07796 n9367 p_14_2_d2jbar n9368 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07795 p_14_8_t_s n9368 n9365 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07794 n9368 n9365 p_14_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07793 p_14_8_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07792 vss p_14_8_t_s p_14_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07791 n9365 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07790 vss a_7 n9367 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07789 n9366 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07788 vss c_14_8_s1_s n9359 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07787 c_15_6_a c_14_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07786 c_14_8_s1_s p_14_8_pi2j c_14_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07785 c_14_8_s2_s n9359 c_12_9_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07784 n9359 c_12_9_cout c_14_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07783 vss p_14_8_pi2j n9355 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07782 n9355 c_14_8_a n9357 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07781 n9357 c_12_9_cout n9356 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07780 vss p_14_8_pi2j n9356 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07779 n9356 c_14_8_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07778 vss n9357 c_15_7_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07777 p_14_8_pi2j c_14_8_a c_14_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07776 vss n9737 c_14_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07775 n9555 p_14_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07774 vss c_14_7_a n9555 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07773 n9737 c_14_7_cin n9555 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07772 n9354 p_14_7_pi2j n9737 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07771 vss c_14_7_a n9354 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07770 n9732 c_14_7_cin c_14_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07769 c_14_7_s2_s n9732 c_14_7_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07768 c_14_7_a p_14_7_pi2j c_14_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07767 c_14_7_s1_s c_14_7_a p_14_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07766 c_15_5_a c_14_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07765 vss c_14_7_s1_s n9732 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07764 n9744 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07763 vss a_5 n9558 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07762 n9558 p_14_2_d2j n9739 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07761 n9739 p_14_2_d2jbar n9559 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07760 n9559 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07759 vss p_14_7_t_s p_14_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07758 p_14_7_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07757 n9739 n9744 p_14_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07756 p_14_7_t_s n9739 n9744 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07755 n10146 p_14_2_d2j n10009 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07754 n10008 p_14_2_d2jbar n10146 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07753 p_14_6_t_s n10146 n10147 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07752 n10146 n10147 p_14_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07751 p_14_6_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07750 vss p_14_6_t_s p_14_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07749 n10147 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07748 vss a_5 n10008 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07747 n10009 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07746 vss c_14_6_s1_s n10007 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07745 c_15_4_a c_14_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07744 c_14_6_s1_s p_14_6_pi2j c_14_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07743 c_14_6_s2_s n10007 c_12_7_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07742 n10007 c_12_7_cout c_14_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07741 vss p_14_6_pi2j n10138 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07740 n10138 c_14_6_a n10139 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07739 n10139 c_12_7_cout n10140 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07738 vss p_14_6_pi2j n10140 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07737 n10140 c_14_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07736 vss n10139 c_15_5_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07735 p_14_6_pi2j c_14_6_a c_14_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07734 vss n10541 c_14_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07733 n10348 c_14_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07732 vss c_14_5_a n10348 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07731 n10541 c_14_5_cin n10348 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07730 n10137 c_14_5_b n10541 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07729 vss c_14_5_a n10137 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07728 n10351 c_14_5_cin c_14_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07727 c_14_5_s2_s n10351 c_14_5_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07726 c_14_5_a c_14_5_b c_14_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07725 c_14_5_s1_s c_14_5_a c_14_5_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07724 c_15_3_a c_14_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07723 vss c_14_5_s1_s n10351 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07722 n10549 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07721 vss a_3 n10148 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07720 n10148 p_14_2_d2j n10544 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07719 n10544 p_14_2_d2jbar n10149 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07718 n10149 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07717 vss p_14_5_t_s c_14_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_07716 c_14_5_b p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_07715 n10544 n10549 p_14_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07714 p_14_5_t_s n10544 n10549 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07713 n10784 p_14_2_d2j n10783 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07712 n10782 p_14_2_d2jbar n10784 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07711 p_14_4_t_s n10784 n10781 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07710 n10784 n10781 p_14_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07709 p_14_4_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07708 vss p_14_4_t_s p_14_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07707 n10781 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07706 vss a_3 n10782 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07705 n10783 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07704 vss c_14_4_s1_s n10779 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07703 c_15_2_a c_14_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07702 c_14_4_s1_s p_14_4_pi2j c_14_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07701 c_14_4_s2_s n10779 c_12_5_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07700 n10779 c_12_5_cout c_14_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07699 vss p_14_4_pi2j n10938 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07698 n10938 c_14_4_a n10775 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07697 n10775 c_12_5_cout n10939 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07696 vss p_14_4_pi2j n10939 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07695 n10939 c_14_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07694 vss n10775 c_15_3_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07693 p_14_4_pi2j c_14_4_a c_14_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07692 vss n11114 c_14_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07691 n10937 c_14_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07690 vss c_14_3_a n10937 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07689 n11114 c_14_3_cin n10937 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07688 n10936 c_14_3_b n11114 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07687 vss c_14_3_a n10936 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07686 n11116 c_14_3_cin c_14_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07685 c_14_3_s2_s n11116 c_14_3_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07684 c_14_3_a c_14_3_b c_14_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07683 c_14_3_s1_s c_14_3_a c_14_3_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07682 c_15_1_a c_14_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07681 vss c_14_3_s1_s n11116 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07680 n11121 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07679 vss a_1 n10943 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07678 n10943 p_14_2_d2j n11124 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07677 n11124 p_14_2_d2jbar n10944 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07676 n10944 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07675 vss p_14_3_t_s c_14_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_07674 c_14_3_b p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_07673 n11124 n11121 p_14_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07672 p_14_3_t_s n11124 n11121 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07671 n11549 p_14_2_d2j n11548 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07670 n11547 p_14_2_d2jbar n11549 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07669 p_14_2_t_s n11549 n11546 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07668 n11549 n11546 p_14_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07667 c_14_2_b p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_07666 vss p_14_2_t_s c_14_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_07665 n11546 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07664 vss a_1 n11547 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07663 n11548 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07662 vss c_14_2_s1_s n11542 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07661 c_14_2_sum c_14_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07660 c_14_2_s1_s c_14_2_b c_14_2_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07659 c_14_2_s2_s n11542 c_12_3_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07658 n11542 c_12_3_cout c_14_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07657 vss c_14_2_b n11538 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07656 n11538 c_14_2_a n11539 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07655 n11539 c_12_3_cout n11537 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07654 vss c_14_2_b n11537 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07653 n11537 c_14_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07652 vss n11539 c_15_1_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07651 c_14_2_b c_14_2_a c_14_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07650 vss n11871 c_14_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07649 n11715 p_14_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07648 vss c_14_1_a n11715 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07647 n11871 c_14_1_cin n11715 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07646 n11714 p_14_1_pi2j n11871 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07645 vss c_14_1_a n11714 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07644 n11867 c_14_1_cin c_14_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07643 c_14_1_s2_s n11867 c_14_1_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07642 c_14_1_a p_14_1_pi2j c_14_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07641 c_14_1_s1_s c_14_1_a p_14_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07640 c_14_1_sum c_14_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07639 vss c_14_1_s1_s n11867 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07638 n11880 p_14_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07637 n11883 p_14_2_d2jbar n11718 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07636 n11718 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07635 vss p_14_1_t_s p_14_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07634 p_14_1_pi2j p_14_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07633 n11883 n11880 p_14_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07632 p_14_1_t_s n11883 n11880 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07631 cl4_14_s1_s n12255 c_12_1_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07630 n12255 c_12_1_sum cl4_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07629 vss cl4_14_s1_s p_20 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_07628 vss c_12_1_sum n12245 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07627 n12245 n12255 n12244 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07626 n12243 n12244 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_07625 n12240 c_12_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_07624 vss c_12_2_sum n12240 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_07623 n12241 c_12_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07622 n12239 c_12_1_cout n12241 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07621 n12238 c_12_1_sum n12239 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07620 n12240 n12255 n12238 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07619 n12236 n12239 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_07618 cl4_14_s2_s c_12_1_cout c_12_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07617 c_12_1_cout c_12_2_sum cl4_14_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07616 vss cl4_14_s2_s n12235 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07615 cl4_14_s3_s n12235 n12243 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07614 n12235 n12243 cl4_14_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07613 vss cl4_14_s3_s p_21 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_07612 vss c_12_33_s1_s n123 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07611 c_14_31_a c_12_33_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07610 c_12_33_s1_s c_12_31_a p_12_33_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07609 c_12_31_a p_12_33_pi2j c_12_33_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07608 c_12_33_s2_s n123 c_12_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07607 n123 c_12_32_cin c_12_33_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07606 vss c_12_31_a n15 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_07605 n15 p_12_33_pi2j n122 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07604 n122 c_12_32_cin n16 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07603 vss c_12_31_a n16 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_07602 n16 p_12_33_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07601 vss n122 c_14_32_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07600 n130 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07599 n131 a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07598 vss p_12_33_t_s p_12_33_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07597 p_12_33_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07596 n131 n130 p_12_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07595 p_12_33_t_s n131 n130 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07594 n477 p_12_2_d2j n475 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07593 n476 p_12_2_d2jbar n477 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07592 p_12_32_t_s n477 n474 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07591 n477 n474 p_12_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07590 p_12_32_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07589 vss p_12_32_t_s p_12_32_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07588 n474 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07587 vss a_31 n476 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07586 n475 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07585 vss c_12_32_s1_s n470 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07584 c_14_30_a c_12_32_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07583 c_12_32_s1_s p_12_32_pi2j c_12_31_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07582 c_12_32_s2_s n470 c_12_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07581 n470 c_12_32_cin c_12_32_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07580 vss p_12_32_pi2j n465 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07579 n465 c_12_31_a n467 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07578 n467 c_12_32_cin n466 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07577 vss p_12_32_pi2j n466 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07576 n466 c_12_31_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07575 vss n467 c_14_31_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07574 p_12_32_pi2j c_12_31_a c_12_32_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07573 vss n799 c_12_31_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07572 n625 p_12_31_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07571 vss c_12_31_a n625 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07570 n799 c_12_31_cin n625 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07569 n626 p_12_31_pi2j n799 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07568 vss c_12_31_a n626 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07567 n794 c_12_31_cin c_12_31_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07566 c_12_31_s2_s n794 c_12_31_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07565 c_12_31_a p_12_31_pi2j c_12_31_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07564 c_12_31_s1_s c_12_31_a p_12_31_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07563 c_14_29_a c_12_31_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07562 vss c_12_31_s1_s n794 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07561 n803 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07560 vss a_29 n627 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07559 n627 p_12_2_d2j n805 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07558 n805 p_12_2_d2jbar n628 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07557 n628 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07556 vss p_12_31_t_s p_12_31_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07555 p_12_31_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07554 n805 n803 p_12_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07553 p_12_31_t_s n805 n803 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07552 n1226 p_12_2_d2j n1224 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07551 n1225 p_12_2_d2jbar n1226 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07550 p_12_30_t_s n1226 n1223 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07549 n1226 n1223 p_12_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07548 p_12_30_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07547 vss p_12_30_t_s p_12_30_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07546 n1223 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07545 vss a_29 n1225 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07544 n1224 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07543 vss c_12_30_s1_s n1218 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07542 c_14_28_a c_12_30_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07541 c_12_30_s1_s p_12_30_pi2j c_12_30_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07540 c_12_30_s2_s n1218 c_11_31_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07539 n1218 c_11_31_cout c_12_30_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07538 vss p_12_30_pi2j n1213 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07537 n1213 c_12_30_a n1215 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07536 n1215 c_11_31_cout n1214 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07535 vss p_12_30_pi2j n1214 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07534 n1214 c_12_30_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07533 vss n1215 c_14_29_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07532 p_12_30_pi2j c_12_30_a c_12_30_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07531 vss n1569 c_12_29_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07530 n1394 p_12_29_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07529 vss c_12_29_a n1394 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07528 n1569 c_12_29_cin n1394 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07527 n1212 p_12_29_pi2j n1569 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07526 vss c_12_29_a n1212 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07525 n1566 c_12_29_cin c_12_29_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07524 c_12_29_s2_s n1566 c_12_29_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07523 c_12_29_a p_12_29_pi2j c_12_29_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07522 c_12_29_s1_s c_12_29_a p_12_29_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07521 c_14_27_a c_12_29_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07520 vss c_12_29_s1_s n1566 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07519 n1573 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07518 vss a_27 n1395 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07517 n1395 p_12_2_d2j n1576 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07516 n1576 p_12_2_d2jbar n1396 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07515 n1396 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07514 vss p_12_29_t_s p_12_29_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07513 p_12_29_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07512 n1576 n1573 p_12_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07511 p_12_29_t_s n1576 n1573 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07510 n1984 p_12_2_d2j n1982 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07509 n1983 p_12_2_d2jbar n1984 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07508 p_12_28_t_s n1984 n1981 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07507 n1984 n1981 p_12_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07506 p_12_28_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07505 vss p_12_28_t_s p_12_28_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07504 n1981 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07503 vss a_27 n1983 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07502 n1982 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07501 vss c_12_28_s1_s n1810 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07500 c_14_26_a c_12_28_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07499 c_12_28_s1_s p_12_28_pi2j c_12_28_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07498 c_12_28_s2_s n1810 c_11_29_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07497 n1810 c_11_29_cout c_12_28_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07496 vss p_12_28_pi2j n1974 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07495 n1974 c_12_28_a n1975 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07494 n1975 c_11_29_cout n1973 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07493 vss p_12_28_pi2j n1973 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07492 n1973 c_12_28_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07491 vss n1975 c_14_27_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07490 p_12_28_pi2j c_12_28_a c_12_28_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07489 vss n2380 c_12_27_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07488 n2169 c_12_27_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07487 vss c_12_27_a n2169 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07486 n2380 c_12_27_cin n2169 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07485 n1972 c_12_27_b n2380 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07484 vss c_12_27_a n1972 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07483 n2372 c_12_27_cin c_12_27_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07482 c_12_27_s2_s n2372 c_12_27_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07481 c_12_27_a c_12_27_b c_12_27_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07480 c_12_27_s1_s c_12_27_a c_12_27_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07479 c_14_25_a c_12_27_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07478 vss c_12_27_s1_s n2372 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07477 n2383 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07476 vss a_25 n2175 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07475 n2175 p_12_2_d2j n2382 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07474 n2382 p_12_2_d2jbar n2174 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07473 n2174 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07472 vss p_12_27_t_s c_12_27_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07471 c_12_27_b p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07470 n2382 n2383 p_12_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07469 p_12_27_t_s n2382 n2383 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07468 n2634 p_12_2_d2j n2633 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07467 n2635 p_12_2_d2jbar n2634 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07466 p_12_26_t_s n2634 n2632 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07465 n2634 n2632 p_12_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07464 p_12_26_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07463 vss p_12_26_t_s p_12_26_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07462 n2632 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07461 vss a_25 n2635 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07460 n2633 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07459 vss c_12_26_s1_s n2631 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07458 c_14_24_a c_12_26_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07457 c_12_26_s1_s p_12_26_pi2j c_12_26_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07456 c_12_26_s2_s n2631 c_11_27_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07455 n2631 c_11_27_cout c_12_26_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07454 vss p_12_26_pi2j n2798 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07453 n2798 c_12_26_a n2799 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07452 n2799 c_11_27_cout n2794 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07451 vss p_12_26_pi2j n2794 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07450 n2794 c_12_26_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07449 vss n2799 c_14_25_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07448 p_12_26_pi2j c_12_26_a c_12_26_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07447 vss n3189 c_12_25_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07446 n2796 c_12_25_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07445 vss c_12_25_a n2796 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07444 n3189 c_12_25_cin n2796 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07443 n2797 c_12_25_b n3189 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07442 vss c_12_25_a n2797 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07441 n2986 c_12_25_cin c_12_25_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07440 c_12_25_s2_s n2986 c_12_25_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07439 c_12_25_a c_12_25_b c_12_25_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07438 c_12_25_s1_s c_12_25_a c_12_25_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07437 c_14_23_a c_12_25_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07436 vss c_12_25_s1_s n2986 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07435 n3191 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07434 vss a_23 n2804 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07433 n2804 p_12_2_d2j n2989 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07432 n2989 p_12_2_d2jbar n2805 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07431 n2805 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07430 vss p_12_25_t_s c_12_25_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07429 c_12_25_b p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07428 n2989 n3191 p_12_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07427 p_12_25_t_s n2989 n3191 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07426 n3417 p_12_2_d2j n3416 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07425 n3418 p_12_2_d2jbar n3417 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07424 p_12_24_t_s n3417 n3415 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07423 n3417 n3415 p_12_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07422 c_12_24_b p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07421 vss p_12_24_t_s c_12_24_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07420 n3415 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07419 vss a_23 n3418 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07418 n3416 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07417 vss c_12_24_s1_s n3412 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07416 c_14_22_a c_12_24_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07415 c_12_24_s1_s c_12_24_b c_12_24_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07414 c_12_24_s2_s n3412 c_11_25_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07413 n3412 c_11_25_cout c_12_24_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07412 vss c_12_24_b n3579 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07411 n3579 c_12_24_a n3408 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07410 n3408 c_11_25_cout n3576 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07409 vss c_12_24_b n3576 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07408 n3576 c_12_24_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07407 vss n3408 c_14_23_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07406 c_12_24_b c_12_24_a c_12_24_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07405 vss n3779 c_12_23_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07404 n3577 c_12_23_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07403 vss c_12_23_a n3577 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07402 n3779 c_12_23_cin n3577 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07401 n3578 c_12_23_b n3779 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07400 vss c_12_23_a n3578 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07399 n3780 c_12_23_cin c_12_23_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07398 c_12_23_s2_s n3780 c_12_23_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07397 c_12_23_a c_12_23_b c_12_23_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07396 c_12_23_s1_s c_12_23_a c_12_23_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07395 c_14_21_a c_12_23_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07394 vss c_12_23_s1_s n3780 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07393 n3783 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07392 vss a_21 n3582 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07391 n3582 p_12_2_d2j n3785 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07390 n3785 p_12_2_d2jbar n3583 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07389 n3583 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07388 vss p_12_23_t_s c_12_23_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07387 c_12_23_b p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07386 n3785 n3783 p_12_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07385 p_12_23_t_s n3785 n3783 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07384 n4210 p_12_2_d2j n4209 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07383 n4211 p_12_2_d2jbar n4210 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07382 p_12_22_t_s n4210 n4208 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07381 n4210 n4208 p_12_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07380 p_12_22_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07379 vss p_12_22_t_s p_12_22_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07378 n4208 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07377 vss a_21 n4211 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07376 n4209 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07375 vss c_12_22_s1_s n4203 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07374 c_14_20_a c_12_22_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07373 c_12_22_s1_s p_12_22_pi2j c_12_22_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07372 c_12_22_s2_s n4203 c_11_23_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07371 n4203 c_11_23_cout c_12_22_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07370 vss p_12_22_pi2j n4198 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07369 n4198 c_12_22_a n4200 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07368 n4200 c_11_23_cout n4199 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07367 vss p_12_22_pi2j n4199 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07366 n4199 c_12_22_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07365 vss n4200 c_14_21_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07364 p_12_22_pi2j c_12_22_a c_12_22_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07363 vss n4546 c_12_21_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07362 n4376 p_12_21_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07361 vss c_12_21_a n4376 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07360 n4546 c_12_21_cin n4376 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07359 n4377 p_12_21_pi2j n4546 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07358 vss c_12_21_a n4377 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07357 n4543 c_12_21_cin c_12_21_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07356 c_12_21_s2_s n4543 c_12_21_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07355 c_12_21_a p_12_21_pi2j c_12_21_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07354 c_12_21_s1_s c_12_21_a p_12_21_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07353 c_14_19_a c_12_21_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07352 vss c_12_21_s1_s n4543 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07351 n4550 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07350 vss a_19 n4378 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07349 n4378 p_12_2_d2j n4552 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07348 n4552 p_12_2_d2jbar n4379 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07347 n4379 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07346 vss p_12_21_t_s p_12_21_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07345 p_12_21_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07344 n4552 n4550 p_12_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07343 p_12_21_t_s n4552 n4550 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07342 n4956 p_12_2_d2j n4955 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07341 n4957 p_12_2_d2jbar n4956 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07340 p_12_20_t_s n4956 n4954 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07339 n4956 n4954 p_12_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07338 p_12_20_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07337 vss p_12_20_t_s p_12_20_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07336 n4954 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07335 vss a_19 n4957 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07334 n4955 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07333 vss c_12_20_s1_s n4951 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07332 c_14_18_a c_12_20_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07331 c_12_20_s1_s p_12_20_pi2j c_12_20_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07330 c_12_20_s2_s n4951 c_11_21_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07329 n4951 c_11_21_cout c_12_20_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07328 vss p_12_20_pi2j n4944 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07327 n4944 c_12_20_a n4946 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07326 n4946 c_11_21_cout n4945 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07325 vss p_12_20_pi2j n4945 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07324 n4945 c_12_20_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07323 vss n4946 c_14_19_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07322 p_12_20_pi2j c_12_20_a c_12_20_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07321 vss n5296 c_12_19_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07320 n5117 p_12_19_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07319 vss c_12_19_a n5117 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07318 n5296 c_12_19_cin n5117 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07317 n5118 p_12_19_pi2j n5296 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07316 vss c_12_19_a n5118 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07315 n5292 c_12_19_cin c_12_19_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07314 c_12_19_s2_s n5292 c_12_19_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07313 c_12_19_a p_12_19_pi2j c_12_19_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07312 c_12_19_s1_s c_12_19_a p_12_19_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07311 c_14_17_a c_12_19_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07310 vss c_12_19_s1_s n5292 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07309 n5300 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07308 vss a_17 n5119 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07307 n5119 p_12_2_d2j n5303 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07306 n5303 p_12_2_d2jbar n5120 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07305 n5120 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07304 vss p_12_19_t_s p_12_19_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07303 p_12_19_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07302 n5303 n5300 p_12_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07301 p_12_19_t_s n5303 n5300 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07300 n5708 p_12_2_d2j n5710 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07299 n5707 p_12_2_d2jbar n5708 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07298 p_12_18_t_s n5708 n5709 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07297 n5708 n5709 p_12_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07296 p_12_18_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07295 vss p_12_18_t_s p_12_18_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07294 n5709 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07293 vss a_17 n5707 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07292 n5710 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07291 vss c_12_18_s1_s n5536 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07290 c_14_16_a c_12_18_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07289 c_12_18_s1_s p_12_18_pi2j c_12_18_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07288 c_12_18_s2_s n5536 c_11_19_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07287 n5536 c_11_19_cout c_12_18_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07286 vss p_12_18_pi2j n5701 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07285 n5701 c_12_18_a n5699 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07284 n5699 c_11_19_cout n5700 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07283 vss p_12_18_pi2j n5700 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07282 n5700 c_12_18_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07281 vss n5699 c_14_17_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07280 p_12_18_pi2j c_12_18_a c_12_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07279 vss n6079 c_12_17_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07278 n5882 p_12_17_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07277 vss c_12_17_a n5882 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07276 n6079 c_12_17_cin n5882 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07275 n5698 p_12_17_pi2j n6079 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07274 vss c_12_17_a n5698 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07273 n6069 c_12_17_cin c_12_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07272 c_12_17_s2_s n6069 c_12_17_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07271 c_12_17_a p_12_17_pi2j c_12_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07270 c_12_17_s1_s c_12_17_a p_12_17_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07269 c_14_15_a c_12_17_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07268 vss c_12_17_s1_s n6069 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07267 n6081 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07266 vss a_15 n5885 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07265 n5885 p_12_2_d2j n6080 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07264 n6080 p_12_2_d2jbar n5886 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07263 n5886 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07262 vss p_12_17_t_s p_12_17_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07261 p_12_17_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07260 n6080 n6081 p_12_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07259 p_12_17_t_s n6080 n6081 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07258 n6339 p_12_2_d2j n6338 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07257 n6340 p_12_2_d2jbar n6339 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07256 p_12_16_t_s n6339 n6493 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07255 n6339 n6493 p_12_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07254 p_12_16_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07253 vss p_12_16_t_s p_12_16_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07252 n6493 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07251 vss a_15 n6340 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07250 n6338 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07249 vss c_12_16_s1_s n6337 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07248 c_14_14_a c_12_16_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07247 c_12_16_s1_s p_12_16_pi2j c_12_16_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07246 c_12_16_s2_s n6337 c_11_17_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07245 n6337 c_11_17_cout c_12_16_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07244 vss p_12_16_pi2j n6488 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07243 n6488 c_12_16_a n6489 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07242 n6489 c_11_17_cout n6484 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07241 vss p_12_16_pi2j n6484 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07240 n6484 c_12_16_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07239 vss n6489 c_14_15_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07238 p_12_16_pi2j c_12_16_a c_12_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07237 vss n6890 c_12_15_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07236 n6487 c_12_15_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07235 vss c_12_15_a n6487 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07234 n6890 c_12_15_cin n6487 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07233 n6486 c_12_15_b n6890 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07232 vss c_12_15_a n6486 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07231 n6687 c_12_15_cin c_12_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07230 c_12_15_s2_s n6687 c_12_15_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07229 c_12_15_a c_12_15_b c_12_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07228 c_12_15_s1_s c_12_15_a c_12_15_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07227 c_14_13_a c_12_15_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07226 vss c_12_15_s1_s n6687 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07225 n6893 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07224 vss a_13 n6495 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07223 n6495 p_12_2_d2j n6690 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07222 n6690 p_12_2_d2jbar n6496 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07221 n6496 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07220 vss p_12_15_t_s c_12_15_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07219 c_12_15_b p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07218 n6690 n6893 p_12_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07217 p_12_15_t_s n6690 n6893 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07216 n7119 p_12_2_d2j n7118 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07215 n7120 p_12_2_d2jbar n7119 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07214 p_12_14_t_s n7119 n7117 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07213 n7119 n7117 p_12_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07212 p_12_14_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07211 vss p_12_14_t_s p_12_14_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07210 n7117 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07209 vss a_13 n7120 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07208 n7118 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07207 vss c_12_14_s1_s n7114 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07206 c_14_12_a c_12_14_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07205 c_12_14_s1_s p_12_14_pi2j c_12_14_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07204 c_12_14_s2_s n7114 c_11_15_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07203 n7114 c_11_15_cout c_12_14_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07202 vss p_12_14_pi2j n7281 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07201 n7281 c_12_14_a n7111 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07200 n7111 c_11_15_cout n7277 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07199 vss p_12_14_pi2j n7277 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07198 n7277 c_12_14_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07197 vss n7111 c_14_13_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07196 p_12_14_pi2j c_12_14_a c_12_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07195 vss n7464 c_12_13_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07194 n7279 c_12_13_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07193 vss c_12_13_a n7279 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07192 n7464 c_12_13_cin n7279 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07191 n7280 c_12_13_b n7464 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07190 vss c_12_13_a n7280 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07189 n7467 c_12_13_cin c_12_13_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07188 c_12_13_s2_s n7467 c_12_13_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07187 c_12_13_a c_12_13_b c_12_13_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07186 c_12_13_s1_s c_12_13_a c_12_13_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07185 c_14_11_a c_12_13_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07184 vss c_12_13_s1_s n7467 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07183 n7469 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07182 vss a_11 n7284 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07181 n7284 p_12_2_d2j n7471 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07180 n7471 p_12_2_d2jbar n7285 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07179 n7285 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07178 vss p_12_13_t_s c_12_13_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07177 c_12_13_b p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07176 n7471 n7469 p_12_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07175 p_12_13_t_s n7471 n7469 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07174 n7898 p_12_2_d2j n7897 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07173 n7899 p_12_2_d2jbar n7898 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07172 p_12_12_t_s n7898 n7896 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07171 n7898 n7896 p_12_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07170 c_12_12_b p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07169 vss p_12_12_t_s c_12_12_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07168 n7896 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07167 vss a_11 n7899 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07166 n7897 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07165 vss c_12_12_s1_s n7892 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07164 c_14_10_a c_12_12_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07163 c_12_12_s1_s c_12_12_b c_12_12_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07162 c_12_12_s2_s n7892 c_11_13_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07161 n7892 c_11_13_cout c_12_12_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07160 vss c_12_12_b n7887 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07159 n7887 c_12_12_a n7889 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07158 n7889 c_11_13_cout n7888 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07157 vss c_12_12_b n7888 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07156 n7888 c_12_12_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07155 vss n7889 c_14_11_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07154 c_12_12_b c_12_12_a c_12_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07153 vss n8232 c_12_11_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07152 n8057 p_12_11_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07151 vss c_12_11_a n8057 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07150 n8232 c_12_11_cin n8057 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07149 n8058 p_12_11_pi2j n8232 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07148 vss c_12_11_a n8058 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07147 n8231 c_12_11_cin c_12_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07146 c_12_11_s2_s n8231 c_12_11_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07145 c_12_11_a p_12_11_pi2j c_12_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07144 c_12_11_s1_s c_12_11_a p_12_11_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07143 c_14_9_a c_12_11_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07142 vss c_12_11_s1_s n8231 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07141 n8238 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07140 vss a_9 n8060 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07139 n8060 p_12_2_d2j n8240 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07138 n8240 p_12_2_d2jbar n8061 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07137 n8061 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07136 vss p_12_11_t_s p_12_11_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07135 p_12_11_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07134 n8240 n8238 p_12_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07133 p_12_11_t_s n8240 n8238 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07132 n8645 p_12_2_d2j n8644 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07131 n8646 p_12_2_d2jbar n8645 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07130 p_12_10_t_s n8645 n8643 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07129 n8645 n8643 p_12_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07128 p_12_10_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07127 vss p_12_10_t_s p_12_10_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07126 n8643 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07125 vss a_9 n8646 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07124 n8644 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07123 vss c_12_10_s1_s n8638 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07122 c_14_8_a c_12_10_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07121 c_12_10_s1_s p_12_10_pi2j c_12_10_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07120 c_12_10_s2_s n8638 c_11_11_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07119 n8638 c_11_11_cout c_12_10_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07118 vss p_12_10_pi2j n8633 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07117 n8633 c_12_10_a n8635 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07116 n8635 c_11_11_cout n8634 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07115 vss p_12_10_pi2j n8634 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07114 n8634 c_12_10_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07113 vss n8635 c_14_9_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07112 p_12_10_pi2j c_12_10_a c_12_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07111 vss n8984 c_12_9_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07110 n8809 p_12_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07109 vss c_12_9_a n8809 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07108 n8984 c_12_9_cin n8809 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07107 n8810 p_12_9_pi2j n8984 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07106 vss c_12_9_a n8810 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07105 n8980 c_12_9_cin c_12_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07104 c_12_9_s2_s n8980 c_12_9_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07103 c_12_9_a p_12_9_pi2j c_12_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07102 c_12_9_s1_s c_12_9_a p_12_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07101 c_14_7_a c_12_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07100 vss c_12_9_s1_s n8980 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07099 n8988 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07098 vss a_7 n8811 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07097 n8811 p_12_2_d2j n8991 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07096 n8991 p_12_2_d2jbar n8812 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07095 n8812 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07094 vss p_12_9_t_s p_12_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07093 p_12_9_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07092 n8991 n8988 p_12_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07091 p_12_9_t_s n8991 n8988 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07090 n9381 p_12_2_d2j n9383 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07089 n9380 p_12_2_d2jbar n9381 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07088 p_12_8_t_s n9381 n9382 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07087 n9381 n9382 p_12_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07086 p_12_8_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07085 vss p_12_8_t_s p_12_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07084 n9382 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07083 vss a_7 n9380 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07082 n9383 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07081 vss c_12_8_s1_s n9369 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07080 c_14_6_a c_12_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07079 c_12_8_s1_s p_12_8_pi2j c_12_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07078 c_12_8_s2_s n9369 c_11_9_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07077 n9369 c_11_9_cout c_12_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07076 vss p_12_8_pi2j n9374 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07075 n9374 c_12_8_a n9372 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07074 n9372 c_11_9_cout n9373 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07073 vss p_12_8_pi2j n9373 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07072 n9373 c_12_8_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07071 vss n9372 c_14_7_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07070 p_12_8_pi2j c_12_8_a c_12_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07069 vss n9763 c_12_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07068 n9560 p_12_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07067 vss c_12_7_a n9560 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07066 n9763 c_12_7_cin n9560 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07065 n9371 p_12_7_pi2j n9763 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07064 vss c_12_7_a n9371 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07063 n9759 c_12_7_cin c_12_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07062 c_12_7_s2_s n9759 c_12_7_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07061 c_12_7_a p_12_7_pi2j c_12_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07060 c_12_7_s1_s c_12_7_a p_12_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07059 c_14_5_a c_12_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07058 vss c_12_7_s1_s n9759 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07057 n9764 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07056 vss a_5 n9563 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07055 n9563 p_12_2_d2j n9765 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07054 n9765 p_12_2_d2jbar n9564 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07053 n9564 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07052 vss p_12_7_t_s p_12_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07051 p_12_7_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07050 n9765 n9764 p_12_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07049 p_12_7_t_s n9765 n9764 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07048 n10160 p_12_2_d2j n10013 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07047 n10014 p_12_2_d2jbar n10160 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07046 p_12_6_t_s n10160 n10159 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07045 n10160 n10159 p_12_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07044 p_12_6_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07043 vss p_12_6_t_s p_12_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07042 n10159 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07041 vss a_5 n10014 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07040 n10013 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07039 vss c_12_6_s1_s n10012 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07038 c_14_4_a c_12_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07037 c_12_6_s1_s p_12_6_pi2j c_12_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07036 c_12_6_s2_s n10012 c_11_7_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07035 n10012 c_11_7_cout c_12_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07034 vss p_12_6_pi2j n10155 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07033 n10155 c_12_6_a n10154 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07032 n10154 c_11_7_cout n10150 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07031 vss p_12_6_pi2j n10150 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07030 n10150 c_12_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07029 vss n10154 c_14_5_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07028 p_12_6_pi2j c_12_6_a c_12_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07027 vss n10562 c_12_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_07026 n10357 c_12_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07025 vss c_12_5_a n10357 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07024 n10562 c_12_5_cin n10357 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07023 n10153 c_12_5_b n10562 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07022 vss c_12_5_a n10153 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_07021 n10362 c_12_5_cin c_12_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07020 c_12_5_s2_s n10362 c_12_5_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07019 c_12_5_a c_12_5_b c_12_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07018 c_12_5_s1_s c_12_5_a c_12_5_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_07017 c_14_3_a c_12_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_07016 vss c_12_5_s1_s n10362 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_07015 n10565 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_07014 vss a_3 n10162 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07013 n10162 p_12_2_d2j n10564 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07012 n10564 p_12_2_d2jbar n10163 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07011 n10163 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_07010 vss p_12_5_t_s c_12_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_07009 c_12_5_b p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_07008 n10564 n10565 p_12_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07007 p_12_5_t_s n10564 n10565 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07006 n10793 p_12_2_d2j n10792 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07005 n10794 p_12_2_d2jbar n10793 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07004 p_12_4_t_s n10793 n10791 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07003 n10793 n10791 p_12_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_07002 p_12_4_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07001 vss p_12_4_t_s p_12_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_07000 n10791 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06999 vss a_3 n10794 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06998 n10792 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06997 vss c_12_4_s1_s n10789 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06996 c_14_2_a c_12_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06995 c_12_4_s1_s p_12_4_pi2j c_12_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06994 c_12_4_s2_s n10789 c_11_5_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06993 n10789 c_11_5_cout c_12_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06992 vss p_12_4_pi2j n10949 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06991 n10949 c_12_4_a n10785 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06990 n10785 c_11_5_cout n10945 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06989 vss p_12_4_pi2j n10945 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06988 n10945 c_12_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06987 vss n10785 c_14_3_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06986 p_12_4_pi2j c_12_4_a c_12_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06985 vss n11129 c_12_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06984 n10947 c_12_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06983 vss c_12_3_a n10947 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06982 n11129 c_12_3_cin n10947 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06981 n10948 c_12_3_b n11129 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06980 vss c_12_3_a n10948 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06979 n11132 c_12_3_cin c_12_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06978 c_12_3_s2_s n11132 c_12_3_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06977 c_12_3_a c_12_3_b c_12_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06976 c_12_3_s1_s c_12_3_a c_12_3_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06975 c_14_1_a c_12_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06974 vss c_12_3_s1_s n11132 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06973 n11134 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06972 vss a_1 n10952 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06971 n10952 p_12_2_d2j n11136 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06970 n11136 p_12_2_d2jbar n10953 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06969 n10953 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06968 vss p_12_3_t_s c_12_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06967 c_12_3_b p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06966 n11136 n11134 p_12_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06965 p_12_3_t_s n11136 n11134 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06964 n11561 p_12_2_d2j n11560 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06963 n11562 p_12_2_d2jbar n11561 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06962 p_12_2_t_s n11561 n11559 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06961 n11561 n11559 p_12_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06960 c_12_2_b p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06959 vss p_12_2_t_s c_12_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06958 n11559 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06957 vss a_1 n11562 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06956 n11560 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06955 vss c_12_2_s1_s n11555 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06954 c_12_2_sum c_12_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06953 c_12_2_s1_s c_12_2_b c_12_2_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06952 c_12_2_s2_s n11555 c_11_3_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06951 n11555 c_11_3_cout c_12_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06950 vss c_12_2_b n11550 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06949 n11550 c_12_2_a n11552 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06948 n11552 c_11_3_cout n11551 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06947 vss c_12_2_b n11551 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06946 n11551 c_12_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06945 vss n11552 c_14_1_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06944 c_12_2_b c_12_2_a c_12_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06943 vss n11894 c_12_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06942 n11719 p_12_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06941 vss c_12_1_a n11719 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06940 n11894 c_12_1_cin n11719 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06939 n11720 p_12_1_pi2j n11894 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06938 vss c_12_1_a n11720 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06937 n11890 c_12_1_cin c_12_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06936 c_12_1_s2_s n11890 c_12_1_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06935 c_12_1_a p_12_1_pi2j c_12_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06934 c_12_1_s1_s c_12_1_a p_12_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06933 c_12_1_sum c_12_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06932 vss c_12_1_s1_s n11890 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06931 n11901 p_12_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06930 n11902 p_12_2_d2jbar n11723 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06929 n11723 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06928 vss p_12_1_t_s p_12_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06927 p_12_1_pi2j p_12_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06926 n11902 n11901 p_12_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06925 p_12_1_t_s n11902 n11901 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06924 cl4_12_s1_s n12272 c_11_1_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06923 n12272 c_11_1_sum cl4_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06922 vss cl4_12_s1_s p_18 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06921 vss c_11_1_sum n12262 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06920 n12262 n12272 n12261 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06919 n12260 n12261 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_06918 n12259 c_11_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_06917 vss c_11_2_sum n12259 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_06916 n12258 c_11_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06915 n12256 c_11_1_cout n12258 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06914 n12254 c_11_1_sum n12256 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06913 n12259 n12272 n12254 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06912 n12255 n12256 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_06911 cl4_12_s2_s c_11_1_cout c_11_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06910 c_11_1_cout c_11_2_sum cl4_12_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06909 vss cl4_12_s2_s n12252 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06908 cl4_12_s3_s n12252 n12260 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06907 n12252 n12260 cl4_12_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06906 vss cl4_12_s3_s p_19 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06905 vss c_11_33_s1_s n141 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06904 c_12_31_a c_11_33_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06903 c_11_33_s1_s c_11_31_a p_11_33_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06902 c_11_31_a p_11_33_pi2j c_11_33_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06901 c_11_33_s2_s n141 c_11_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06900 n141 c_11_32_cin c_11_33_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06899 vss c_11_31_a n17 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_06898 n17 p_11_33_pi2j n133 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06897 n133 c_11_32_cin n18 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06896 vss c_11_31_a n18 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_06895 n18 p_11_33_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06894 vss n133 c_12_32_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06893 n142 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06892 n145 a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06891 vss p_11_33_t_s p_11_33_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06890 p_11_33_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06889 n145 n142 p_11_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06888 p_11_33_t_s n145 n142 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06887 n489 p_11_2_d2j n490 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06886 n488 p_11_2_d2jbar n489 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06885 p_11_32_t_s n489 n486 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06884 n489 n486 p_11_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06883 p_11_32_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06882 vss p_11_32_t_s p_11_32_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06881 n486 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06880 vss a_31 n488 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06879 n490 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06878 vss c_11_32_s1_s n484 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06877 c_12_30_a c_11_32_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06876 c_11_32_s1_s p_11_32_pi2j c_11_31_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06875 c_11_32_s2_s n484 c_11_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06874 n484 c_11_32_cin c_11_32_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06873 vss p_11_32_pi2j n479 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06872 n479 c_11_31_a n478 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06871 n478 c_11_32_cin n480 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06870 vss p_11_32_pi2j n480 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06869 n480 c_11_31_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06868 vss n478 c_12_31_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06867 p_11_32_pi2j c_11_31_a c_11_32_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06866 vss n810 c_11_31_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06865 n630 p_11_31_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06864 vss c_11_31_a n630 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06863 n810 c_11_31_cin n630 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06862 n629 p_11_31_pi2j n810 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06861 vss c_11_31_a n629 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06860 n815 c_11_31_cin c_11_31_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06859 c_11_31_s2_s n815 c_11_31_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06858 c_11_31_a p_11_31_pi2j c_11_31_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06857 c_11_31_s1_s c_11_31_a p_11_31_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06856 c_12_29_a c_11_31_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06855 vss c_11_31_s1_s n815 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06854 n821 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06853 vss a_29 n631 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06852 n631 p_11_2_d2j n823 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06851 n823 p_11_2_d2jbar n632 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06850 n632 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06849 vss p_11_31_t_s p_11_31_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06848 p_11_31_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06847 n823 n821 p_11_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06846 p_11_31_t_s n823 n821 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06845 n1241 p_11_2_d2j n1239 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06844 n1240 p_11_2_d2jbar n1241 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06843 p_11_30_t_s n1241 n1237 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06842 n1241 n1237 p_11_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06841 p_11_30_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06840 vss p_11_30_t_s p_11_30_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06839 n1237 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06838 vss a_29 n1240 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06837 n1239 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06836 vss c_11_30_s1_s n1233 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06835 c_12_28_a c_11_30_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06834 c_11_30_s1_s p_11_30_pi2j c_11_30_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06833 c_11_30_s2_s n1233 c_10_31_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06832 n1233 c_10_31_cout c_11_30_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06831 vss p_11_30_pi2j n1230 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06830 n1230 c_11_30_a n1228 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06829 n1228 c_10_31_cout n1229 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06828 vss p_11_30_pi2j n1229 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06827 n1229 c_11_30_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06826 vss n1228 c_12_29_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06825 p_11_30_pi2j c_11_30_a c_11_30_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06824 vss n1583 c_11_29_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06823 n1397 p_11_29_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06822 vss c_11_29_a n1397 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06821 n1583 c_11_29_cin n1397 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06820 n1227 p_11_29_pi2j n1583 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06819 vss c_11_29_a n1227 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06818 n1589 c_11_29_cin c_11_29_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06817 c_11_29_s2_s n1589 c_11_29_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06816 c_11_29_a p_11_29_pi2j c_11_29_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06815 c_11_29_s1_s c_11_29_a p_11_29_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06814 c_12_27_a c_11_29_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06813 vss c_11_29_s1_s n1589 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06812 n1593 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06811 vss a_27 n1398 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06810 n1398 p_11_2_d2j n1594 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06809 n1594 p_11_2_d2jbar n1399 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06808 n1399 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06807 vss p_11_29_t_s p_11_29_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06806 p_11_29_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06805 n1594 n1593 p_11_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06804 p_11_29_t_s n1594 n1593 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06803 n1998 p_11_2_d2j n1996 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06802 n1997 p_11_2_d2jbar n1998 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06801 p_11_28_t_s n1998 n1994 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06800 n1998 n1994 p_11_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06799 p_11_28_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06798 vss p_11_28_t_s p_11_28_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06797 n1994 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06796 vss a_27 n1997 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06795 n1996 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06794 vss c_11_28_s1_s n1817 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06793 c_12_26_a c_11_28_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06792 c_11_28_s1_s p_11_28_pi2j c_11_28_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06791 c_11_28_s2_s n1817 c_10_29_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06790 n1817 c_10_29_cout c_11_28_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06789 vss p_11_28_pi2j n1988 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06788 n1988 c_11_28_a n1987 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06787 n1987 c_10_29_cout n1986 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06786 vss p_11_28_pi2j n1986 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06785 n1986 c_11_28_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06784 vss n1987 c_12_27_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06783 p_11_28_pi2j c_11_28_a c_11_28_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06782 vss n2395 c_11_27_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06781 n2176 c_11_27_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06780 vss c_11_27_a n2176 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06779 n2395 c_11_27_cin n2176 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06778 n1985 c_11_27_b n2395 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06777 vss c_11_27_a n1985 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06776 n2392 c_11_27_cin c_11_27_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06775 c_11_27_s2_s n2392 c_11_27_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06774 c_11_27_a c_11_27_b c_11_27_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06773 c_11_27_s1_s c_11_27_a c_11_27_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06772 c_12_25_a c_11_27_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06771 vss c_11_27_s1_s n2392 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06770 n2403 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06769 vss a_25 n2182 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06768 n2182 p_11_2_d2j n2402 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06767 n2402 p_11_2_d2jbar n2181 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06766 n2181 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06765 vss p_11_27_t_s c_11_27_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06764 c_11_27_b p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06763 n2402 n2403 p_11_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06762 p_11_27_t_s n2402 n2403 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06761 n2642 p_11_2_d2j n2643 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06760 n2641 p_11_2_d2jbar n2642 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06759 p_11_26_t_s n2642 n2640 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06758 n2642 n2640 p_11_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06757 p_11_26_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06756 vss p_11_26_t_s p_11_26_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06755 n2640 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06754 vss a_25 n2641 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06753 n2643 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06752 vss c_11_26_s1_s n2639 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06751 c_12_24_a c_11_26_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06750 c_11_26_s1_s p_11_26_pi2j c_11_26_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06749 c_11_26_s2_s n2639 c_10_27_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06748 n2639 c_10_27_cout c_11_26_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06747 vss p_11_26_pi2j n2809 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06746 n2809 c_11_26_a n2808 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06745 n2808 c_10_27_cout n2810 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06744 vss p_11_26_pi2j n2810 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06743 n2810 c_11_26_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06742 vss n2808 c_12_25_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06741 p_11_26_pi2j c_11_26_a c_11_26_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06740 vss n3199 c_11_25_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06739 n2807 c_11_25_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06738 vss c_11_25_a n2807 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06737 n3199 c_11_25_cin n2807 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06736 n2806 c_11_25_b n3199 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06735 vss c_11_25_a n2806 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06734 n2995 c_11_25_cin c_11_25_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06733 c_11_25_s2_s n2995 c_11_25_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06732 c_11_25_a c_11_25_b c_11_25_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06731 c_11_25_s1_s c_11_25_a c_11_25_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06730 c_12_23_a c_11_25_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06729 vss c_11_25_s1_s n2995 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06728 n3207 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06727 vss a_23 n2816 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06726 n2816 p_11_2_d2j n2998 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06725 n2998 p_11_2_d2jbar n2817 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06724 n2817 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06723 vss p_11_25_t_s c_11_25_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06722 c_11_25_b p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06721 n2998 n3207 p_11_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06720 p_11_25_t_s n2998 n3207 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06719 n3428 p_11_2_d2j n3429 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06718 n3427 p_11_2_d2jbar n3428 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06717 p_11_24_t_s n3428 n3426 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06716 n3428 n3426 p_11_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06715 c_11_24_b p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06714 vss p_11_24_t_s c_11_24_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06713 n3426 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06712 vss a_23 n3427 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06711 n3429 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06710 vss c_11_24_s1_s n3425 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06709 c_12_22_a c_11_24_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06708 c_11_24_s1_s c_11_24_b c_11_24_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06707 c_11_24_s2_s n3425 c_10_25_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06706 n3425 c_10_25_cout c_11_24_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06705 vss c_11_24_b n3586 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06704 n3586 c_11_24_a n3419 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06703 n3419 c_10_25_cout n3587 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06702 vss c_11_24_b n3587 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06701 n3587 c_11_24_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06700 vss n3419 c_12_23_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06699 c_11_24_b c_11_24_a c_11_24_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06698 vss n3789 c_11_23_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06697 n3585 c_11_23_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06696 vss c_11_23_a n3585 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06695 n3789 c_11_23_cin n3585 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06694 n3584 c_11_23_b n3789 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06693 vss c_11_23_a n3584 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06692 n3796 c_11_23_cin c_11_23_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06691 c_11_23_s2_s n3796 c_11_23_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06690 c_11_23_a c_11_23_b c_11_23_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06689 c_11_23_s1_s c_11_23_a c_11_23_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06688 c_12_21_a c_11_23_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06687 vss c_11_23_s1_s n3796 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06686 n3799 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06685 vss a_21 n3590 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06684 n3590 p_11_2_d2j n3801 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06683 n3801 p_11_2_d2jbar n3591 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06682 n3591 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06681 vss p_11_23_t_s c_11_23_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06680 c_11_23_b p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06679 n3801 n3799 p_11_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06678 p_11_23_t_s n3801 n3799 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06677 n4224 p_11_2_d2j n4225 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06676 n4223 p_11_2_d2jbar n4224 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06675 p_11_22_t_s n4224 n4221 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06674 n4224 n4221 p_11_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06673 p_11_22_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06672 vss p_11_22_t_s p_11_22_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06671 n4221 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06670 vss a_21 n4223 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06669 n4225 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06668 vss c_11_22_s1_s n4219 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06667 c_12_20_a c_11_22_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06666 c_11_22_s1_s p_11_22_pi2j c_11_22_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06665 c_11_22_s2_s n4219 c_10_23_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06664 n4219 c_10_23_cout c_11_22_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06663 vss p_11_22_pi2j n4213 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06662 n4213 c_11_22_a n4212 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06661 n4212 c_10_23_cout n4214 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06660 vss p_11_22_pi2j n4214 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06659 n4214 c_11_22_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06658 vss n4212 c_12_21_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06657 p_11_22_pi2j c_11_22_a c_11_22_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06656 vss n4558 c_11_21_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06655 n4381 p_11_21_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06654 vss c_11_21_a n4381 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06653 n4558 c_11_21_cin n4381 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06652 n4380 p_11_21_pi2j n4558 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06651 vss c_11_21_a n4380 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06650 n4563 c_11_21_cin c_11_21_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06649 c_11_21_s2_s n4563 c_11_21_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06648 c_11_21_a p_11_21_pi2j c_11_21_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06647 c_11_21_s1_s c_11_21_a p_11_21_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06646 c_12_19_a c_11_21_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06645 vss c_11_21_s1_s n4563 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06644 n4568 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06643 vss a_19 n4382 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06642 n4382 p_11_2_d2j n4570 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06641 n4570 p_11_2_d2jbar n4383 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06640 n4383 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06639 vss p_11_21_t_s p_11_21_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06638 p_11_21_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06637 n4570 n4568 p_11_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06636 p_11_21_t_s n4570 n4568 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06635 n4970 p_11_2_d2j n4971 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06634 n4969 p_11_2_d2jbar n4970 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06633 p_11_20_t_s n4970 n4967 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06632 n4970 n4967 p_11_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06631 p_11_20_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06630 vss p_11_20_t_s p_11_20_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06629 n4967 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06628 vss a_19 n4969 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06627 n4971 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06626 vss c_11_20_s1_s n4963 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06625 c_12_18_a c_11_20_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06624 c_11_20_s1_s p_11_20_pi2j c_11_20_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06623 c_11_20_s2_s n4963 c_10_21_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06622 n4963 c_10_21_cout c_11_20_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06621 vss p_11_20_pi2j n4959 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06620 n4959 c_11_20_a n4960 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06619 n4960 c_10_21_cout n4958 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06618 vss p_11_20_pi2j n4958 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06617 n4958 c_11_20_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06616 vss n4960 c_12_19_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06615 p_11_20_pi2j c_11_20_a c_11_20_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06614 vss n5309 c_11_19_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06613 n5122 p_11_19_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06612 vss c_11_19_a n5122 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06611 n5309 c_11_19_cin n5122 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06610 n5121 p_11_19_pi2j n5309 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06609 vss c_11_19_a n5121 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06608 n5315 c_11_19_cin c_11_19_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06607 c_11_19_s2_s n5315 c_11_19_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06606 c_11_19_a p_11_19_pi2j c_11_19_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06605 c_11_19_s1_s c_11_19_a p_11_19_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06604 c_12_17_a c_11_19_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06603 vss c_11_19_s1_s n5315 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06602 n5320 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06601 vss a_17 n5123 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06600 n5123 p_11_2_d2j n5321 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06599 n5321 p_11_2_d2jbar n5124 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06598 n5124 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06597 vss p_11_19_t_s p_11_19_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06596 p_11_19_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06595 n5321 n5320 p_11_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06594 p_11_19_t_s n5321 n5320 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06593 n5723 p_11_2_d2j n5724 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06592 n5722 p_11_2_d2jbar n5723 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06591 p_11_18_t_s n5723 n5720 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06590 n5723 n5720 p_11_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06589 p_11_18_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06588 vss p_11_18_t_s p_11_18_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06587 n5720 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06586 vss a_17 n5722 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06585 n5724 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06584 vss c_11_18_s1_s n5543 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06583 c_12_16_a c_11_18_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06582 c_11_18_s1_s p_11_18_pi2j c_11_18_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06581 c_11_18_s2_s n5543 c_10_19_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06580 n5543 c_10_19_cout c_11_18_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06579 vss p_11_18_pi2j n5712 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06578 n5712 c_11_18_a n5714 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06577 n5714 c_10_19_cout n5713 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06576 vss p_11_18_pi2j n5713 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06575 n5713 c_11_18_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06574 vss n5714 c_12_17_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06573 p_11_18_pi2j c_11_18_a c_11_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06572 vss n6095 c_11_17_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06571 n5887 p_11_17_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06570 vss c_11_17_a n5887 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06569 n6095 c_11_17_cin n5887 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06568 n5711 p_11_17_pi2j n6095 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06567 vss c_11_17_a n5711 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06566 n6090 c_11_17_cin c_11_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06565 c_11_17_s2_s n6090 c_11_17_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06564 c_11_17_a p_11_17_pi2j c_11_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06563 c_11_17_s1_s c_11_17_a p_11_17_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06562 c_12_15_a c_11_17_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06561 vss c_11_17_s1_s n6090 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06560 n6104 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06559 vss a_15 n5890 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06558 n5890 p_11_2_d2j n6103 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06557 n6103 p_11_2_d2jbar n5891 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06556 n5891 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06555 vss p_11_17_t_s p_11_17_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06554 p_11_17_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06553 n6103 n6104 p_11_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06552 p_11_17_t_s n6103 n6104 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06551 n6346 p_11_2_d2j n6347 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06550 n6345 p_11_2_d2jbar n6346 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06549 p_11_16_t_s n6346 n6507 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06548 n6346 n6507 p_11_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06547 p_11_16_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06546 vss p_11_16_t_s p_11_16_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06545 n6507 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06544 vss a_15 n6345 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06543 n6347 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06542 vss c_11_16_s1_s n6344 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06541 c_12_14_a c_11_16_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06540 c_11_16_s1_s p_11_16_pi2j c_11_16_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06539 c_11_16_s2_s n6344 c_10_17_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06538 n6344 c_10_17_cout c_11_16_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06537 vss p_11_16_pi2j n6500 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06536 n6500 c_11_16_a n6501 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06535 n6501 c_10_17_cout n6499 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06534 vss p_11_16_pi2j n6499 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06533 n6499 c_11_16_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06532 vss n6501 c_12_15_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06531 p_11_16_pi2j c_11_16_a c_11_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06530 vss n6902 c_11_15_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06529 n6498 c_11_15_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06528 vss c_11_15_a n6498 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06527 n6902 c_11_15_cin n6498 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06526 n6497 c_11_15_b n6902 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06525 vss c_11_15_a n6497 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06524 n6696 c_11_15_cin c_11_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06523 c_11_15_s2_s n6696 c_11_15_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06522 c_11_15_a c_11_15_b c_11_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06521 c_11_15_s1_s c_11_15_a c_11_15_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06520 c_12_13_a c_11_15_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06519 vss c_11_15_s1_s n6696 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06518 n6909 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06517 vss a_13 n6508 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06516 n6508 p_11_2_d2j n6699 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06515 n6699 p_11_2_d2jbar n6509 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06514 n6509 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06513 vss p_11_15_t_s c_11_15_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06512 c_11_15_b p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06511 n6699 n6909 p_11_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06510 p_11_15_t_s n6699 n6909 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06509 n7129 p_11_2_d2j n7130 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06508 n7128 p_11_2_d2jbar n7129 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06507 p_11_14_t_s n7129 n7127 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06506 n7129 n7127 p_11_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06505 p_11_14_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06504 vss p_11_14_t_s p_11_14_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06503 n7127 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06502 vss a_13 n7128 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06501 n7130 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06500 vss c_11_14_s1_s n7126 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06499 c_12_12_a c_11_14_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06498 c_11_14_s1_s p_11_14_pi2j c_11_14_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06497 c_11_14_s2_s n7126 c_10_15_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06496 n7126 c_10_15_cout c_11_14_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06495 vss p_11_14_pi2j n7288 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06494 n7288 c_11_14_a n7121 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06493 n7121 c_10_15_cout n7289 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06492 vss p_11_14_pi2j n7289 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06491 n7289 c_11_14_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06490 vss n7121 c_12_13_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06489 p_11_14_pi2j c_11_14_a c_11_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06488 vss n7473 c_11_13_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06487 n7287 c_11_13_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06486 vss c_11_13_a n7287 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06485 n7473 c_11_13_cin n7287 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06484 n7286 c_11_13_b n7473 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06483 vss c_11_13_a n7286 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06482 n7480 c_11_13_cin c_11_13_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06481 c_11_13_s2_s n7480 c_11_13_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06480 c_11_13_a c_11_13_b c_11_13_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06479 c_11_13_s1_s c_11_13_a c_11_13_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06478 c_12_11_a c_11_13_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06477 vss c_11_13_s1_s n7480 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06476 n7482 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06475 vss a_11 n7293 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06474 n7293 p_11_2_d2j n7484 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06473 n7484 p_11_2_d2jbar n7294 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06472 n7294 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06471 vss p_11_13_t_s c_11_13_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06470 c_11_13_b p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06469 n7484 n7482 p_11_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06468 p_11_13_t_s n7484 n7482 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06467 n7911 p_11_2_d2j n7912 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06466 n7910 p_11_2_d2jbar n7911 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06465 p_11_12_t_s n7911 n7908 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06464 n7911 n7908 p_11_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06463 c_11_12_b p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06462 vss p_11_12_t_s c_11_12_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06461 n7908 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06460 vss a_11 n7910 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06459 n7912 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06458 vss c_11_12_s1_s n7907 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06457 c_12_10_a c_11_12_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06456 c_11_12_s1_s c_11_12_b c_11_12_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06455 c_11_12_s2_s n7907 c_10_13_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06454 n7907 c_10_13_cout c_11_12_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06453 vss c_11_12_b n7901 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06452 n7901 c_11_12_a n7902 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06451 n7902 c_10_13_cout n7900 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06450 vss c_11_12_b n7900 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06449 n7900 c_11_12_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06448 vss n7902 c_12_11_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06447 c_11_12_b c_11_12_a c_11_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06446 vss n8247 c_11_11_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06445 n8063 p_11_11_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06444 vss c_11_11_a n8063 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06443 n8247 c_11_11_cin n8063 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06442 n8062 p_11_11_pi2j n8247 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06441 vss c_11_11_a n8062 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06440 n8251 c_11_11_cin c_11_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06439 c_11_11_s2_s n8251 c_11_11_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06438 c_11_11_a p_11_11_pi2j c_11_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06437 c_11_11_s1_s c_11_11_a p_11_11_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06436 c_12_9_a c_11_11_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06435 vss c_11_11_s1_s n8251 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06434 n8256 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06433 vss a_9 n8065 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06432 n8065 p_11_2_d2j n8258 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06431 n8258 p_11_2_d2jbar n8066 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06430 n8066 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06429 vss p_11_11_t_s p_11_11_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06428 p_11_11_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06427 n8258 n8256 p_11_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06426 p_11_11_t_s n8258 n8256 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06425 n8659 p_11_2_d2j n8660 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06424 n8658 p_11_2_d2jbar n8659 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06423 p_11_10_t_s n8659 n8657 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06422 n8659 n8657 p_11_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06421 p_11_10_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06420 vss p_11_10_t_s p_11_10_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06419 n8657 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06418 vss a_9 n8658 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06417 n8660 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06416 vss c_11_10_s1_s n8653 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06415 c_12_8_a c_11_10_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06414 c_11_10_s1_s p_11_10_pi2j c_11_10_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06413 c_11_10_s2_s n8653 c_10_11_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06412 n8653 c_10_11_cout c_11_10_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06411 vss p_11_10_pi2j n8649 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06410 n8649 c_11_10_a n8647 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06409 n8647 c_10_11_cout n8648 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06408 vss p_11_10_pi2j n8648 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06407 n8648 c_11_10_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06406 vss n8647 c_12_9_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06405 p_11_10_pi2j c_11_10_a c_11_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06404 vss n8997 c_11_9_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06403 n8814 p_11_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06402 vss c_11_9_a n8814 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06401 n8997 c_11_9_cin n8814 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06400 n8813 p_11_9_pi2j n8997 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06399 vss c_11_9_a n8813 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06398 n9003 c_11_9_cin c_11_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06397 c_11_9_s2_s n9003 c_11_9_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06396 c_11_9_a p_11_9_pi2j c_11_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06395 c_11_9_s1_s c_11_9_a p_11_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06394 c_12_7_a c_11_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06393 vss c_11_9_s1_s n9003 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06392 n9008 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06391 vss a_7 n8815 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06390 n8815 p_11_2_d2j n9010 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06389 n9010 p_11_2_d2jbar n8816 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06388 n8816 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06387 vss p_11_9_t_s p_11_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06386 p_11_9_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06385 n9010 n9008 p_11_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06384 p_11_9_t_s n9010 n9008 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06383 n9397 p_11_2_d2j n9398 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06382 n9396 p_11_2_d2jbar n9397 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06381 p_11_8_t_s n9397 n9394 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06380 n9397 n9394 p_11_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06379 p_11_8_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06378 vss p_11_8_t_s p_11_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06377 n9394 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06376 vss a_7 n9396 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06375 n9398 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06374 vss c_11_8_s1_s n9389 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06373 c_12_6_a c_11_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06372 c_11_8_s1_s p_11_8_pi2j c_11_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06371 c_11_8_s2_s n9389 c_10_9_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06370 n9389 c_10_9_cout c_11_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06369 vss p_11_8_pi2j n9385 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06368 n9385 c_11_8_a n9386 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06367 n9386 c_10_9_cout n9387 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06366 vss p_11_8_pi2j n9387 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06365 n9387 c_11_8_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06364 vss n9386 c_12_7_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06363 p_11_8_pi2j c_11_8_a c_11_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06362 vss n9777 c_11_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06361 n9565 p_11_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06360 vss c_11_7_a n9565 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06359 n9777 c_11_7_cin n9565 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06358 n9384 p_11_7_pi2j n9777 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06357 vss c_11_7_a n9384 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06356 n9785 c_11_7_cin c_11_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06355 c_11_7_s2_s n9785 c_11_7_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06354 c_11_7_a p_11_7_pi2j c_11_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06353 c_11_7_s1_s c_11_7_a p_11_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06352 c_12_5_a c_11_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06351 vss c_11_7_s1_s n9785 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06350 n9788 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06349 vss a_5 n9568 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06348 n9568 p_11_2_d2j n9787 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06347 n9787 p_11_2_d2jbar n9569 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06346 n9569 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06345 vss p_11_7_t_s p_11_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06344 p_11_7_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06343 n9787 n9788 p_11_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06342 p_11_7_t_s n9787 n9788 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06341 n10174 p_11_2_d2j n10019 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06340 n10018 p_11_2_d2jbar n10174 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06339 p_11_6_t_s n10174 n10175 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06338 n10174 n10175 p_11_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06337 c_11_6_b p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06336 vss p_11_6_t_s c_11_6_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06335 n10175 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06334 vss a_5 n10018 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06333 n10019 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06332 vss c_11_6_s1_s n10017 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06331 c_12_4_a c_11_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06330 c_11_6_s1_s c_11_6_b c_11_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06329 c_11_6_s2_s n10017 c_10_7_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06328 n10017 c_10_7_cout c_11_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06327 vss c_11_6_b n10166 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06326 n10166 c_11_6_a n10167 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06325 n10167 c_10_7_cout n10165 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06324 vss c_11_6_b n10165 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06323 n10165 c_11_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06322 vss n10167 c_12_5_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06321 c_11_6_b c_11_6_a c_11_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06320 vss n10574 c_11_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06319 n10366 c_11_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06318 vss c_11_5_a n10366 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06317 n10574 c_11_5_cin n10366 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06316 n10164 c_11_5_b n10574 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06315 vss c_11_5_a n10164 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06314 n10371 c_11_5_cin c_11_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06313 c_11_5_s2_s n10371 c_11_5_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06312 c_11_5_a c_11_5_b c_11_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06311 c_11_5_s1_s c_11_5_a c_11_5_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06310 c_12_3_a c_11_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06309 vss c_11_5_s1_s n10371 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06308 n10583 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06307 vss a_3 n10176 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06306 n10176 p_11_2_d2j n10581 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06305 n10581 p_11_2_d2jbar n10177 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06304 n10177 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06303 vss p_11_5_t_s c_11_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06302 c_11_5_b p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06301 n10581 n10583 p_11_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06300 p_11_5_t_s n10581 n10583 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06299 n10803 p_11_2_d2j n10804 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06298 n10802 p_11_2_d2jbar n10803 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06297 p_11_4_t_s n10803 n10801 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06296 n10803 n10801 p_11_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06295 p_11_4_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06294 vss p_11_4_t_s p_11_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06293 n10801 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06292 vss a_3 n10802 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06291 n10804 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06290 vss c_11_4_s1_s n10800 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06289 c_12_2_a c_11_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06288 c_11_4_s1_s p_11_4_pi2j c_11_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06287 c_11_4_s2_s n10800 c_10_5_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06286 n10800 c_10_5_cout c_11_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06285 vss p_11_4_pi2j n10956 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06284 n10956 c_11_4_a n10795 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06283 n10795 c_10_5_cout n10957 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06282 vss p_11_4_pi2j n10957 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06281 n10957 c_11_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06280 vss n10795 c_12_3_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06279 p_11_4_pi2j c_11_4_a c_11_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06278 vss n11138 c_11_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06277 n10955 c_11_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06276 vss c_11_3_a n10955 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06275 n11138 c_11_3_cin n10955 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06274 n10954 c_11_3_b n11138 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06273 vss c_11_3_a n10954 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06272 n11144 c_11_3_cin c_11_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06271 c_11_3_s2_s n11144 c_11_3_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06270 c_11_3_a c_11_3_b c_11_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06269 c_11_3_s1_s c_11_3_a c_11_3_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06268 c_12_1_a c_11_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06267 vss c_11_3_s1_s n11144 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06266 n11147 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06265 vss a_1 n10961 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06264 n10961 p_11_2_d2j n11149 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06263 n11149 p_11_2_d2jbar n10962 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06262 n10962 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06261 vss p_11_3_t_s c_11_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06260 c_11_3_b p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06259 n11149 n11147 p_11_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06258 p_11_3_t_s n11149 n11147 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06257 n11574 p_11_2_d2j n11575 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06256 n11573 p_11_2_d2jbar n11574 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06255 p_11_2_t_s n11574 n11571 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06254 n11574 n11571 p_11_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06253 c_11_2_b p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06252 vss p_11_2_t_s c_11_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06251 n11571 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06250 vss a_1 n11573 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06249 n11575 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06248 vss c_11_2_s1_s n11570 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06247 c_11_2_sum c_11_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06246 c_11_2_s1_s c_11_2_b c_11_2_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06245 c_11_2_s2_s n11570 c_10_3_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06244 n11570 c_10_3_cout c_11_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06243 vss c_11_2_b n11564 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06242 n11564 c_11_2_a n11565 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06241 n11565 c_10_3_cout n11563 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06240 vss c_11_2_b n11563 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06239 n11563 c_11_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06238 vss n11565 c_12_1_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06237 c_11_2_b c_11_2_a c_11_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06236 vss n11907 c_11_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06235 n11725 p_11_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06234 vss c_11_1_a n11725 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06233 n11907 c_11_1_cin n11725 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06232 n11724 p_11_1_pi2j n11907 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06231 vss c_11_1_a n11724 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06230 n11915 c_11_1_cin c_11_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06229 c_11_1_s2_s n11915 c_11_1_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06228 c_11_1_a p_11_1_pi2j c_11_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06227 c_11_1_s1_s c_11_1_a p_11_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06226 c_11_1_sum c_11_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06225 vss c_11_1_s1_s n11915 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06224 n11917 p_11_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06223 n11921 p_11_2_d2jbar n11728 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06222 n11728 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06221 vss p_11_1_t_s p_11_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06220 p_11_1_pi2j p_11_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06219 n11921 n11917 p_11_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06218 p_11_1_t_s n11921 n11917 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06217 cl4_11_s1_s n12287 c_10_1_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06216 n12287 c_10_1_sum cl4_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06215 vss cl4_11_s1_s p_16 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06214 vss c_10_1_sum n12277 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06213 n12277 n12287 n12278 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06212 n12279 n12278 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_06211 n12276 c_10_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_06210 vss c_10_2_sum n12276 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_06209 n12273 c_10_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06208 n12274 c_10_1_cout n12273 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06207 n12271 c_10_1_sum n12274 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06206 n12276 n12287 n12271 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06205 n12272 n12274 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_06204 cl4_11_s2_s c_10_1_cout c_10_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06203 c_10_1_cout c_10_2_sum cl4_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06202 vss cl4_11_s2_s n12270 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06201 cl4_11_s3_s n12270 n12279 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06200 n12270 n12279 cl4_11_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06199 vss cl4_11_s3_s p_17 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_06198 vss c_10_33_s1_s n149 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06197 c_11_31_a c_10_33_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06196 c_10_33_s1_s c_10_31_a p_10_33_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06195 c_10_31_a p_10_33_pi2j c_10_33_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06194 c_10_33_s2_s n149 c_10_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06193 n149 c_10_32_cin c_10_33_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06192 vss c_10_31_a n19 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_06191 n19 p_10_33_pi2j n148 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06190 n148 c_10_32_cin n20 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06189 vss c_10_31_a n20 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_06188 n20 p_10_33_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06187 vss n148 c_11_32_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06186 n156 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06185 n159 a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06184 vss p_10_33_t_s p_10_33_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06183 p_10_33_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06182 n159 n156 p_10_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06181 p_10_33_t_s n159 n156 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06180 n503 p_10_2_d2j n501 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06179 n502 p_10_2_d2jbar n503 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06178 p_10_32_t_s n503 n499 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06177 n503 n499 p_10_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06176 p_10_32_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06175 vss p_10_32_t_s p_10_32_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06174 n499 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06173 vss a_31 n502 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06172 n501 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06171 vss c_10_32_s1_s n496 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06170 c_11_30_a c_10_32_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06169 c_10_32_s1_s p_10_32_pi2j c_10_31_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06168 c_10_32_s2_s n496 c_10_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06167 n496 c_10_32_cin c_10_32_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06166 vss p_10_32_pi2j n492 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06165 n492 c_10_31_a n491 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06164 n491 c_10_32_cin n493 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06163 vss p_10_32_pi2j n493 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06162 n493 c_10_31_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06161 vss n491 c_11_31_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06160 p_10_32_pi2j c_10_31_a c_10_32_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06159 vss n833 c_10_31_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06158 n634 p_10_31_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06157 vss c_10_31_a n634 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06156 n833 c_10_31_cin n634 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06155 n633 p_10_31_pi2j n833 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06154 vss c_10_31_a n633 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06153 n829 c_10_31_cin c_10_31_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06152 c_10_31_s2_s n829 c_10_31_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06151 c_10_31_a p_10_31_pi2j c_10_31_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06150 c_10_31_s1_s c_10_31_a p_10_31_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06149 c_11_29_a c_10_31_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06148 vss c_10_31_s1_s n829 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06147 n839 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06146 vss a_29 n635 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06145 n635 p_10_2_d2j n841 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06144 n841 p_10_2_d2jbar n636 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06143 n636 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06142 vss p_10_31_t_s p_10_31_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06141 p_10_31_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06140 n841 n839 p_10_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06139 p_10_31_t_s n841 n839 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06138 n1255 p_10_2_d2j n1256 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06137 n1254 p_10_2_d2jbar n1255 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06136 p_10_30_t_s n1255 n1253 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06135 n1255 n1253 p_10_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06134 p_10_30_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06133 vss p_10_30_t_s p_10_30_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06132 n1253 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06131 vss a_29 n1254 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06130 n1256 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06129 vss c_10_30_s1_s n1249 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06128 c_11_28_a c_10_30_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06127 c_10_30_s1_s p_10_30_pi2j c_10_30_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06126 c_10_30_s2_s n1249 c_9_31_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06125 n1249 c_9_31_cout c_10_30_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06124 vss p_10_30_pi2j n1245 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06123 n1245 c_10_30_a n1243 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06122 n1243 c_9_31_cout n1244 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06121 vss p_10_30_pi2j n1244 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06120 n1244 c_10_30_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06119 vss n1243 c_11_29_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06118 p_10_30_pi2j c_10_30_a c_10_30_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06117 vss n1606 c_10_29_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06116 n1400 p_10_29_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06115 vss c_10_29_a n1400 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06114 n1606 c_10_29_cin n1400 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06113 n1242 p_10_29_pi2j n1606 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06112 vss c_10_29_a n1242 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06111 n1601 c_10_29_cin c_10_29_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06110 c_10_29_s2_s n1601 c_10_29_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06109 c_10_29_a p_10_29_pi2j c_10_29_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06108 c_10_29_s1_s c_10_29_a p_10_29_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06107 c_11_27_a c_10_29_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06106 vss c_10_29_s1_s n1601 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06105 n1613 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06104 vss a_27 n1401 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06103 n1401 p_10_2_d2j n1615 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06102 n1615 p_10_2_d2jbar n1402 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06101 n1402 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06100 vss p_10_29_t_s p_10_29_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06099 p_10_29_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06098 n1615 n1613 p_10_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06097 p_10_29_t_s n1615 n1613 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06096 n2011 p_10_2_d2j n2012 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06095 n2010 p_10_2_d2jbar n2011 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06094 p_10_28_t_s n2011 n2009 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06093 n2011 n2009 p_10_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06092 p_10_28_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06091 vss p_10_28_t_s p_10_28_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06090 n2009 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06089 vss a_27 n2010 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06088 n2012 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06087 vss c_10_28_s1_s n1823 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06086 c_11_26_a c_10_28_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06085 c_10_28_s1_s p_10_28_pi2j c_10_28_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06084 c_10_28_s2_s n1823 c_9_29_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06083 n1823 c_9_29_cout c_10_28_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06082 vss p_10_28_pi2j n2001 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06081 n2001 c_10_28_a n2000 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06080 n2000 c_9_29_cout n2002 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06079 vss p_10_28_pi2j n2002 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06078 n2002 c_10_28_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06077 vss n2000 c_11_27_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06076 p_10_28_pi2j c_10_28_a c_10_28_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06075 vss n2418 c_10_27_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06074 n2183 c_10_27_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06073 vss c_10_27_a n2183 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06072 n2418 c_10_27_cin n2183 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06071 n1999 c_10_27_b n2418 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06070 vss c_10_27_a n1999 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06069 n2410 c_10_27_cin c_10_27_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06068 c_10_27_s2_s n2410 c_10_27_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06067 c_10_27_a c_10_27_b c_10_27_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06066 c_10_27_s1_s c_10_27_a c_10_27_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06065 c_11_25_a c_10_27_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06064 vss c_10_27_s1_s n2410 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06063 n2423 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06062 vss a_25 n2188 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06061 n2188 p_10_2_d2j n2419 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06060 n2419 p_10_2_d2jbar n2189 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06059 n2189 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06058 vss p_10_27_t_s c_10_27_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06057 c_10_27_b p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06056 n2419 n2423 p_10_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06055 p_10_27_t_s n2419 n2423 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06054 n2650 p_10_2_d2j n2649 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06053 n2651 p_10_2_d2jbar n2650 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06052 p_10_26_t_s n2650 n2648 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06051 n2650 n2648 p_10_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06050 p_10_26_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06049 vss p_10_26_t_s p_10_26_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06048 n2648 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06047 vss a_25 n2651 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06046 n2649 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06045 vss c_10_26_s1_s n2647 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06044 c_11_24_a c_10_26_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06043 c_10_26_s1_s p_10_26_pi2j c_10_26_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06042 c_10_26_s2_s n2647 c_9_27_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06041 n2647 c_9_27_cout c_10_26_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06040 vss p_10_26_pi2j n2821 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06039 n2821 c_10_26_a n2820 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06038 n2820 c_9_27_cout n2822 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06037 vss p_10_26_pi2j n2822 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06036 n2822 c_10_26_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06035 vss n2820 c_11_25_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06034 p_10_26_pi2j c_10_26_a c_10_26_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06033 vss n3218 c_10_25_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_06032 n2819 c_10_25_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06031 vss c_10_25_a n2819 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06030 n3218 c_10_25_cin n2819 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06029 n2818 c_10_25_b n3218 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06028 vss c_10_25_a n2818 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_06027 n3001 c_10_25_cin c_10_25_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06026 c_10_25_s2_s n3001 c_10_25_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06025 c_10_25_a c_10_25_b c_10_25_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06024 c_10_25_s1_s c_10_25_a c_10_25_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06023 c_11_23_a c_10_25_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06022 vss c_10_25_s1_s n3001 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06021 n3224 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06020 vss a_23 n2829 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06019 n2829 p_10_2_d2j n3007 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06018 n3007 p_10_2_d2jbar n2828 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06017 n2828 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06016 vss p_10_25_t_s c_10_25_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06015 c_10_25_b p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06014 n3007 n3224 p_10_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06013 p_10_25_t_s n3007 n3224 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06012 n3439 p_10_2_d2j n3440 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06011 n3438 p_10_2_d2jbar n3439 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_06010 p_10_24_t_s n3439 n3437 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06009 n3439 n3437 p_10_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06008 c_10_24_b p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06007 vss p_10_24_t_s c_10_24_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_06006 n3437 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_06005 vss a_23 n3438 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06004 n3440 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_06003 vss c_10_24_s1_s n3434 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_06002 c_11_22_a c_10_24_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_06001 c_10_24_s1_s c_10_24_b c_10_24_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_06000 c_10_24_s2_s n3434 c_9_25_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05999 n3434 c_9_25_cout c_10_24_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05998 vss c_10_24_b n3595 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05997 n3595 c_10_24_a n3430 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05996 n3430 c_9_25_cout n3594 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05995 vss c_10_24_b n3594 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05994 n3594 c_10_24_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05993 vss n3430 c_11_23_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05992 c_10_24_b c_10_24_a c_10_24_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05991 vss n3807 c_10_23_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05990 n3593 c_10_23_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05989 vss c_10_23_a n3593 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05988 n3807 c_10_23_cin n3593 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05987 n3592 c_10_23_b n3807 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05986 vss c_10_23_a n3592 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05985 n3810 c_10_23_cin c_10_23_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05984 c_10_23_s2_s n3810 c_10_23_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05983 c_10_23_a c_10_23_b c_10_23_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05982 c_10_23_s1_s c_10_23_a c_10_23_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05981 c_11_21_a c_10_23_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05980 vss c_10_23_s1_s n3810 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05979 n3815 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05978 vss a_21 n3598 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05977 n3598 p_10_2_d2j n3817 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05976 n3817 p_10_2_d2jbar n3599 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05975 n3599 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05974 vss p_10_23_t_s c_10_23_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05973 c_10_23_b p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05972 n3817 n3815 p_10_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05971 p_10_23_t_s n3817 n3815 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05970 n4239 p_10_2_d2j n4237 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05969 n4238 p_10_2_d2jbar n4239 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05968 p_10_22_t_s n4239 n4236 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05967 n4239 n4236 p_10_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05966 p_10_22_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05965 vss p_10_22_t_s p_10_22_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05964 n4236 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05963 vss a_21 n4238 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05962 n4237 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05961 vss c_10_22_s1_s n4231 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05960 c_11_20_a c_10_22_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05959 c_10_22_s1_s p_10_22_pi2j c_10_22_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05958 c_10_22_s2_s n4231 c_9_23_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05957 n4231 c_9_23_cout c_10_22_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05956 vss p_10_22_pi2j n4227 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05955 n4227 c_10_22_a n4226 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05954 n4226 c_9_23_cout n4228 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05953 vss p_10_22_pi2j n4228 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05952 n4228 c_10_22_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05951 vss n4226 c_11_21_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05950 p_10_22_pi2j c_10_22_a c_10_22_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05949 vss n4578 c_10_21_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05948 n4385 p_10_21_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05947 vss c_10_21_a n4385 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05946 n4578 c_10_21_cin n4385 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05945 n4384 p_10_21_pi2j n4578 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05944 vss c_10_21_a n4384 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05943 n4574 c_10_21_cin c_10_21_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05942 c_10_21_s2_s n4574 c_10_21_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05941 c_10_21_a p_10_21_pi2j c_10_21_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05940 c_10_21_s1_s c_10_21_a p_10_21_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05939 c_11_19_a c_10_21_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05938 vss c_10_21_s1_s n4574 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05937 n4586 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05936 vss a_19 n4386 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05935 n4386 p_10_2_d2j n4588 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05934 n4588 p_10_2_d2jbar n4387 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05933 n4387 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05932 vss p_10_21_t_s p_10_21_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05931 p_10_21_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05930 n4588 n4586 p_10_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05929 p_10_21_t_s n4588 n4586 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05928 n4985 p_10_2_d2j n4984 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05927 n4983 p_10_2_d2jbar n4985 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05926 p_10_20_t_s n4985 n4982 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05925 n4985 n4982 p_10_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05924 p_10_20_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05923 vss p_10_20_t_s p_10_20_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05922 n4982 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05921 vss a_19 n4983 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05920 n4984 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05919 vss c_10_20_s1_s n4978 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05918 c_11_18_a c_10_20_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05917 c_10_20_s1_s p_10_20_pi2j c_10_20_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05916 c_10_20_s2_s n4978 c_9_21_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05915 n4978 c_9_21_cout c_10_20_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05914 vss p_10_20_pi2j n4973 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05913 n4973 c_10_20_a n4974 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05912 n4974 c_9_21_cout n4972 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05911 vss p_10_20_pi2j n4972 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05910 n4972 c_10_20_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05909 vss n4974 c_11_19_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05908 p_10_20_pi2j c_10_20_a c_10_20_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05907 vss n5332 c_10_19_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05906 n5126 p_10_19_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05905 vss c_10_19_a n5126 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05904 n5332 c_10_19_cin n5126 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05903 n5125 p_10_19_pi2j n5332 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05902 vss c_10_19_a n5125 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05901 n5328 c_10_19_cin c_10_19_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05900 c_10_19_s2_s n5328 c_10_19_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05899 c_10_19_a p_10_19_pi2j c_10_19_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05898 c_10_19_s1_s c_10_19_a p_10_19_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05897 c_11_17_a c_10_19_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05896 vss c_10_19_s1_s n5328 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05895 n5340 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05894 vss a_17 n5127 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05893 n5127 p_10_2_d2j n5342 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05892 n5342 p_10_2_d2jbar n5128 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05891 n5128 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05890 vss p_10_19_t_s p_10_19_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05889 p_10_19_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05888 n5342 n5340 p_10_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05887 p_10_19_t_s n5342 n5340 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05886 n5737 p_10_2_d2j n5736 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05885 n5738 p_10_2_d2jbar n5737 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05884 p_10_18_t_s n5737 n5735 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05883 n5737 n5735 p_10_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05882 p_10_18_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05881 vss p_10_18_t_s p_10_18_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05880 n5735 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05879 vss a_17 n5738 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05878 n5736 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05877 vss c_10_18_s1_s n5549 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05876 c_11_16_a c_10_18_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05875 c_10_18_s1_s p_10_18_pi2j c_10_18_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05874 c_10_18_s2_s n5549 c_9_19_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05873 n5549 c_9_19_cout c_10_18_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05872 vss p_10_18_pi2j n5726 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05871 n5726 c_10_18_a n5728 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05870 n5728 c_9_19_cout n5727 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05869 vss p_10_18_pi2j n5727 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05868 n5727 c_10_18_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05867 vss n5728 c_11_17_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05866 p_10_18_pi2j c_10_18_a c_10_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05865 vss n6119 c_10_17_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05864 n5892 p_10_17_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05863 vss c_10_17_a n5892 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05862 n6119 c_10_17_cin n5892 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05861 n5725 p_10_17_pi2j n6119 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05860 vss c_10_17_a n5725 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05859 n6112 c_10_17_cin c_10_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05858 c_10_17_s2_s n6112 c_10_17_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05857 c_10_17_a p_10_17_pi2j c_10_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05856 c_10_17_s1_s c_10_17_a p_10_17_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05855 c_11_15_a c_10_17_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05854 vss c_10_17_s1_s n6112 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05853 n6126 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05852 vss a_15 n5896 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05851 n5896 p_10_2_d2j n6121 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05850 n6121 p_10_2_d2jbar n5895 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05849 n5895 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05848 vss p_10_17_t_s p_10_17_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05847 p_10_17_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05846 n6121 n6126 p_10_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05845 p_10_17_t_s n6121 n6126 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05844 n6354 p_10_2_d2j n6353 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05843 n6352 p_10_2_d2jbar n6354 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05842 p_10_16_t_s n6354 n6520 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05841 n6354 n6520 p_10_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05840 p_10_16_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05839 vss p_10_16_t_s p_10_16_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05838 n6520 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05837 vss a_15 n6352 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05836 n6353 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05835 vss c_10_16_s1_s n6351 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05834 c_11_14_a c_10_16_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05833 c_10_16_s1_s p_10_16_pi2j c_10_16_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05832 c_10_16_s2_s n6351 c_9_17_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05831 n6351 c_9_17_cout c_10_16_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05830 vss p_10_16_pi2j n6512 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05829 n6512 c_10_16_a n6513 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05828 n6513 c_9_17_cout n6514 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05827 vss p_10_16_pi2j n6514 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05826 n6514 c_10_16_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05825 vss n6513 c_11_15_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05824 p_10_16_pi2j c_10_16_a c_10_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05823 vss n6921 c_10_15_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05822 n6511 c_10_15_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05821 vss c_10_15_a n6511 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05820 n6921 c_10_15_cin n6511 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05819 n6510 c_10_15_b n6921 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05818 vss c_10_15_a n6510 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05817 n6702 c_10_15_cin c_10_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05816 c_10_15_s2_s n6702 c_10_15_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05815 c_10_15_a c_10_15_b c_10_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05814 c_10_15_s1_s c_10_15_a c_10_15_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05813 c_11_13_a c_10_15_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05812 vss c_10_15_s1_s n6702 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05811 n6926 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05810 vss a_13 n6521 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05809 n6521 p_10_2_d2j n6708 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05808 n6708 p_10_2_d2jbar n6522 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05807 n6522 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05806 vss p_10_15_t_s c_10_15_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05805 c_10_15_b p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05804 n6708 n6926 p_10_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05803 p_10_15_t_s n6708 n6926 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05802 n7139 p_10_2_d2j n7140 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05801 n7138 p_10_2_d2jbar n7139 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05800 p_10_14_t_s n7139 n7137 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05799 n7139 n7137 p_10_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05798 p_10_14_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05797 vss p_10_14_t_s p_10_14_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05796 n7137 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05795 vss a_13 n7138 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05794 n7140 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05793 vss c_10_14_s1_s n7134 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05792 c_11_12_a c_10_14_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05791 c_10_14_s1_s p_10_14_pi2j c_10_14_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05790 c_10_14_s2_s n7134 c_9_15_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05789 n7134 c_9_15_cout c_10_14_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05788 vss p_10_14_pi2j n7297 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05787 n7297 c_10_14_a n7131 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05786 n7131 c_9_15_cout n7298 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05785 vss p_10_14_pi2j n7298 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05784 n7298 c_10_14_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05783 vss n7131 c_11_13_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05782 p_10_14_pi2j c_10_14_a c_10_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05781 vss n7487 c_10_13_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05780 n7296 c_10_13_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05779 vss c_10_13_a n7296 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05778 n7487 c_10_13_cin n7296 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05777 n7295 c_10_13_b n7487 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05776 vss c_10_13_a n7295 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05775 n7491 c_10_13_cin c_10_13_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05774 c_10_13_s2_s n7491 c_10_13_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05773 c_10_13_a c_10_13_b c_10_13_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05772 c_10_13_s1_s c_10_13_a c_10_13_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05771 c_11_11_a c_10_13_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05770 vss c_10_13_s1_s n7491 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05769 n7495 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05768 vss a_11 n7303 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05767 n7303 p_10_2_d2j n7497 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05766 n7497 p_10_2_d2jbar n7302 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05765 n7302 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05764 vss p_10_13_t_s c_10_13_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05763 c_10_13_b p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05762 n7497 n7495 p_10_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05761 p_10_13_t_s n7497 n7495 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05760 n7925 p_10_2_d2j n7923 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05759 n7924 p_10_2_d2jbar n7925 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05758 p_10_12_t_s n7925 n7922 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05757 n7925 n7922 p_10_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05756 c_10_12_b p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05755 vss p_10_12_t_s c_10_12_b vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05754 n7922 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05753 vss a_11 n7924 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05752 n7923 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05751 vss c_10_12_s1_s n7918 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05750 c_11_10_a c_10_12_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05749 c_10_12_s1_s c_10_12_b c_10_12_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05748 c_10_12_s2_s n7918 c_9_13_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05747 n7918 c_9_13_cout c_10_12_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05746 vss c_10_12_b n7914 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05745 n7914 c_10_12_a n7915 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05744 n7915 c_9_13_cout n7913 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05743 vss c_10_12_b n7913 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05742 n7913 c_10_12_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05741 vss n7915 c_11_11_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05740 c_10_12_b c_10_12_a c_10_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05739 vss n8267 c_10_11_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05738 n8068 p_10_11_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05737 vss c_10_11_a n8068 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05736 n8267 c_10_11_cin n8068 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05735 n8067 p_10_11_pi2j n8267 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05734 vss c_10_11_a n8067 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05733 n8262 c_10_11_cin c_10_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05732 c_10_11_s2_s n8262 c_10_11_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05731 c_10_11_a p_10_11_pi2j c_10_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05730 c_10_11_s1_s c_10_11_a p_10_11_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05729 c_11_9_a c_10_11_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05728 vss c_10_11_s1_s n8262 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05727 n8274 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05726 vss a_9 n8070 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05725 n8070 p_10_2_d2j n8276 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05724 n8276 p_10_2_d2jbar n8071 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05723 n8071 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05722 vss p_10_11_t_s p_10_11_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05721 p_10_11_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05720 n8276 n8274 p_10_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05719 p_10_11_t_s n8276 n8274 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05718 n8673 p_10_2_d2j n8674 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05717 n8672 p_10_2_d2jbar n8673 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05716 p_10_10_t_s n8673 n8671 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05715 n8673 n8671 p_10_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05714 p_10_10_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05713 vss p_10_10_t_s p_10_10_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05712 n8671 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05711 vss a_9 n8672 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05710 n8674 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05709 vss c_10_10_s1_s n8667 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05708 c_11_8_a c_10_10_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05707 c_10_10_s1_s p_10_10_pi2j c_10_10_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05706 c_10_10_s2_s n8667 c_9_11_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05705 n8667 c_9_11_cout c_10_10_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05704 vss p_10_10_pi2j n8663 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05703 n8663 c_10_10_a n8661 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05702 n8661 c_9_11_cout n8662 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05701 vss p_10_10_pi2j n8662 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05700 n8662 c_10_10_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05699 vss n8661 c_11_9_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05698 p_10_10_pi2j c_10_10_a c_10_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05697 vss n9020 c_10_9_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05696 n8818 p_10_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05695 vss c_10_9_a n8818 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05694 n9020 c_10_9_cin n8818 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05693 n8817 p_10_9_pi2j n9020 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05692 vss c_10_9_a n8817 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05691 n9016 c_10_9_cin c_10_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05690 c_10_9_s2_s n9016 c_10_9_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05689 c_10_9_a p_10_9_pi2j c_10_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05688 c_10_9_s1_s c_10_9_a p_10_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05687 c_11_7_a c_10_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05686 vss c_10_9_s1_s n9016 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05685 n9028 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05684 vss a_7 n8819 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05683 n8819 p_10_2_d2j n9030 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05682 n9030 p_10_2_d2jbar n8820 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05681 n8820 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05680 vss p_10_9_t_s p_10_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05679 p_10_9_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05678 n9030 n9028 p_10_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05677 p_10_9_t_s n9030 n9028 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05676 n9413 p_10_2_d2j n9411 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05675 n9412 p_10_2_d2jbar n9413 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05674 p_10_8_t_s n9413 n9410 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05673 n9413 n9410 p_10_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05672 p_10_8_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05671 vss p_10_8_t_s p_10_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05670 n9410 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05669 vss a_7 n9412 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05668 n9411 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05667 vss c_10_8_s1_s n9405 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05666 c_11_6_a c_10_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05665 c_10_8_s1_s p_10_8_pi2j c_10_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05664 c_10_8_s2_s n9405 c_9_9_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05663 n9405 c_9_9_cout c_10_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05662 vss p_10_8_pi2j n9400 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05661 n9400 c_10_8_a n9402 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05660 n9402 c_9_9_cout n9401 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05659 vss p_10_8_pi2j n9401 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05658 n9401 c_10_8_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05657 vss n9402 c_11_7_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05656 p_10_8_pi2j c_10_8_a c_10_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05655 vss n9803 c_10_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05654 n9570 p_10_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05653 vss c_10_7_a n9570 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05652 n9803 c_10_7_cin n9570 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05651 n9399 p_10_7_pi2j n9803 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05650 vss c_10_7_a n9399 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05649 n9798 c_10_7_cin c_10_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05648 c_10_7_s2_s n9798 c_10_7_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05647 c_10_7_a p_10_7_pi2j c_10_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05646 c_10_7_s1_s c_10_7_a p_10_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05645 c_11_5_a c_10_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05644 vss c_10_7_s1_s n9798 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05643 n9810 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05642 vss a_5 n9573 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05641 n9573 p_10_2_d2j n9805 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05640 n9805 p_10_2_d2jbar n9574 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05639 n9574 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05638 vss p_10_7_t_s p_10_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05637 p_10_7_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05636 n9805 n9810 p_10_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05635 p_10_7_t_s n9805 n9810 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05634 n10188 p_10_2_d2j n10024 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05633 n10023 p_10_2_d2jbar n10188 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05632 p_10_6_t_s n10188 n10189 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05631 n10188 n10189 p_10_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05630 p_10_6_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05629 vss p_10_6_t_s p_10_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05628 n10189 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05627 vss a_5 n10023 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05626 n10024 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05625 vss c_10_6_s1_s n10022 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05624 c_11_4_a c_10_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05623 c_10_6_s1_s p_10_6_pi2j c_10_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05622 c_10_6_s2_s n10022 c_9_7_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05621 n10022 c_9_7_cout c_10_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05620 vss p_10_6_pi2j n10180 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05619 n10180 c_10_6_a n10181 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05618 n10181 c_9_7_cout n10182 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05617 vss p_10_6_pi2j n10182 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05616 n10182 c_10_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05615 vss n10181 c_11_5_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05614 p_10_6_pi2j c_10_6_a c_10_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05613 vss n10592 c_10_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05612 n10375 c_10_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05611 vss c_10_5_a n10375 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05610 n10592 c_10_5_cin n10375 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05609 n10179 c_10_5_b n10592 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05608 vss c_10_5_a n10179 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05607 n10377 c_10_5_cin c_10_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05606 c_10_5_s2_s n10377 c_10_5_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05605 c_10_5_a c_10_5_b c_10_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05604 c_10_5_s1_s c_10_5_a c_10_5_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05603 c_11_3_a c_10_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05602 vss c_10_5_s1_s n10377 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05601 n10600 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05600 vss a_3 n10190 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05599 n10190 p_10_2_d2j n10595 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05598 n10595 p_10_2_d2jbar n10191 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05597 n10191 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05596 vss p_10_5_t_s c_10_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05595 c_10_5_b p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05594 n10595 n10600 p_10_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05593 p_10_5_t_s n10595 n10600 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05592 n10814 p_10_2_d2j n10812 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05591 n10813 p_10_2_d2jbar n10814 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05590 p_10_4_t_s n10814 n10811 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05589 n10814 n10811 p_10_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05588 p_10_4_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05587 vss p_10_4_t_s p_10_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05586 n10811 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05585 vss a_3 n10813 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05584 n10812 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05583 vss c_10_4_s1_s n10809 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05582 c_11_2_a c_10_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05581 c_10_4_s1_s p_10_4_pi2j c_10_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05580 c_10_4_s2_s n10809 c_9_5_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05579 n10809 c_9_5_cout c_10_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05578 vss p_10_4_pi2j n10965 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05577 n10965 c_10_4_a n10805 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05576 n10805 c_9_5_cout n10966 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05575 vss p_10_4_pi2j n10966 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05574 n10966 c_10_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05573 vss n10805 c_11_3_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05572 p_10_4_pi2j c_10_4_a c_10_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05571 vss n11152 c_10_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05570 n10964 c_10_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05569 vss c_10_3_a n10964 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05568 n11152 c_10_3_cin n10964 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05567 n10963 c_10_3_b n11152 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05566 vss c_10_3_a n10963 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05565 n11155 c_10_3_cin c_10_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05564 c_10_3_s2_s n11155 c_10_3_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05563 c_10_3_a c_10_3_b c_10_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05562 c_10_3_s1_s c_10_3_a c_10_3_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05561 c_11_1_a c_10_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05560 vss c_10_3_s1_s n11155 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05559 n11160 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05558 vss a_1 n10971 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05557 n10971 p_10_2_d2j n11162 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05556 n11162 p_10_2_d2jbar n10970 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05555 n10970 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05554 vss p_10_3_t_s c_10_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05553 c_10_3_b p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05552 n11162 n11160 p_10_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05551 p_10_3_t_s n11162 n11160 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05550 n11587 p_10_2_d2j n11588 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05549 n11586 p_10_2_d2jbar n11587 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05548 p_10_2_t_s n11587 n11585 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05547 n11587 n11585 p_10_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05546 c_10_2_b p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05545 vss p_10_2_t_s c_10_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05544 n11585 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05543 vss a_1 n11586 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05542 n11588 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05541 vss c_10_2_s1_s n11581 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05540 c_10_2_sum c_10_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05539 c_10_2_s1_s c_10_2_b c_10_2_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05538 c_10_2_s2_s n11581 c_9_3_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05537 n11581 c_9_3_cout c_10_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05536 vss c_10_2_b n11577 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05535 n11577 c_10_2_a n11578 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05534 n11578 c_9_3_cout n11576 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05533 vss c_10_2_b n11576 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05532 n11576 c_10_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05531 vss n11578 c_11_1_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05530 c_10_2_b c_10_2_a c_10_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05529 vss n11928 c_10_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05528 n11730 p_10_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05527 vss c_10_1_a n11730 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05526 n11928 c_10_1_cin n11730 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05525 n11729 p_10_1_pi2j n11928 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05524 vss c_10_1_a n11729 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05523 n11924 c_10_1_cin c_10_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05522 c_10_1_s2_s n11924 c_10_1_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05521 c_10_1_a p_10_1_pi2j c_10_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05520 c_10_1_s1_s c_10_1_a p_10_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05519 c_10_1_sum c_10_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05518 vss c_10_1_s1_s n11924 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05517 n11938 p_10_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05516 n11940 p_10_2_d2jbar n11733 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05515 n11733 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05514 vss p_10_1_t_s p_10_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05513 p_10_1_pi2j p_10_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05512 n11940 n11938 p_10_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05511 p_10_1_t_s n11940 n11938 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05510 cl4_10_s1_s n12305 c_9_1_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05509 n12305 c_9_1_sum cl4_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05508 vss cl4_10_s1_s p_14 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05507 vss c_9_1_sum n12295 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05506 n12295 n12305 n12296 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05505 n12293 n12296 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_05504 n12294 c_9_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_05503 vss c_9_2_sum n12294 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_05502 n12291 c_9_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05501 n12290 c_9_1_cout n12291 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05500 n12289 c_9_1_sum n12290 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05499 n12294 n12305 n12289 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05498 n12287 n12290 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_05497 cl4_10_s2_s c_9_1_cout c_9_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05496 c_9_1_cout c_9_2_sum cl4_10_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05495 vss cl4_10_s2_s n12286 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05494 cl4_10_s3_s n12286 n12293 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05493 n12286 n12293 cl4_10_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05492 vss cl4_10_s3_s p_15 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05491 vss c_9_33_s1_s n163 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05490 c_10_31_a c_9_33_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05489 c_9_33_s1_s c_9_31_a p_9_33_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05488 c_9_31_a p_9_33_pi2j c_9_33_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05487 c_9_33_s2_s n163 c_9_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05486 n163 c_9_32_cin c_9_33_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05485 vss c_9_31_a n22 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_05484 n22 p_9_33_pi2j n162 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05483 n162 c_9_32_cin n21 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05482 vss c_9_31_a n21 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_05481 n21 p_9_33_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05480 vss n162 c_10_32_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05479 n172 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05478 n173 a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05477 vss p_9_33_t_s p_9_33_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05476 p_9_33_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05475 n173 n172 p_9_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05474 p_9_33_t_s n173 n172 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05473 n515 p_9_2_d2j n516 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05472 n514 p_9_2_d2jbar n515 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05471 p_9_32_t_s n515 n513 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05470 n515 n513 p_9_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05469 p_9_32_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05468 vss p_9_32_t_s p_9_32_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05467 n513 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05466 vss a_31 n514 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05465 n516 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05464 vss c_9_32_s1_s n510 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05463 c_10_30_a c_9_32_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05462 c_9_32_s1_s p_9_32_pi2j c_9_31_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05461 c_9_32_s2_s n510 c_9_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05460 n510 c_9_32_cin c_9_32_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05459 vss p_9_32_pi2j n504 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05458 n504 c_9_31_a n505 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05457 n505 c_9_32_cin n506 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05456 vss p_9_32_pi2j n506 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05455 n506 c_9_31_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_05454 vss n505 c_10_31_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05453 p_9_32_pi2j c_9_31_a c_9_32_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05452 vss n852 c_9_31_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05451 n638 p_9_31_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05450 vss c_9_31_a n638 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_05449 n852 c_9_31_cin n638 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05448 n637 p_9_31_pi2j n852 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05447 vss c_9_31_a n637 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_05446 n848 c_9_31_cin c_9_31_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05445 c_9_31_s2_s n848 c_9_31_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05444 c_9_31_a p_9_31_pi2j c_9_31_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05443 c_9_31_s1_s c_9_31_a p_9_31_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05442 c_10_29_a c_9_31_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05441 vss c_9_31_s1_s n848 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05440 n858 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05439 vss a_29 n639 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05438 n639 p_9_2_d2j n857 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05437 n857 p_9_2_d2jbar n640 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05436 n640 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05435 vss p_9_31_t_s p_9_31_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05434 p_9_31_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05433 n857 n858 p_9_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05432 p_9_31_t_s n857 n858 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05431 n1270 p_9_2_d2j n1271 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05430 n1269 p_9_2_d2jbar n1270 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05429 p_9_30_t_s n1270 n1268 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05428 n1270 n1268 p_9_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05427 p_9_30_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05426 vss p_9_30_t_s p_9_30_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05425 n1268 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05424 vss a_29 n1269 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05423 n1271 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05422 vss c_9_30_s1_s n1263 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05421 c_10_28_a c_9_30_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05420 c_9_30_s1_s p_9_30_pi2j c_9_30_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05419 c_9_30_s2_s n1263 c_8_31_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05418 n1263 c_8_31_cout c_9_30_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05417 vss p_9_30_pi2j n1259 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05416 n1259 c_9_30_a n1260 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05415 n1260 c_8_31_cout n1258 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05414 vss p_9_30_pi2j n1258 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05413 n1258 c_9_30_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05412 vss n1260 c_10_29_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05411 p_9_30_pi2j c_9_30_a c_9_30_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05410 vss n1627 c_9_29_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05409 n1403 p_9_29_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05408 vss c_9_29_a n1403 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05407 n1627 c_9_29_cin n1403 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05406 n1257 p_9_29_pi2j n1627 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05405 vss c_9_29_a n1257 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05404 n1624 c_9_29_cin c_9_29_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05403 c_9_29_s2_s n1624 c_9_29_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05402 c_9_29_a p_9_29_pi2j c_9_29_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05401 c_9_29_s1_s c_9_29_a p_9_29_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05400 c_10_27_a c_9_29_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05399 vss c_9_29_s1_s n1624 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05398 n1635 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05397 vss a_27 n1404 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05396 n1404 p_9_2_d2j n1633 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05395 n1633 p_9_2_d2jbar n1405 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05394 n1405 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05393 vss p_9_29_t_s p_9_29_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05392 p_9_29_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05391 n1633 n1635 p_9_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05390 p_9_29_t_s n1633 n1635 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05389 n2025 p_9_2_d2j n2026 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05388 n2024 p_9_2_d2jbar n2025 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05387 p_9_28_t_s n2025 n2023 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05386 n2025 n2023 p_9_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05385 p_9_28_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05384 vss p_9_28_t_s p_9_28_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05383 n2023 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05382 vss a_27 n2024 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05381 n2026 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05380 vss c_9_28_s1_s n1830 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05379 c_10_26_a c_9_28_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05378 c_9_28_s1_s p_9_28_pi2j c_9_28_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05377 c_9_28_s2_s n1830 c_8_29_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05376 n1830 c_8_29_cout c_9_28_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05375 vss p_9_28_pi2j n2016 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05374 n2016 c_9_28_a n2015 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05373 n2015 c_8_29_cout n2014 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05372 vss p_9_28_pi2j n2014 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05371 n2014 c_9_28_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05370 vss n2015 c_10_27_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05369 p_9_28_pi2j c_9_28_a c_9_28_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05368 vss n2438 c_9_27_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05367 n2190 c_9_27_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05366 vss c_9_27_a n2190 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05365 n2438 c_9_27_cin n2190 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05364 n2013 c_9_27_b n2438 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05363 vss c_9_27_a n2013 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05362 n2431 c_9_27_cin c_9_27_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05361 c_9_27_s2_s n2431 c_9_27_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05360 c_9_27_a c_9_27_b c_9_27_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05359 c_9_27_s1_s c_9_27_a c_9_27_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05358 c_10_25_a c_9_27_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05357 vss c_9_27_s1_s n2431 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05356 n2445 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05355 vss a_25 n2194 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05354 n2194 p_9_2_d2j n2441 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05353 n2441 p_9_2_d2jbar n2196 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05352 n2196 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05351 vss p_9_27_t_s c_9_27_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05350 c_9_27_b p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05349 n2441 n2445 p_9_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05348 p_9_27_t_s n2441 n2445 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05347 n2657 p_9_2_d2j n2659 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05346 n2658 p_9_2_d2jbar n2657 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05345 p_9_26_t_s n2657 n2656 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05344 n2657 n2656 p_9_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05343 p_9_26_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05342 vss p_9_26_t_s p_9_26_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05341 n2656 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05340 vss a_25 n2658 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05339 n2659 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05338 vss c_9_26_s1_s n2655 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05337 c_10_24_a c_9_26_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05336 c_9_26_s1_s p_9_26_pi2j c_9_26_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05335 c_9_26_s2_s n2655 c_8_27_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05334 n2655 c_8_27_cout c_9_26_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05333 vss p_9_26_pi2j n2833 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05332 n2833 c_9_26_a n2832 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05331 n2832 c_8_27_cout n2834 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05330 vss p_9_26_pi2j n2834 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05329 n2834 c_9_26_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05328 vss n2832 c_10_25_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05327 p_9_26_pi2j c_9_26_a c_9_26_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05326 vss n3236 c_9_25_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05325 n2831 c_9_25_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05324 vss c_9_25_a n2831 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05323 n3236 c_9_25_cin n2831 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05322 n2830 c_9_25_b n3236 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05321 vss c_9_25_a n2830 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05320 n3012 c_9_25_cin c_9_25_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05319 c_9_25_s2_s n3012 c_9_25_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05318 c_9_25_a c_9_25_b c_9_25_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05317 c_9_25_s1_s c_9_25_a c_9_25_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05316 c_10_23_a c_9_25_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05315 vss c_9_25_s1_s n3012 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05314 n3240 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05313 vss a_23 n2840 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05312 n2840 p_9_2_d2j n3015 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05311 n3015 p_9_2_d2jbar n2841 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05310 n2841 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05309 vss p_9_25_t_s c_9_25_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05308 c_9_25_b p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05307 n3015 n3240 p_9_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05306 p_9_25_t_s n3015 n3240 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05305 n3449 p_9_2_d2j n3451 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05304 n3450 p_9_2_d2jbar n3449 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05303 p_9_24_t_s n3449 n3448 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05302 n3449 n3448 p_9_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05301 c_9_24_b p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05300 vss p_9_24_t_s c_9_24_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05299 n3448 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05298 vss a_23 n3450 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05297 n3451 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05296 vss c_9_24_s1_s n3447 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05295 c_10_22_a c_9_24_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05294 c_9_24_s1_s c_9_24_b c_9_24_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05293 c_9_24_s2_s n3447 c_8_25_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05292 n3447 c_8_25_cout c_9_24_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05291 vss c_9_24_b n3602 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05290 n3602 c_9_24_a n3441 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05289 n3441 c_8_25_cout n3603 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05288 vss c_9_24_b n3603 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05287 n3603 c_9_24_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05286 vss n3441 c_10_23_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05285 c_9_24_b c_9_24_a c_9_24_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05284 vss n3825 c_9_23_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05283 n3601 c_9_23_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05282 vss c_9_23_a n3601 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05281 n3825 c_9_23_cin n3601 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05280 n3600 c_9_23_b n3825 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05279 vss c_9_23_a n3600 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05278 n3827 c_9_23_cin c_9_23_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05277 c_9_23_s2_s n3827 c_9_23_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05276 c_9_23_a c_9_23_b c_9_23_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05275 c_9_23_s1_s c_9_23_a c_9_23_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05274 c_10_21_a c_9_23_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05273 vss c_9_23_s1_s n3827 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05272 n3832 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05271 vss a_21 n3606 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05270 n3606 p_9_2_d2j n3831 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05269 n3831 p_9_2_d2jbar n3608 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05268 n3608 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05267 vss p_9_23_t_s c_9_23_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05266 c_9_23_b p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05265 n3831 n3832 p_9_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05264 p_9_23_t_s n3831 n3832 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05263 n4251 p_9_2_d2j n4253 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05262 n4252 p_9_2_d2jbar n4251 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05261 p_9_22_t_s n4251 n4249 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05260 n4251 n4249 p_9_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05259 p_9_22_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05258 vss p_9_22_t_s p_9_22_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05257 n4249 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05256 vss a_21 n4252 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05255 n4253 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05254 vss c_9_22_s1_s n4247 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05253 c_10_20_a c_9_22_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05252 c_9_22_s1_s p_9_22_pi2j c_9_22_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05251 c_9_22_s2_s n4247 c_8_23_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05250 n4247 c_8_23_cout c_9_22_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05249 vss p_9_22_pi2j n4240 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05248 n4240 c_9_22_a n4241 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05247 n4241 c_8_23_cout n4242 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05246 vss p_9_22_pi2j n4242 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05245 n4242 c_9_22_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05244 vss n4241 c_10_21_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05243 p_9_22_pi2j c_9_22_a c_9_22_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05242 vss n4596 c_9_21_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05241 n4389 p_9_21_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05240 vss c_9_21_a n4389 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05239 n4596 c_9_21_cin n4389 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05238 n4388 p_9_21_pi2j n4596 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05237 vss c_9_21_a n4388 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05236 n4593 c_9_21_cin c_9_21_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05235 c_9_21_s2_s n4593 c_9_21_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05234 c_9_21_a p_9_21_pi2j c_9_21_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05233 c_9_21_s1_s c_9_21_a p_9_21_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05232 c_10_19_a c_9_21_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05231 vss c_9_21_s1_s n4593 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05230 n4605 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05229 vss a_19 n4390 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05228 n4390 p_9_2_d2j n4604 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05227 n4604 p_9_2_d2jbar n4391 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05226 n4391 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05225 vss p_9_21_t_s p_9_21_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05224 p_9_21_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05223 n4604 n4605 p_9_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05222 p_9_21_t_s n4604 n4605 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05221 n4997 p_9_2_d2j n4999 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05220 n4998 p_9_2_d2jbar n4997 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05219 p_9_20_t_s n4997 n4995 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05218 n4997 n4995 p_9_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05217 p_9_20_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05216 vss p_9_20_t_s p_9_20_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05215 n4995 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05214 vss a_19 n4998 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05213 n4999 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05212 vss c_9_20_s1_s n4993 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05211 c_10_18_a c_9_20_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05210 c_9_20_s1_s p_9_20_pi2j c_9_20_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05209 c_9_20_s2_s n4993 c_8_21_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05208 n4993 c_8_21_cout c_9_20_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05207 vss p_9_20_pi2j n4988 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05206 n4988 c_9_20_a n4987 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05205 n4987 c_8_21_cout n4986 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05204 vss p_9_20_pi2j n4986 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05203 n4986 c_9_20_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05202 vss n4987 c_10_19_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05201 p_9_20_pi2j c_9_20_a c_9_20_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05200 vss n5355 c_9_19_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05199 n5130 p_9_19_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05198 vss c_9_19_a n5130 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05197 n5355 c_9_19_cin n5130 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05196 n5129 p_9_19_pi2j n5355 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05195 vss c_9_19_a n5129 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05194 n5351 c_9_19_cin c_9_19_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05193 c_9_19_s2_s n5351 c_9_19_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05192 c_9_19_a p_9_19_pi2j c_9_19_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05191 c_9_19_s1_s c_9_19_a p_9_19_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05190 c_10_17_a c_9_19_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05189 vss c_9_19_s1_s n5351 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05188 n5362 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05187 vss a_17 n5131 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05186 n5131 p_9_2_d2j n5360 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05185 n5360 p_9_2_d2jbar n5132 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05184 n5132 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05183 vss p_9_19_t_s p_9_19_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05182 p_9_19_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05181 n5360 n5362 p_9_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05180 p_9_19_t_s n5360 n5362 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05179 n5749 p_9_2_d2j n5752 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05178 n5748 p_9_2_d2jbar n5749 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05177 p_9_18_t_s n5749 n5750 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05176 n5749 n5750 p_9_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05175 p_9_18_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05174 vss p_9_18_t_s p_9_18_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05173 n5750 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05172 vss a_17 n5748 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05171 n5752 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05170 vss c_9_18_s1_s n5556 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05169 c_10_16_a c_9_18_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05168 c_9_18_s1_s p_9_18_pi2j c_9_18_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05167 c_9_18_s2_s n5556 c_8_19_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05166 n5556 c_8_19_cout c_9_18_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05165 vss p_9_18_pi2j n5741 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05164 n5741 c_9_18_a n5740 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05163 n5740 c_8_19_cout n5742 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05162 vss p_9_18_pi2j n5742 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05161 n5742 c_9_18_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05160 vss n5740 c_10_17_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05159 p_9_18_pi2j c_9_18_a c_9_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05158 vss n6143 c_9_17_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05157 n5897 p_9_17_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05156 vss c_9_17_a n5897 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05155 n6143 c_9_17_cin n5897 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05154 n5739 p_9_17_pi2j n6143 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05153 vss c_9_17_a n5739 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05152 n6133 c_9_17_cin c_9_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05151 c_9_17_s2_s n6133 c_9_17_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05150 c_9_17_a p_9_17_pi2j c_9_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05149 c_9_17_s1_s c_9_17_a p_9_17_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05148 c_10_15_a c_9_17_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05147 vss c_9_17_s1_s n6133 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05146 n6150 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05145 vss a_15 n5899 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05144 n5899 p_9_2_d2j n6144 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05143 n6144 p_9_2_d2jbar n5901 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05142 n5901 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05141 vss p_9_17_t_s p_9_17_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05140 p_9_17_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05139 n6144 n6150 p_9_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05138 p_9_17_t_s n6144 n6150 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05137 n6359 p_9_2_d2j n6361 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05136 n6360 p_9_2_d2jbar n6359 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05135 p_9_16_t_s n6359 n6533 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05134 n6359 n6533 p_9_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05133 p_9_16_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05132 vss p_9_16_t_s p_9_16_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05131 n6533 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05130 vss a_15 n6360 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05129 n6361 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05128 vss c_9_16_s1_s n6358 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05127 c_10_14_a c_9_16_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05126 c_9_16_s1_s p_9_16_pi2j c_9_16_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05125 c_9_16_s2_s n6358 c_8_17_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05124 n6358 c_8_17_cout c_9_16_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05123 vss p_9_16_pi2j n6525 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05122 n6525 c_9_16_a n6526 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05121 n6526 c_8_17_cout n6527 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05120 vss p_9_16_pi2j n6527 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05119 n6527 c_9_16_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05118 vss n6526 c_10_15_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05117 p_9_16_pi2j c_9_16_a c_9_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05116 vss n6939 c_9_15_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05115 n6524 c_9_15_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05114 vss c_9_15_a n6524 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05113 n6939 c_9_15_cin n6524 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05112 n6523 c_9_15_b n6939 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05111 vss c_9_15_a n6523 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05110 n6713 c_9_15_cin c_9_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05109 c_9_15_s2_s n6713 c_9_15_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05108 c_9_15_a c_9_15_b c_9_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05107 c_9_15_s1_s c_9_15_a c_9_15_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05106 c_10_13_a c_9_15_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05105 vss c_9_15_s1_s n6713 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05104 n6942 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05103 vss a_13 n6534 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05102 n6534 p_9_2_d2j n6716 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05101 n6716 p_9_2_d2jbar n6535 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05100 n6535 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05099 vss p_9_15_t_s c_9_15_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05098 c_9_15_b p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05097 n6716 n6942 p_9_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05096 p_9_15_t_s n6716 n6942 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05095 n7148 p_9_2_d2j n7150 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05094 n7149 p_9_2_d2jbar n7148 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05093 p_9_14_t_s n7148 n7147 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05092 n7148 n7147 p_9_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05091 p_9_14_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05090 vss p_9_14_t_s p_9_14_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05089 n7147 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05088 vss a_13 n7149 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05087 n7150 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05086 vss c_9_14_s1_s n7146 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05085 c_10_12_a c_9_14_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05084 c_9_14_s1_s p_9_14_pi2j c_9_14_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05083 c_9_14_s2_s n7146 c_8_15_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05082 n7146 c_8_15_cout c_9_14_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05081 vss p_9_14_pi2j n7306 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05080 n7306 c_9_14_a n7141 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05079 n7141 c_8_15_cout n7307 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05078 vss p_9_14_pi2j n7307 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05077 n7307 c_9_14_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05076 vss n7141 c_10_13_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05075 p_9_14_pi2j c_9_14_a c_9_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05074 vss n7503 c_9_13_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05073 n7305 c_9_13_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05072 vss c_9_13_a n7305 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05071 n7503 c_9_13_cin n7305 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05070 n7304 c_9_13_b n7503 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05069 vss c_9_13_a n7304 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05068 n7505 c_9_13_cin c_9_13_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05067 c_9_13_s2_s n7505 c_9_13_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05066 c_9_13_a c_9_13_b c_9_13_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05065 c_9_13_s1_s c_9_13_a c_9_13_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05064 c_10_11_a c_9_13_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05063 vss c_9_13_s1_s n7505 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05062 n7509 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05061 vss a_11 n7311 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05060 n7311 p_9_2_d2j n7508 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05059 n7508 p_9_2_d2jbar n7312 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05058 n7312 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05057 vss p_9_13_t_s c_9_13_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05056 c_9_13_b p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05055 n7508 n7509 p_9_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05054 p_9_13_t_s n7508 n7509 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05053 n7936 p_9_2_d2j n7938 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05052 n7937 p_9_2_d2jbar n7936 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05051 p_9_12_t_s n7936 n7934 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05050 n7936 n7934 p_9_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05049 c_9_12_b p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05048 vss p_9_12_t_s c_9_12_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_05047 n7934 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05046 vss a_11 n7937 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05045 n7938 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05044 vss c_9_12_s1_s n7933 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05043 c_10_10_a c_9_12_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05042 c_9_12_s1_s c_9_12_b c_9_12_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05041 c_9_12_s2_s n7933 c_8_13_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05040 n7933 c_8_13_cout c_9_12_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05039 vss c_9_12_b n7926 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05038 n7926 c_9_12_a n7928 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05037 n7928 c_8_13_cout n7927 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05036 vss c_9_12_b n7927 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05035 n7927 c_9_12_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05034 vss n7928 c_10_11_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05033 c_9_12_b c_9_12_a c_9_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05032 vss n8286 c_9_11_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_05031 n8073 p_9_11_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05030 vss c_9_11_a n8073 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05029 n8286 c_9_11_cin n8073 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05028 n8072 p_9_11_pi2j n8286 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05027 vss c_9_11_a n8072 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_05026 n8281 c_9_11_cin c_9_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05025 c_9_11_s2_s n8281 c_9_11_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05024 c_9_11_a p_9_11_pi2j c_9_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05023 c_9_11_s1_s c_9_11_a p_9_11_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_05022 c_10_9_a c_9_11_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05021 vss c_9_11_s1_s n8281 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05020 n8293 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05019 vss a_9 n8075 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05018 n8075 p_9_2_d2j n8292 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05017 n8292 p_9_2_d2jbar n8076 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05016 n8076 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05015 vss p_9_11_t_s p_9_11_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05014 p_9_11_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05013 n8292 n8293 p_9_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05012 p_9_11_t_s n8292 n8293 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05011 n8686 p_9_2_d2j n8688 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05010 n8687 p_9_2_d2jbar n8686 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_05009 p_9_10_t_s n8686 n8684 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05008 n8686 n8684 p_9_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05007 p_9_10_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05006 vss p_9_10_t_s p_9_10_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_05005 n8684 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_05004 vss a_9 n8687 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05003 n8688 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_05002 vss c_9_10_s1_s n8680 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_05001 c_10_8_a c_9_10_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_05000 c_9_10_s1_s p_9_10_pi2j c_9_10_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04999 c_9_10_s2_s n8680 c_8_11_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04998 n8680 c_8_11_cout c_9_10_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04997 vss p_9_10_pi2j n8677 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04996 n8677 c_9_10_a n8676 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04995 n8676 c_8_11_cout n8675 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04994 vss p_9_10_pi2j n8675 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04993 n8675 c_9_10_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04992 vss n8676 c_10_9_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04991 p_9_10_pi2j c_9_10_a c_9_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04990 vss n9043 c_9_9_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04989 n8822 p_9_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04988 vss c_9_9_a n8822 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04987 n9043 c_9_9_cin n8822 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04986 n8821 p_9_9_pi2j n9043 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04985 vss c_9_9_a n8821 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04984 n9039 c_9_9_cin c_9_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04983 c_9_9_s2_s n9039 c_9_9_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04982 c_9_9_a p_9_9_pi2j c_9_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04981 c_9_9_s1_s c_9_9_a p_9_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04980 c_10_7_a c_9_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04979 vss c_9_9_s1_s n9039 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04978 n9050 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04977 vss a_7 n8823 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04976 n8823 p_9_2_d2j n9048 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04975 n9048 p_9_2_d2jbar n8824 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04974 n8824 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04973 vss p_9_9_t_s p_9_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04972 p_9_9_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04971 n9048 n9050 p_9_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04970 p_9_9_t_s n9048 n9050 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04969 n9425 p_9_2_d2j n9428 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04968 n9424 p_9_2_d2jbar n9425 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04967 p_9_8_t_s n9425 n9426 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04966 n9425 n9426 p_9_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04965 p_9_8_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04964 vss p_9_8_t_s p_9_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04963 n9426 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04962 vss a_7 n9424 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04961 n9428 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04960 vss c_9_8_s1_s n9414 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04959 c_10_6_a c_9_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04958 c_9_8_s1_s p_9_8_pi2j c_9_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04957 c_9_8_s2_s n9414 c_8_9_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04956 n9414 c_8_9_cout c_9_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04955 vss p_9_8_pi2j n9417 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04954 n9417 c_9_8_a n9416 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04953 n9416 c_8_9_cout n9418 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04952 vss p_9_8_pi2j n9418 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04951 n9418 c_9_8_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04950 vss n9416 c_10_7_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04949 p_9_8_pi2j c_9_8_a c_9_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04948 vss n9826 c_9_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04947 n9575 p_9_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04946 vss c_9_7_a n9575 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04945 n9826 c_9_7_cin n9575 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04944 n9415 p_9_7_pi2j n9826 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04943 vss c_9_7_a n9415 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04942 n9821 c_9_7_cin c_9_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04941 c_9_7_s2_s n9821 c_9_7_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04940 c_9_7_a p_9_7_pi2j c_9_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04939 c_9_7_s1_s c_9_7_a p_9_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04938 c_10_5_a c_9_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04937 vss c_9_7_s1_s n9821 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04936 n9834 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04935 vss a_5 n9577 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04934 n9577 p_9_2_d2j n9828 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04933 n9828 p_9_2_d2jbar n9579 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04932 n9579 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04931 vss p_9_7_t_s p_9_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04930 p_9_7_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04929 n9828 n9834 p_9_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04928 p_9_7_t_s n9828 n9834 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04927 n10203 p_9_2_d2j n10029 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04926 n10028 p_9_2_d2jbar n10203 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04925 p_9_6_t_s n10203 n10202 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04924 n10203 n10202 p_9_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04923 p_9_6_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04922 vss p_9_6_t_s p_9_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04921 n10202 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04920 vss a_5 n10028 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04919 n10029 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04918 vss c_9_6_s1_s n10027 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04917 c_10_4_a c_9_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04916 c_9_6_s1_s p_9_6_pi2j c_9_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04915 c_9_6_s2_s n10027 c_8_7_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04914 n10027 c_8_7_cout c_9_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04913 vss p_9_6_pi2j n10194 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04912 n10194 c_9_6_a n10195 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04911 n10195 c_8_7_cout n10196 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04910 vss p_9_6_pi2j n10196 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04909 n10196 c_9_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04908 vss n10195 c_10_5_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04907 p_9_6_pi2j c_9_6_a c_9_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04906 vss n10611 c_9_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04905 n10384 c_9_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04904 vss c_9_5_a n10384 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04903 n10611 c_9_5_cin n10384 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04902 n10193 c_9_5_b n10611 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04901 vss c_9_5_a n10193 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04900 n10388 c_9_5_cin c_9_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04899 c_9_5_s2_s n10388 c_9_5_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04898 c_9_5_a c_9_5_b c_9_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04897 c_9_5_s1_s c_9_5_a c_9_5_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04896 c_10_3_a c_9_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04895 vss c_9_5_s1_s n10388 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04894 n10617 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04893 vss a_3 n10204 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04892 n10204 p_9_2_d2j n10614 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04891 n10614 p_9_2_d2jbar n10205 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04890 n10205 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04889 vss p_9_5_t_s c_9_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04888 c_9_5_b p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04887 n10614 n10617 p_9_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04886 p_9_5_t_s n10614 n10617 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04885 n10822 p_9_2_d2j n10824 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04884 n10823 p_9_2_d2jbar n10822 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04883 p_9_4_t_s n10822 n10821 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04882 n10822 n10821 p_9_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04881 p_9_4_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04880 vss p_9_4_t_s p_9_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04879 n10821 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04878 vss a_3 n10823 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04877 n10824 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04876 vss c_9_4_s1_s n10820 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04875 c_10_2_a c_9_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04874 c_9_4_s1_s p_9_4_pi2j c_9_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04873 c_9_4_s2_s n10820 c_8_5_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04872 n10820 c_8_5_cout c_9_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04871 vss p_9_4_pi2j n10974 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04870 n10974 c_9_4_a n10815 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04869 n10815 c_8_5_cout n10975 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04868 vss p_9_4_pi2j n10975 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04867 n10975 c_9_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04866 vss n10815 c_10_3_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04865 p_9_4_pi2j c_9_4_a c_9_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04864 vss n11168 c_9_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04863 n10973 c_9_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04862 vss c_9_3_a n10973 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04861 n11168 c_9_3_cin n10973 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04860 n10972 c_9_3_b n11168 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04859 vss c_9_3_a n10972 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04858 n11170 c_9_3_cin c_9_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04857 c_9_3_s2_s n11170 c_9_3_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04856 c_9_3_a c_9_3_b c_9_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04855 c_9_3_s1_s c_9_3_a c_9_3_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04854 c_10_1_a c_9_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04853 vss c_9_3_s1_s n11170 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04852 n11174 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04851 vss a_1 n10979 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04850 n10979 p_9_2_d2j n11173 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04849 n11173 p_9_2_d2jbar n10980 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04848 n10980 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04847 vss p_9_3_t_s c_9_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04846 c_9_3_b p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04845 n11173 n11174 p_9_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04844 p_9_3_t_s n11173 n11174 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04843 n11599 p_9_2_d2j n11601 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04842 n11600 p_9_2_d2jbar n11599 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04841 p_9_2_t_s n11599 n11597 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04840 n11599 n11597 p_9_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04839 c_9_2_b p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04838 vss p_9_2_t_s c_9_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04837 n11597 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04836 vss a_1 n11600 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04835 n11601 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04834 vss c_9_2_s1_s n11596 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04833 c_9_2_sum c_9_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04832 c_9_2_s1_s c_9_2_b c_9_2_a vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04831 c_9_2_s2_s n11596 c_8_3_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04830 n11596 c_8_3_cout c_9_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04829 vss c_9_2_b n11589 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04828 n11589 c_9_2_a n11590 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04827 n11590 c_8_3_cout n11591 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04826 vss c_9_2_b n11591 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04825 n11591 c_9_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04824 vss n11590 c_10_1_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04823 c_9_2_b c_9_2_a c_9_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04822 vss n11947 c_9_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04821 n11735 p_9_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04820 vss c_9_1_a n11735 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04819 n11947 c_9_1_cin n11735 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04818 n11734 p_9_1_pi2j n11947 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04817 vss c_9_1_a n11734 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04816 n11944 c_9_1_cin c_9_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04815 c_9_1_s2_s n11944 c_9_1_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04814 c_9_1_a p_9_1_pi2j c_9_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04813 c_9_1_s1_s c_9_1_a p_9_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04812 c_9_1_sum c_9_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04811 vss c_9_1_s1_s n11944 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04810 n11957 p_9_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04809 n11958 p_9_2_d2jbar n11738 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04808 n11738 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04807 vss p_9_1_t_s p_9_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04806 p_9_1_pi2j p_9_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04805 n11958 n11957 p_9_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04804 p_9_1_t_s n11958 n11957 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04803 cl4_9_s1_s n12323 c_8_1_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04802 n12323 c_8_1_sum cl4_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04801 vss cl4_9_s1_s p_12 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04800 vss c_8_1_sum n12313 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04799 n12313 n12323 n12312 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04798 n12311 n12312 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04797 n12310 c_8_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_04796 vss c_8_2_sum n12310 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_04795 n12307 c_8_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04794 n12309 c_8_1_cout n12307 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04793 n12308 c_8_1_sum n12309 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04792 n12310 n12323 n12308 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04791 n12305 n12309 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04790 cl4_9_s2_s c_8_1_cout c_8_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04789 c_8_1_cout c_8_2_sum cl4_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04788 vss cl4_9_s2_s n12304 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04787 cl4_9_s3_s n12304 n12311 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04786 n12304 n12311 cl4_9_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04785 vss cl4_9_s3_s p_13 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04784 vss c_8_33_s1_s n181 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04783 c_9_31_a c_8_33_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04782 c_8_33_s1_s c_8_31_a p_8_33_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04781 c_8_31_a p_8_33_pi2j c_8_33_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04780 c_8_33_s2_s n181 c_8_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04779 n181 c_8_32_cin c_8_33_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04778 vss c_8_31_a n23 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04777 n23 p_8_33_pi2j n178 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04776 n178 c_8_32_cin n24 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04775 vss c_8_31_a n24 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04774 n24 p_8_33_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04773 vss n178 c_9_32_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04772 n186 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04771 n187 a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04770 vss p_8_33_t_s p_8_33_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04769 p_8_33_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04768 n187 n186 p_8_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04767 p_8_33_t_s n187 n186 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04766 n529 p_8_2_d2j n527 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04765 n528 p_8_2_d2jbar n529 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04764 p_8_32_t_s n529 n526 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04763 n529 n526 p_8_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04762 p_8_32_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04761 vss p_8_32_t_s p_8_32_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04760 n526 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04759 vss a_31 n528 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04758 n527 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04757 vss c_8_32_s1_s n522 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04756 c_9_30_a c_8_32_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04755 c_8_32_s1_s p_8_32_pi2j c_8_31_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04754 c_8_32_s2_s n522 c_8_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04753 n522 c_8_32_cin c_8_32_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04752 vss p_8_32_pi2j n519 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04751 n519 c_8_31_a n517 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04750 n517 c_8_32_cin n518 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04749 vss p_8_32_pi2j n518 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04748 n518 c_8_31_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04747 vss n517 c_9_31_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04746 p_8_32_pi2j c_8_31_a c_8_32_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04745 vss n871 c_8_31_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04744 n642 p_8_31_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04743 vss c_8_31_a n642 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04742 n871 c_8_31_cin n642 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04741 n641 p_8_31_pi2j n871 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04740 vss c_8_31_a n641 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04739 n868 c_8_31_cin c_8_31_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04738 c_8_31_s2_s n868 c_8_31_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04737 c_8_31_a p_8_31_pi2j c_8_31_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04736 c_8_31_s1_s c_8_31_a p_8_31_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04735 c_9_29_a c_8_31_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04734 vss c_8_31_s1_s n868 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04733 n878 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04732 vss a_29 n644 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04731 n644 p_8_2_d2j n875 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04730 n875 p_8_2_d2jbar n643 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04729 n643 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04728 vss p_8_31_t_s p_8_31_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04727 p_8_31_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04726 n875 n878 p_8_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04725 p_8_31_t_s n875 n878 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04724 n1286 p_8_2_d2j n1284 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04723 n1285 p_8_2_d2jbar n1286 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04722 p_8_30_t_s n1286 n1283 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04721 n1286 n1283 p_8_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04720 p_8_30_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04719 vss p_8_30_t_s p_8_30_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04718 n1283 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04717 vss a_29 n1285 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04716 n1284 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04715 vss c_8_30_s1_s n1280 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04714 c_9_28_a c_8_30_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04713 c_8_30_s1_s p_8_30_pi2j c_8_30_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04712 c_8_30_s2_s n1280 c_6_31_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04711 n1280 c_6_31_cout c_8_30_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04710 vss p_8_30_pi2j n1274 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04709 n1274 c_8_30_a n1275 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04708 n1275 c_6_31_cout n1273 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04707 vss p_8_30_pi2j n1273 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04706 n1273 c_8_30_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04705 vss n1275 c_9_29_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04704 p_8_30_pi2j c_8_30_a c_8_30_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04703 vss n1649 c_8_29_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04702 n1406 p_8_29_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04701 vss c_8_29_a n1406 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04700 n1649 c_8_29_cin n1406 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04699 n1272 p_8_29_pi2j n1649 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04698 vss c_8_29_a n1272 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04697 n1644 c_8_29_cin c_8_29_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04696 c_8_29_s2_s n1644 c_8_29_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04695 c_8_29_a p_8_29_pi2j c_8_29_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04694 c_8_29_s1_s c_8_29_a p_8_29_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04693 c_9_27_a c_8_29_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04692 vss c_8_29_s1_s n1644 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04691 n1656 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04690 vss a_27 n1408 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04689 n1408 p_8_2_d2j n1654 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04688 n1654 p_8_2_d2jbar n1407 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04687 n1407 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04686 vss p_8_29_t_s p_8_29_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04685 p_8_29_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04684 n1654 n1656 p_8_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04683 p_8_29_t_s n1654 n1656 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04682 n2039 p_8_2_d2j n2037 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04681 n2038 p_8_2_d2jbar n2039 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04680 p_8_28_t_s n2039 n2040 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04679 n2039 n2040 p_8_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04678 p_8_28_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04677 vss p_8_28_t_s p_8_28_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04676 n2040 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04675 vss a_27 n2038 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04674 n2037 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04673 vss c_8_28_s1_s n1838 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04672 c_9_26_a c_8_28_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04671 c_8_28_s1_s p_8_28_pi2j c_8_28_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04670 c_8_28_s2_s n1838 c_6_29_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04669 n1838 c_6_29_cout c_8_28_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04668 vss p_8_28_pi2j n2029 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04667 n2029 c_8_28_a n2031 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04666 n2031 c_6_29_cout n2030 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04665 vss p_8_28_pi2j n2030 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04664 n2030 c_8_28_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04663 vss n2031 c_9_27_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04662 p_8_28_pi2j c_8_28_a c_8_28_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04661 vss n2461 c_8_27_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04660 n2197 c_8_27_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04659 vss c_8_27_a n2197 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04658 n2461 c_8_27_cin n2197 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04657 n2028 c_8_27_b n2461 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04656 vss c_8_27_a n2028 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04655 n2451 c_8_27_cin c_8_27_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04654 c_8_27_s2_s n2451 c_8_27_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04653 c_8_27_a c_8_27_b c_8_27_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04652 c_8_27_s1_s c_8_27_a c_8_27_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04651 c_9_25_a c_8_27_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04650 vss c_8_27_s1_s n2451 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04649 n2466 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04648 vss a_25 n2202 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04647 n2202 p_8_2_d2j n2462 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04646 n2462 p_8_2_d2jbar n2203 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04645 n2203 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04644 vss p_8_27_t_s c_8_27_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04643 c_8_27_b p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04642 n2462 n2466 p_8_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04641 p_8_27_t_s n2462 n2466 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04640 n2667 p_8_2_d2j n2665 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04639 n2666 p_8_2_d2jbar n2667 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04638 p_8_26_t_s n2667 n2664 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04637 n2667 n2664 p_8_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04636 p_8_26_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04635 vss p_8_26_t_s p_8_26_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04634 n2664 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04633 vss a_25 n2666 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04632 n2665 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04631 vss c_8_26_s1_s n2663 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04630 c_9_24_a c_8_26_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04629 c_8_26_s1_s p_8_26_pi2j c_8_26_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04628 c_8_26_s2_s n2663 c_6_27_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04627 n2663 c_6_27_cout c_8_26_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04626 vss p_8_26_pi2j n2847 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04625 n2847 c_8_26_a n2845 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04624 n2845 c_6_27_cout n2842 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04623 vss p_8_26_pi2j n2842 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04622 n2842 c_8_26_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04621 vss n2845 c_9_25_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04620 p_8_26_pi2j c_8_26_a c_8_26_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04619 vss n3254 c_8_25_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04618 n2846 c_8_25_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04617 vss c_8_25_a n2846 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04616 n3254 c_8_25_cin n2846 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04615 n2844 c_8_25_b n3254 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04614 vss c_8_25_a n2844 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04613 n3022 c_8_25_cin c_8_25_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04612 c_8_25_s2_s n3022 c_8_25_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04611 c_8_25_a c_8_25_b c_8_25_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04610 c_8_25_s1_s c_8_25_a c_8_25_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04609 c_9_23_a c_8_25_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04608 vss c_8_25_s1_s n3022 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04607 n3257 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04606 vss a_23 n2853 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04605 n2853 p_8_2_d2j n3024 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04604 n3024 p_8_2_d2jbar n2852 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04603 n2852 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04602 vss p_8_25_t_s c_8_25_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04601 c_8_25_b p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04600 n3024 n3257 p_8_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04599 p_8_25_t_s n3024 n3257 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04598 n3462 p_8_2_d2j n3460 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04597 n3461 p_8_2_d2jbar n3462 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04596 p_8_24_t_s n3462 n3459 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04595 n3462 n3459 p_8_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04594 c_8_24_b p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04593 vss p_8_24_t_s c_8_24_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04592 n3459 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04591 vss a_23 n3461 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04590 n3460 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04589 vss c_8_24_s1_s n3456 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04588 c_9_22_a c_8_24_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04587 c_8_24_s1_s c_8_24_b c_8_24_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04586 c_8_24_s2_s n3456 c_6_25_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04585 n3456 c_6_25_cout c_8_24_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04584 vss c_8_24_b n3611 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04583 n3611 c_8_24_a n3452 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04582 n3452 c_6_25_cout n3607 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04581 vss c_8_24_b n3607 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04580 n3607 c_8_24_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04579 vss n3452 c_9_23_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04578 c_8_24_b c_8_24_a c_8_24_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04577 vss n3843 c_8_23_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04576 n3610 c_8_23_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04575 vss c_8_23_a n3610 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04574 n3843 c_8_23_cin n3610 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04573 n3609 c_8_23_b n3843 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04572 vss c_8_23_a n3609 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04571 n3844 c_8_23_cin c_8_23_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04570 c_8_23_s2_s n3844 c_8_23_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04569 c_8_23_a c_8_23_b c_8_23_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04568 c_8_23_s1_s c_8_23_a c_8_23_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04567 c_9_21_a c_8_23_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04566 vss c_8_23_s1_s n3844 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04565 n3850 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04564 vss a_21 n3615 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04563 n3615 p_8_2_d2j n3847 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04562 n3847 p_8_2_d2jbar n3614 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04561 n3614 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04560 vss p_8_23_t_s c_8_23_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04559 c_8_23_b p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04558 n3847 n3850 p_8_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04557 p_8_23_t_s n3847 n3850 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04556 n4267 p_8_2_d2j n4265 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04555 n4266 p_8_2_d2jbar n4267 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04554 p_8_22_t_s n4267 n4264 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04553 n4267 n4264 p_8_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04552 p_8_22_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04551 vss p_8_22_t_s p_8_22_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04550 n4264 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04549 vss a_21 n4266 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04548 n4265 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04547 vss c_8_22_s1_s n4259 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04546 c_9_20_a c_8_22_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04545 c_8_22_s1_s p_8_22_pi2j c_8_22_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04544 c_8_22_s2_s n4259 c_6_23_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04543 n4259 c_6_23_cout c_8_22_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04542 vss p_8_22_pi2j n4256 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04541 n4256 c_8_22_a n4254 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04540 n4254 c_6_23_cout n4255 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04539 vss p_8_22_pi2j n4255 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04538 n4255 c_8_22_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04537 vss n4254 c_9_21_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04536 p_8_22_pi2j c_8_22_a c_8_22_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04535 vss n4617 c_8_21_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04534 n4393 p_8_21_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04533 vss c_8_21_a n4393 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04532 n4617 c_8_21_cin n4393 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04531 n4392 p_8_21_pi2j n4617 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04530 vss c_8_21_a n4392 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04529 n4613 c_8_21_cin c_8_21_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04528 c_8_21_s2_s n4613 c_8_21_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04527 c_8_21_a p_8_21_pi2j c_8_21_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04526 c_8_21_s1_s c_8_21_a p_8_21_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04525 c_9_19_a c_8_21_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04524 vss c_8_21_s1_s n4613 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04523 n4625 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04522 vss a_19 n4395 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04521 n4395 p_8_2_d2j n4622 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04520 n4622 p_8_2_d2jbar n4394 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04519 n4394 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04518 vss p_8_21_t_s p_8_21_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04517 p_8_21_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04516 n4622 n4625 p_8_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04515 p_8_21_t_s n4622 n4625 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04514 n5013 p_8_2_d2j n5011 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04513 n5012 p_8_2_d2jbar n5013 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04512 p_8_20_t_s n5013 n5010 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04511 n5013 n5010 p_8_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04510 p_8_20_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04509 vss p_8_20_t_s p_8_20_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04508 n5010 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04507 vss a_19 n5012 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04506 n5011 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04505 vss c_8_20_s1_s n5006 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04504 c_9_18_a c_8_20_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04503 c_8_20_s1_s p_8_20_pi2j c_8_20_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04502 c_8_20_s2_s n5006 c_6_21_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04501 n5006 c_6_21_cout c_8_20_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04500 vss p_8_20_pi2j n5001 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04499 n5001 c_8_20_a n5002 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04498 n5002 c_6_21_cout n5000 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04497 vss p_8_20_pi2j n5000 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04496 n5000 c_8_20_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04495 vss n5002 c_9_19_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04494 p_8_20_pi2j c_8_20_a c_8_20_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04493 vss n5376 c_8_19_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04492 n5133 p_8_19_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04491 vss c_8_19_a n5133 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04490 n5376 c_8_19_cin n5133 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04489 n5134 p_8_19_pi2j n5376 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04488 vss c_8_19_a n5134 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04487 n5371 c_8_19_cin c_8_19_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04486 c_8_19_s2_s n5371 c_8_19_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04485 c_8_19_a p_8_19_pi2j c_8_19_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04484 c_8_19_s1_s c_8_19_a p_8_19_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04483 c_9_17_a c_8_19_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04482 vss c_8_19_s1_s n5371 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04481 n5383 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04480 vss a_17 n5136 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04479 n5136 p_8_2_d2j n5381 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04478 n5381 p_8_2_d2jbar n5135 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04477 n5135 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04476 vss p_8_19_t_s p_8_19_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04475 p_8_19_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04474 n5381 n5383 p_8_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04473 p_8_19_t_s n5381 n5383 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04472 n5766 p_8_2_d2j n5765 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04471 n5763 p_8_2_d2jbar n5766 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04470 p_8_18_t_s n5766 n5764 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04469 n5766 n5764 p_8_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04468 p_8_18_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04467 vss p_8_18_t_s p_8_18_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04466 n5764 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04465 vss a_17 n5763 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04464 n5765 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04463 vss c_8_18_s1_s n5564 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04462 c_9_16_a c_8_18_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04461 c_8_18_s1_s p_8_18_pi2j c_8_18_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04460 c_8_18_s2_s n5564 c_6_19_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04459 n5564 c_6_19_cout c_8_18_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04458 vss p_8_18_pi2j n5755 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04457 n5755 c_8_18_a n5757 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04456 n5757 c_6_19_cout n5756 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04455 vss p_8_18_pi2j n5756 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04454 n5756 c_8_18_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04453 vss n5757 c_9_17_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04452 p_8_18_pi2j c_8_18_a c_8_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04451 vss n6167 c_8_17_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04450 n5902 p_8_17_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04449 vss c_8_17_a n5902 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04448 n6167 c_8_17_cin n5902 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04447 n5754 p_8_17_pi2j n6167 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04446 vss c_8_17_a n5754 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04445 n6156 c_8_17_cin c_8_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04444 c_8_17_s2_s n6156 c_8_17_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04443 c_8_17_a p_8_17_pi2j c_8_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04442 c_8_17_s1_s c_8_17_a p_8_17_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04441 c_9_15_a c_8_17_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04440 vss c_8_17_s1_s n6156 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04439 n6173 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04438 vss a_15 n5905 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04437 n5905 p_8_2_d2j n6168 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04436 n6168 p_8_2_d2jbar n5906 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04435 n5906 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04434 vss p_8_17_t_s p_8_17_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04433 p_8_17_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04432 n6168 n6173 p_8_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04431 p_8_17_t_s n6168 n6173 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04430 n6368 p_8_2_d2j n6366 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04429 n6367 p_8_2_d2jbar n6368 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04428 p_8_16_t_s n6368 n6546 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04427 n6368 n6546 p_8_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04426 p_8_16_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04425 vss p_8_16_t_s p_8_16_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04424 n6546 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04423 vss a_15 n6367 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04422 n6366 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04421 vss c_8_16_s1_s n6365 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04420 c_9_14_a c_8_16_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04419 c_8_16_s1_s p_8_16_pi2j c_8_16_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04418 c_8_16_s2_s n6365 c_6_17_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04417 n6365 c_6_17_cout c_8_16_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04416 vss p_8_16_pi2j n6541 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04415 n6541 c_8_16_a n6540 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04414 n6540 c_6_17_cout n6536 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04413 vss p_8_16_pi2j n6536 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04412 n6536 c_8_16_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04411 vss n6540 c_9_15_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04410 p_8_16_pi2j c_8_16_a c_8_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04409 vss n6955 c_8_15_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04408 n6538 c_8_15_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04407 vss c_8_15_a n6538 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04406 n6955 c_8_15_cin n6538 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04405 n6539 c_8_15_b n6955 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04404 vss c_8_15_a n6539 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04403 n6723 c_8_15_cin c_8_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04402 c_8_15_s2_s n6723 c_8_15_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04401 c_8_15_a c_8_15_b c_8_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04400 c_8_15_s1_s c_8_15_a c_8_15_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04399 c_9_13_a c_8_15_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04398 vss c_8_15_s1_s n6723 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04397 n6959 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04396 vss a_13 n6548 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04395 n6548 p_8_2_d2j n6725 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04394 n6725 p_8_2_d2jbar n6547 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04393 n6547 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04392 vss p_8_15_t_s c_8_15_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04391 c_8_15_b p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04390 n6725 n6959 p_8_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04389 p_8_15_t_s n6725 n6959 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04388 n7160 p_8_2_d2j n7158 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04387 n7159 p_8_2_d2jbar n7160 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04386 p_8_14_t_s n7160 n7157 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04385 n7160 n7157 p_8_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04384 p_8_14_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04383 vss p_8_14_t_s p_8_14_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04382 n7157 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04381 vss a_13 n7159 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04380 n7158 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04379 vss c_8_14_s1_s n7154 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04378 c_9_12_a c_8_14_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04377 c_8_14_s1_s p_8_14_pi2j c_8_14_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04376 c_8_14_s2_s n7154 c_6_15_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04375 n7154 c_6_15_cout c_8_14_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04374 vss p_8_14_pi2j n7317 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04373 n7317 c_8_14_a n7151 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04372 n7151 c_6_15_cout n7313 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04371 vss p_8_14_pi2j n7313 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04370 n7313 c_8_14_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04369 vss n7151 c_9_13_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04368 p_8_14_pi2j c_8_14_a c_8_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04367 vss n7517 c_8_13_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04366 n7316 c_8_13_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04365 vss c_8_13_a n7316 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04364 n7517 c_8_13_cin n7316 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04363 n7315 c_8_13_b n7517 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04362 vss c_8_13_a n7315 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04361 n7519 c_8_13_cin c_8_13_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04360 c_8_13_s2_s n7519 c_8_13_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04359 c_8_13_a c_8_13_b c_8_13_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04358 c_8_13_s1_s c_8_13_a c_8_13_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04357 c_9_11_a c_8_13_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04356 vss c_8_13_s1_s n7519 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04355 n7524 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04354 vss a_11 n7321 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04353 n7321 p_8_2_d2j n7521 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04352 n7521 p_8_2_d2jbar n7320 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04351 n7320 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04350 vss p_8_13_t_s c_8_13_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04349 c_8_13_b p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04348 n7521 n7524 p_8_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04347 p_8_13_t_s n7521 n7524 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04346 n7951 p_8_2_d2j n7949 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04345 n7950 p_8_2_d2jbar n7951 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04344 p_8_12_t_s n7951 n7948 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04343 n7951 n7948 p_8_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04342 c_8_12_b p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04341 vss p_8_12_t_s c_8_12_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04340 n7948 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04339 vss a_11 n7950 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04338 n7949 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04337 vss c_8_12_s1_s n7944 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04336 c_9_10_a c_8_12_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04335 c_8_12_s1_s c_8_12_b c_8_12_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04334 c_8_12_s2_s n7944 c_6_13_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04333 n7944 c_6_13_cout c_8_12_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04332 vss c_8_12_b n7939 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04331 n7939 c_8_12_a n7941 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04330 n7941 c_6_13_cout n7940 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04329 vss c_8_12_b n7940 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04328 n7940 c_8_12_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04327 vss n7941 c_9_11_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04326 c_8_12_b c_8_12_a c_8_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04325 vss n8306 c_8_11_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04324 n8078 p_8_11_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04323 vss c_8_11_a n8078 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04322 n8306 c_8_11_cin n8078 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04321 n8077 p_8_11_pi2j n8306 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04320 vss c_8_11_a n8077 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04319 n8301 c_8_11_cin c_8_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04318 c_8_11_s2_s n8301 c_8_11_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04317 c_8_11_a p_8_11_pi2j c_8_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04316 c_8_11_s1_s c_8_11_a p_8_11_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04315 c_9_9_a c_8_11_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04314 vss c_8_11_s1_s n8301 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04313 n8313 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04312 vss a_9 n8081 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04311 n8081 p_8_2_d2j n8310 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04310 n8310 p_8_2_d2jbar n8080 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04309 n8080 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04308 vss p_8_11_t_s p_8_11_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04307 p_8_11_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04306 n8310 n8313 p_8_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04305 p_8_11_t_s n8310 n8313 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04304 n8702 p_8_2_d2j n8700 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04303 n8701 p_8_2_d2jbar n8702 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04302 p_8_10_t_s n8702 n8699 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04301 n8702 n8699 p_8_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04300 p_8_10_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04299 vss p_8_10_t_s p_8_10_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04298 n8699 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04297 vss a_9 n8701 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04296 n8700 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04295 vss c_8_10_s1_s n8696 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04294 c_9_8_a c_8_10_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04293 c_8_10_s1_s p_8_10_pi2j c_8_10_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04292 c_8_10_s2_s n8696 c_6_11_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04291 n8696 c_6_11_cout c_8_10_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04290 vss p_8_10_pi2j n8690 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04289 n8690 c_8_10_a n8691 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04288 n8691 c_6_11_cout n8689 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04287 vss p_8_10_pi2j n8689 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04286 n8689 c_8_10_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04285 vss n8691 c_9_9_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04284 p_8_10_pi2j c_8_10_a c_8_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04283 vss n9064 c_8_9_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04282 n8826 p_8_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04281 vss c_8_9_a n8826 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04280 n9064 c_8_9_cin n8826 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04279 n8825 p_8_9_pi2j n9064 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04278 vss c_8_9_a n8825 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04277 n9059 c_8_9_cin c_8_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04276 c_8_9_s2_s n9059 c_8_9_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04275 c_8_9_a p_8_9_pi2j c_8_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04274 c_8_9_s1_s c_8_9_a p_8_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04273 c_9_7_a c_8_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04272 vss c_8_9_s1_s n9059 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04271 n9071 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04270 vss a_7 n8828 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04269 n8828 p_8_2_d2j n9069 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04268 n9069 p_8_2_d2jbar n8827 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04267 n8827 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04266 vss p_8_9_t_s p_8_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04265 p_8_9_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04264 n9069 n9071 p_8_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04263 p_8_9_t_s n9069 n9071 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04262 n9443 p_8_2_d2j n9442 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04261 n9440 p_8_2_d2jbar n9443 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04260 p_8_8_t_s n9443 n9441 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04259 n9443 n9441 p_8_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04258 p_8_8_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04257 vss p_8_8_t_s p_8_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04256 n9441 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04255 vss a_7 n9440 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04254 n9442 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04253 vss c_8_8_s1_s n9429 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04252 c_9_6_a c_8_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04251 c_8_8_s1_s p_8_8_pi2j c_8_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04250 c_8_8_s2_s n9429 c_6_9_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04249 n9429 c_6_9_cout c_8_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04248 vss p_8_8_pi2j n9433 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04247 n9433 c_8_8_a n9432 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04246 n9432 c_6_9_cout n9434 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04245 vss p_8_8_pi2j n9434 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04244 n9434 c_8_8_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04243 vss n9432 c_9_7_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04242 p_8_8_pi2j c_8_8_a c_8_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04241 vss n9851 c_8_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04240 n9580 p_8_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04239 vss c_8_7_a n9580 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04238 n9851 c_8_7_cin n9580 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04237 n9431 p_8_7_pi2j n9851 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04236 vss c_8_7_a n9431 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04235 n9846 c_8_7_cin c_8_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04234 c_8_7_s2_s n9846 c_8_7_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04233 c_8_7_a p_8_7_pi2j c_8_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04232 c_8_7_s1_s c_8_7_a p_8_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04231 c_9_5_a c_8_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04230 vss c_8_7_s1_s n9846 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04229 n9857 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04228 vss a_5 n9584 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04227 n9584 p_8_2_d2j n9852 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04226 n9852 p_8_2_d2jbar n9583 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04225 n9583 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04224 vss p_8_7_t_s p_8_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04223 p_8_7_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04222 n9852 n9857 p_8_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04221 p_8_7_t_s n9852 n9857 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04220 n10215 p_8_2_d2j n10033 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04219 n10034 p_8_2_d2jbar n10215 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04218 p_8_6_t_s n10215 n10217 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04217 n10215 n10217 p_8_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04216 p_8_6_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04215 vss p_8_6_t_s p_8_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04214 n10217 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04213 vss a_5 n10034 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04212 n10033 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04211 vss c_8_6_s1_s n10032 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04210 c_9_4_a c_8_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04209 c_8_6_s1_s p_8_6_pi2j c_8_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04208 c_8_6_s2_s n10032 c_6_7_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04207 n10032 c_6_7_cout c_8_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04206 vss p_8_6_pi2j n10211 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04205 n10211 c_8_6_a n10210 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04204 n10210 c_6_7_cout n10206 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04203 vss p_8_6_pi2j n10206 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04202 n10206 c_8_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04201 vss n10210 c_9_5_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04200 p_8_6_pi2j c_8_6_a c_8_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04199 vss n10631 c_8_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04198 n10393 c_8_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04197 vss c_8_5_a n10393 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04196 n10631 c_8_5_cin n10393 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04195 n10209 c_8_5_b n10631 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04194 vss c_8_5_a n10209 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04193 n10398 c_8_5_cin c_8_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04192 c_8_5_s2_s n10398 c_8_5_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04191 c_8_5_a c_8_5_b c_8_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04190 c_8_5_s1_s c_8_5_a c_8_5_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04189 c_9_3_a c_8_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04188 vss c_8_5_s1_s n10398 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04187 n10635 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04186 vss a_3 n10219 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04185 n10219 p_8_2_d2j n10632 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04184 n10632 p_8_2_d2jbar n10218 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04183 n10218 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04182 vss p_8_5_t_s c_8_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04181 c_8_5_b p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04180 n10632 n10635 p_8_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04179 p_8_5_t_s n10632 n10635 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04178 n10834 p_8_2_d2j n10832 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04177 n10833 p_8_2_d2jbar n10834 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04176 p_8_4_t_s n10834 n10831 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04175 n10834 n10831 p_8_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04174 p_8_4_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04173 vss p_8_4_t_s p_8_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04172 n10831 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04171 vss a_3 n10833 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04170 n10832 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04169 vss c_8_4_s1_s n10830 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04168 c_9_2_a c_8_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04167 c_8_4_s1_s p_8_4_pi2j c_8_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04166 c_8_4_s2_s n10830 c_6_5_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04165 n10830 c_6_5_cout c_8_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04164 vss p_8_4_pi2j n10985 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04163 n10985 c_8_4_a n10825 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04162 n10825 c_6_5_cout n10981 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04161 vss p_8_4_pi2j n10981 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04160 n10981 c_8_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04159 vss n10825 c_9_3_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04158 p_8_4_pi2j c_8_4_a c_8_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04157 vss n11182 c_8_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04156 n10984 c_8_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04155 vss c_8_3_a n10984 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04154 n11182 c_8_3_cin n10984 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04153 n10983 c_8_3_b n11182 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04152 vss c_8_3_a n10983 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04151 n11184 c_8_3_cin c_8_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04150 c_8_3_s2_s n11184 c_8_3_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04149 c_8_3_a c_8_3_b c_8_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04148 c_8_3_s1_s c_8_3_a c_8_3_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04147 c_9_1_a c_8_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04146 vss c_8_3_s1_s n11184 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04145 n11189 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04144 vss a_1 n10989 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04143 n10989 p_8_2_d2j n11186 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04142 n11186 p_8_2_d2jbar n10988 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04141 n10988 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04140 vss p_8_3_t_s c_8_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04139 c_8_3_b p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04138 n11186 n11189 p_8_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04137 p_8_3_t_s n11186 n11189 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04136 n11614 p_8_2_d2j n11612 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04135 n11613 p_8_2_d2jbar n11614 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04134 p_8_2_t_s n11614 n11611 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04133 n11614 n11611 p_8_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04132 c_8_2_b p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04131 vss p_8_2_t_s c_8_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04130 n11611 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04129 vss a_1 n11613 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04128 n11612 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04127 vss c_8_2_s1_s n11607 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04126 c_8_2_sum c_8_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04125 c_8_2_s1_s c_8_2_b c_8_2_a vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04124 c_8_2_s2_s n11607 c_6_3_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04123 n11607 c_6_3_cout c_8_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04122 vss c_8_2_b n11602 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04121 n11602 c_8_2_a n11604 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04120 n11604 c_6_3_cout n11603 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04119 vss c_8_2_b n11603 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04118 n11603 c_8_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04117 vss n11604 c_9_1_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04116 c_8_2_b c_8_2_a c_8_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04115 vss n11968 c_8_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04114 n11740 p_8_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04113 vss c_8_1_a n11740 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04112 n11968 c_8_1_cin n11740 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04111 n11739 p_8_1_pi2j n11968 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04110 vss c_8_1_a n11739 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04109 n11967 c_8_1_cin c_8_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04108 c_8_1_s2_s n11967 c_8_1_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04107 c_8_1_a p_8_1_pi2j c_8_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04106 c_8_1_s1_s c_8_1_a p_8_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04105 c_8_1_sum c_8_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04104 vss c_8_1_s1_s n11967 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04103 n11977 p_8_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04102 n11978 p_8_2_d2jbar n11743 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04101 n11743 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04100 vss p_8_1_t_s p_8_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04099 p_8_1_pi2j p_8_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04098 n11978 n11977 p_8_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04097 p_8_1_t_s n11978 n11977 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04096 cl4_8_s1_s n12339 c_6_1_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04095 n12339 c_6_1_sum cl4_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04094 vss cl4_8_s1_s p_10 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04093 vss c_6_1_sum n12330 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04092 n12330 n12339 n12329 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04091 n12328 n12329 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04090 n12327 c_6_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_04089 vss c_6_2_sum n12327 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_04088 n12326 c_6_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04087 n12324 c_6_1_cout n12326 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04086 n12322 c_6_1_sum n12324 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04085 n12327 n12339 n12322 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04084 n12323 n12324 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04083 cl4_8_s2_s c_6_1_cout c_6_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04082 c_6_1_cout c_6_2_sum cl4_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04081 vss cl4_8_s2_s n12320 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04080 cl4_8_s3_s n12320 n12328 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04079 n12320 n12328 cl4_8_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04078 vss cl4_8_s3_s p_11 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_04077 vss c_6_33_s1_s n191 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04076 c_8_31_a c_6_33_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04075 c_6_33_s1_s c_6_31_a p_6_33_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04074 c_6_31_a p_6_33_pi2j c_6_33_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04073 c_6_33_s2_s n191 c_6_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04072 n191 c_6_32_cin c_6_33_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04071 vss c_6_31_a n25 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04070 n25 p_6_33_pi2j n190 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04069 n190 c_6_32_cin n26 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04068 vss c_6_31_a n26 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04067 n26 p_6_33_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04066 vss n190 c_8_32_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04065 n198 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04064 n201 a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04063 vss p_6_33_t_s p_6_33_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04062 p_6_33_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04061 n201 n198 p_6_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04060 p_6_33_t_s n201 n198 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04059 n541 p_6_2_d2j n542 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04058 n540 p_6_2_d2jbar n541 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04057 p_6_32_t_s n541 n538 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04056 n541 n538 p_6_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04055 p_6_32_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04054 vss p_6_32_t_s p_6_32_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04053 n538 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04052 vss a_31 n540 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04051 n542 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04050 vss c_6_32_s1_s n535 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04049 c_8_30_a c_6_32_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04048 c_6_32_s1_s p_6_32_pi2j c_6_31_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04047 c_6_32_s2_s n535 c_6_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04046 n535 c_6_32_cin c_6_32_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04045 vss p_6_32_pi2j n531 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04044 n531 c_6_31_a n530 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04043 n530 c_6_32_cin n532 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04042 vss p_6_32_pi2j n532 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04041 n532 c_6_31_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04040 vss n530 c_8_31_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04039 p_6_32_pi2j c_6_31_a c_6_32_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04038 vss n887 c_6_31_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_04037 n646 p_6_31_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04036 vss c_6_31_a n646 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04035 n887 c_6_31_cin n646 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04034 n645 p_6_31_pi2j n887 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04033 vss c_6_31_a n645 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_04032 n883 c_6_31_cin c_6_31_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04031 c_6_31_s2_s n883 c_6_31_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04030 c_6_31_a p_6_31_pi2j c_6_31_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04029 c_6_31_s1_s c_6_31_a p_6_31_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04028 c_8_29_a c_6_31_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04027 vss c_6_31_s1_s n883 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04026 n893 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04025 vss a_29 n648 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04024 n648 p_6_2_d2j n895 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04023 n895 p_6_2_d2jbar n647 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04022 n647 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04021 vss p_6_31_t_s p_6_31_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04020 p_6_31_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04019 n895 n893 p_6_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04018 p_6_31_t_s n895 n893 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04017 n1301 p_6_2_d2j n1300 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04016 n1299 p_6_2_d2jbar n1301 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_04015 p_6_30_t_s n1301 n1298 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04014 n1301 n1298 p_6_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04013 p_6_30_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04012 vss p_6_30_t_s p_6_30_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_04011 n1298 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_04010 vss a_29 n1299 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04009 n1300 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_04008 vss c_6_30_s1_s n1293 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_04007 c_8_28_a c_6_30_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_04006 c_6_30_s1_s p_6_30_pi2j c_6_30_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04005 c_6_30_s2_s n1293 c_5_31_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04004 n1293 c_5_31_cout c_6_30_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_04003 vss p_6_30_pi2j n1290 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04002 n1290 c_6_30_a n1288 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04001 n1288 c_5_31_cout n1289 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_04000 vss p_6_30_pi2j n1289 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03999 n1289 c_6_30_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03998 vss n1288 c_8_29_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03997 p_6_30_pi2j c_6_30_a c_6_30_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03996 vss n1666 c_6_29_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03995 n1409 p_6_29_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03994 vss c_6_29_a n1409 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03993 n1666 c_6_29_cin n1409 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03992 n1287 p_6_29_pi2j n1666 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03991 vss c_6_29_a n1287 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03990 n1661 c_6_29_cin c_6_29_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03989 c_6_29_s2_s n1661 c_6_29_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03988 c_6_29_a p_6_29_pi2j c_6_29_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03987 c_6_29_s1_s c_6_29_a p_6_29_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03986 c_8_27_a c_6_29_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03985 vss c_6_29_s1_s n1661 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03984 n1673 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03983 vss a_27 n1410 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03982 n1410 p_6_2_d2j n1675 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03981 n1675 p_6_2_d2jbar n1411 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03980 n1411 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03979 vss p_6_29_t_s p_6_29_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03978 p_6_29_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03977 n1675 n1673 p_6_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03976 p_6_29_t_s n1675 n1673 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03975 n2054 p_6_2_d2j n2053 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03974 n2052 p_6_2_d2jbar n2054 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03973 p_6_28_t_s n2054 n2051 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03972 n2054 n2051 p_6_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03971 p_6_28_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03970 vss p_6_28_t_s p_6_28_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03969 n2051 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03968 vss a_27 n2052 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03967 n2053 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03966 vss c_6_28_s1_s n1844 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03965 c_8_26_a c_6_28_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03964 c_6_28_s1_s p_6_28_pi2j c_6_28_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03963 c_6_28_s2_s n1844 c_5_29_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03962 n1844 c_5_29_cout c_6_28_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03961 vss p_6_28_pi2j n2043 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03960 n2043 c_6_28_a n2044 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03959 n2044 c_5_29_cout n2042 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03958 vss p_6_28_pi2j n2042 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03957 n2042 c_6_28_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03956 vss n2044 c_8_27_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03955 p_6_28_pi2j c_6_28_a c_6_28_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03954 vss n2478 c_6_27_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03953 n2204 c_6_27_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03952 vss c_6_27_a n2204 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03951 n2478 c_6_27_cin n2204 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03950 n2041 c_6_27_b n2478 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03949 vss c_6_27_a n2041 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03948 n2470 c_6_27_cin c_6_27_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03947 c_6_27_s2_s n2470 c_6_27_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03946 c_6_27_a c_6_27_b c_6_27_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03945 c_6_27_s1_s c_6_27_a c_6_27_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03944 c_8_25_a c_6_27_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03943 vss c_6_27_s1_s n2470 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03942 n2483 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03941 vss a_25 n2209 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03940 n2209 p_6_2_d2j n2479 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03939 n2479 p_6_2_d2jbar n2210 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03938 n2210 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03937 vss p_6_27_t_s c_6_27_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03936 c_6_27_b p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03935 n2479 n2483 p_6_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03934 p_6_27_t_s n2479 n2483 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03933 n2675 p_6_2_d2j n2673 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03932 n2674 p_6_2_d2jbar n2675 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03931 p_6_26_t_s n2675 n2672 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03930 n2675 n2672 p_6_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03929 p_6_26_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03928 vss p_6_26_t_s p_6_26_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03927 n2672 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03926 vss a_25 n2674 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03925 n2673 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03924 vss c_6_26_s1_s n2671 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03923 c_8_24_a c_6_26_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03922 c_6_26_s1_s p_6_26_pi2j c_6_26_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03921 c_6_26_s2_s n2671 c_5_27_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03920 n2671 c_5_27_cout c_6_26_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03919 vss p_6_26_pi2j n2858 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03918 n2858 c_6_26_a n2857 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03917 n2857 c_5_27_cout n2856 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03916 vss p_6_26_pi2j n2856 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03915 n2856 c_6_26_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03914 vss n2857 c_8_25_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03913 p_6_26_pi2j c_6_26_a c_6_26_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03912 vss n3266 c_6_25_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03911 n2855 c_6_25_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03910 vss c_6_25_a n2855 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03909 n3266 c_6_25_cin n2855 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03908 n2854 c_6_25_b n3266 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03907 vss c_6_25_a n2854 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03906 n3028 c_6_25_cin c_6_25_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03905 c_6_25_s2_s n3028 c_6_25_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03904 c_6_25_a c_6_25_b c_6_25_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03903 c_6_25_s1_s c_6_25_a c_6_25_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03902 c_8_23_a c_6_25_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03901 vss c_6_25_s1_s n3028 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03900 n3272 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03899 vss a_23 n2865 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03898 n2865 p_6_2_d2j n3034 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03897 n3034 p_6_2_d2jbar n2864 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03896 n2864 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03895 vss p_6_25_t_s c_6_25_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03894 c_6_25_b p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03893 n3034 n3272 p_6_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03892 p_6_25_t_s n3034 n3272 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03891 n3471 p_6_2_d2j n3473 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03890 n3472 p_6_2_d2jbar n3471 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03889 p_6_24_t_s n3471 n3470 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03888 n3471 n3470 p_6_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03887 c_6_24_b p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03886 vss p_6_24_t_s c_6_24_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03885 n3470 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03884 vss a_23 n3472 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03883 n3473 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03882 vss c_6_24_s1_s n3467 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03881 c_8_22_a c_6_24_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03880 c_6_24_s1_s c_6_24_b c_6_24_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03879 c_6_24_s2_s n3467 c_5_25_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03878 n3467 c_5_25_cout c_6_24_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03877 vss c_6_24_b n3618 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03876 n3618 c_6_24_a n3463 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03875 n3463 c_5_25_cout n3619 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03874 vss c_6_24_b n3619 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03873 n3619 c_6_24_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03872 vss n3463 c_8_23_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03871 c_6_24_b c_6_24_a c_6_24_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03870 vss n3855 c_6_23_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03869 n3617 c_6_23_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03868 vss c_6_23_a n3617 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03867 n3855 c_6_23_cin n3617 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03866 n3616 c_6_23_b n3855 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03865 vss c_6_23_a n3616 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03864 n3858 c_6_23_cin c_6_23_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03863 c_6_23_s2_s n3858 c_6_23_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03862 c_6_23_a c_6_23_b c_6_23_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03861 c_6_23_s1_s c_6_23_a c_6_23_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03860 c_8_21_a c_6_23_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03859 vss c_6_23_s1_s n3858 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03858 n3863 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03857 vss a_21 n3623 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03856 n3623 p_6_2_d2j n3865 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03855 n3865 p_6_2_d2jbar n3622 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03854 n3622 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03853 vss p_6_23_t_s c_6_23_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03852 c_6_23_b p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03851 n3865 n3863 p_6_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03850 p_6_23_t_s n3865 n3863 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03849 n4280 p_6_2_d2j n4281 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03848 n4279 p_6_2_d2jbar n4280 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03847 p_6_22_t_s n4280 n4278 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03846 n4280 n4278 p_6_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03845 p_6_22_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03844 vss p_6_22_t_s p_6_22_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03843 n4278 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03842 vss a_21 n4279 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03841 n4281 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03840 vss c_6_22_s1_s n4273 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03839 c_8_20_a c_6_22_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03838 c_6_22_s1_s p_6_22_pi2j c_6_22_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03837 c_6_22_s2_s n4273 c_5_23_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03836 n4273 c_5_23_cout c_6_22_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03835 vss p_6_22_pi2j n4269 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03834 n4269 c_6_22_a n4268 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03833 n4268 c_5_23_cout n4270 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03832 vss p_6_22_pi2j n4270 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03831 n4270 c_6_22_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03830 vss n4268 c_8_21_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03829 p_6_22_pi2j c_6_22_a c_6_22_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03828 vss n4632 c_6_21_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03827 n4397 p_6_21_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03826 vss c_6_21_a n4397 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03825 n4632 c_6_21_cin n4397 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03824 n4396 p_6_21_pi2j n4632 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03823 vss c_6_21_a n4396 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03822 n4628 c_6_21_cin c_6_21_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03821 c_6_21_s2_s n4628 c_6_21_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03820 c_6_21_a p_6_21_pi2j c_6_21_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03819 c_6_21_s1_s c_6_21_a p_6_21_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03818 c_8_19_a c_6_21_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03817 vss c_6_21_s1_s n4628 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03816 n4640 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03815 vss a_19 n4398 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03814 n4398 p_6_2_d2j n4642 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03813 n4642 p_6_2_d2jbar n4399 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03812 n4399 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03811 vss p_6_21_t_s p_6_21_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03810 p_6_21_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03809 n4642 n4640 p_6_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03808 p_6_21_t_s n4642 n4640 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03807 n5027 p_6_2_d2j n5026 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03806 n5025 p_6_2_d2jbar n5027 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03805 p_6_20_t_s n5027 n5024 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03804 n5027 n5024 p_6_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03803 p_6_20_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03802 vss p_6_20_t_s p_6_20_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03801 n5024 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03800 vss a_19 n5025 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03799 n5026 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03798 vss c_6_20_s1_s n5019 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03797 c_8_18_a c_6_20_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03796 c_6_20_s1_s p_6_20_pi2j c_6_20_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03795 c_6_20_s2_s n5019 c_5_21_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03794 n5019 c_5_21_cout c_6_20_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03793 vss p_6_20_pi2j n5015 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03792 n5015 c_6_20_a n5016 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03791 n5016 c_5_21_cout n5014 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03790 vss p_6_20_pi2j n5014 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03789 n5014 c_6_20_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03788 vss n5016 c_8_19_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03787 p_6_20_pi2j c_6_20_a c_6_20_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03786 vss n5392 c_6_19_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03785 n5138 p_6_19_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03784 vss c_6_19_a n5138 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03783 n5392 c_6_19_cin n5138 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03782 n5137 p_6_19_pi2j n5392 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03781 vss c_6_19_a n5137 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03780 n5388 c_6_19_cin c_6_19_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03779 c_6_19_s2_s n5388 c_6_19_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03778 c_6_19_a p_6_19_pi2j c_6_19_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03777 c_6_19_s1_s c_6_19_a p_6_19_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03776 c_8_17_a c_6_19_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03775 vss c_6_19_s1_s n5388 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03774 n5400 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03773 vss a_17 n5139 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03772 n5139 p_6_2_d2j n5402 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03771 n5402 p_6_2_d2jbar n5140 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03770 n5140 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03769 vss p_6_19_t_s p_6_19_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03768 p_6_19_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03767 n5402 n5400 p_6_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03766 p_6_19_t_s n5402 n5400 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03765 n5780 p_6_2_d2j n5778 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03764 n5779 p_6_2_d2jbar n5780 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03763 p_6_18_t_s n5780 n5777 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03762 n5780 n5777 p_6_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03761 p_6_18_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03760 vss p_6_18_t_s p_6_18_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03759 n5777 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03758 vss a_17 n5779 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03757 n5778 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03756 vss c_6_18_s1_s n5570 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03755 c_8_16_a c_6_18_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03754 c_6_18_s1_s p_6_18_pi2j c_6_18_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03753 c_6_18_s2_s n5570 c_5_19_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03752 n5570 c_5_19_cout c_6_18_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03751 vss p_6_18_pi2j n5770 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03750 n5770 c_6_18_a n5769 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03749 n5769 c_5_19_cout n5768 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03748 vss p_6_18_pi2j n5768 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03747 n5768 c_6_18_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03746 vss n5769 c_8_17_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03745 p_6_18_pi2j c_6_18_a c_6_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03744 vss n6185 c_6_17_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03743 n5907 p_6_17_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03742 vss c_6_17_a n5907 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03741 n6185 c_6_17_cin n5907 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03740 n5767 p_6_17_pi2j n6185 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03739 vss c_6_17_a n5767 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03738 n6178 c_6_17_cin c_6_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03737 c_6_17_s2_s n6178 c_6_17_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03736 c_6_17_a p_6_17_pi2j c_6_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03735 c_6_17_s1_s c_6_17_a p_6_17_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03734 c_8_15_a c_6_17_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03733 vss c_6_17_s1_s n6178 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03732 n6192 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03731 vss a_15 n5911 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03730 n5911 p_6_2_d2j n6187 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03729 n6187 p_6_2_d2jbar n5910 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03728 n5910 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03727 vss p_6_17_t_s p_6_17_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03726 p_6_17_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03725 n6187 n6192 p_6_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03724 p_6_17_t_s n6187 n6192 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03723 n6374 p_6_2_d2j n6373 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03722 n6375 p_6_2_d2jbar n6374 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03721 p_6_16_t_s n6374 n6559 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03720 n6374 n6559 p_6_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03719 p_6_16_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03718 vss p_6_16_t_s p_6_16_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03717 n6559 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03716 vss a_15 n6375 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03715 n6373 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03714 vss c_6_16_s1_s n6372 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03713 c_8_14_a c_6_16_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03712 c_6_16_s1_s p_6_16_pi2j c_6_16_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03711 c_6_16_s2_s n6372 c_5_17_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03710 n6372 c_5_17_cout c_6_16_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03709 vss p_6_16_pi2j n6553 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03708 n6553 c_6_16_a n6552 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03707 n6552 c_5_17_cout n6551 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03706 vss p_6_16_pi2j n6551 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03705 n6551 c_6_16_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03704 vss n6552 c_8_15_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03703 p_6_16_pi2j c_6_16_a c_6_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03702 vss n6969 c_6_15_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03701 n6550 c_6_15_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03700 vss c_6_15_a n6550 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03699 n6969 c_6_15_cin n6550 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03698 n6549 c_6_15_b n6969 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03697 vss c_6_15_a n6549 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03696 n6729 c_6_15_cin c_6_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03695 c_6_15_s2_s n6729 c_6_15_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03694 c_6_15_a c_6_15_b c_6_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03693 c_6_15_s1_s c_6_15_a c_6_15_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03692 c_8_13_a c_6_15_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03691 vss c_6_15_s1_s n6729 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03690 n6974 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03689 vss a_13 n6561 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03688 n6561 p_6_2_d2j n6735 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03687 n6735 p_6_2_d2jbar n6560 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03686 n6560 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03685 vss p_6_15_t_s c_6_15_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03684 c_6_15_b p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03683 n6735 n6974 p_6_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03682 p_6_15_t_s n6735 n6974 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03681 n7168 p_6_2_d2j n7169 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03680 n7170 p_6_2_d2jbar n7168 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03679 p_6_14_t_s n7168 n7167 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03678 n7168 n7167 p_6_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03677 p_6_14_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03676 vss p_6_14_t_s p_6_14_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03675 n7167 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03674 vss a_13 n7170 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03673 n7169 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03672 vss c_6_14_s1_s n7164 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03671 c_8_12_a c_6_14_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03670 c_6_14_s1_s p_6_14_pi2j c_6_14_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03669 c_6_14_s2_s n7164 c_5_15_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03668 n7164 c_5_15_cout c_6_14_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03667 vss p_6_14_pi2j n7325 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03666 n7325 c_6_14_a n7161 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03665 n7161 c_5_15_cout n7324 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03664 vss p_6_14_pi2j n7324 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03663 n7324 c_6_14_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03662 vss n7161 c_8_13_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03661 p_6_14_pi2j c_6_14_a c_6_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03660 vss n7526 c_6_13_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03659 n7323 c_6_13_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03658 vss c_6_13_a n7323 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03657 n7526 c_6_13_cin n7323 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03656 n7322 c_6_13_b n7526 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03655 vss c_6_13_a n7322 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03654 n7529 c_6_13_cin c_6_13_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03653 c_6_13_s2_s n7529 c_6_13_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03652 c_6_13_a c_6_13_b c_6_13_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03651 c_6_13_s1_s c_6_13_a c_6_13_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03650 c_8_11_a c_6_13_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03649 vss c_6_13_s1_s n7529 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03648 n7534 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03647 vss a_11 n7330 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03646 n7330 p_6_2_d2j n7536 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03645 n7536 p_6_2_d2jbar n7329 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03644 n7329 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03643 vss p_6_13_t_s c_6_13_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03642 c_6_13_b p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03641 n7536 n7534 p_6_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03640 p_6_13_t_s n7536 n7534 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03639 n7964 p_6_2_d2j n7962 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03638 n7963 p_6_2_d2jbar n7964 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03637 p_6_12_t_s n7964 n7961 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03636 n7964 n7961 p_6_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03635 c_6_12_b p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03634 vss p_6_12_t_s c_6_12_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03633 n7961 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03632 vss a_11 n7963 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03631 n7962 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03630 vss c_6_12_s1_s n7957 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03629 c_8_10_a c_6_12_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03628 c_6_12_s1_s c_6_12_b c_6_12_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03627 c_6_12_s2_s n7957 c_5_13_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03626 n7957 c_5_13_cout c_6_12_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03625 vss c_6_12_b n7953 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03624 n7953 c_6_12_a n7954 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03623 n7954 c_5_13_cout n7952 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03622 vss c_6_12_b n7952 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03621 n7952 c_6_12_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03620 vss n7954 c_8_11_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03619 c_6_12_b c_6_12_a c_6_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03618 vss n8321 c_6_11_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03617 n8083 p_6_11_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03616 vss c_6_11_a n8083 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03615 n8321 c_6_11_cin n8083 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03614 n8082 p_6_11_pi2j n8321 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03613 vss c_6_11_a n8082 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03612 n8316 c_6_11_cin c_6_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03611 c_6_11_s2_s n8316 c_6_11_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03610 c_6_11_a p_6_11_pi2j c_6_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03609 c_6_11_s1_s c_6_11_a p_6_11_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03608 c_8_9_a c_6_11_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03607 vss c_6_11_s1_s n8316 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03606 n8328 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03605 vss a_9 n8085 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03604 n8085 p_6_2_d2j n8330 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03603 n8330 p_6_2_d2jbar n8086 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03602 n8086 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03601 vss p_6_11_t_s p_6_11_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03600 p_6_11_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03599 n8330 n8328 p_6_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03598 p_6_11_t_s n8330 n8328 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03597 n8716 p_6_2_d2j n8715 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03596 n8714 p_6_2_d2jbar n8716 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03595 p_6_10_t_s n8716 n8713 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03594 n8716 n8713 p_6_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03593 p_6_10_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03592 vss p_6_10_t_s p_6_10_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03591 n8713 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03590 vss a_9 n8714 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03589 n8715 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03588 vss c_6_10_s1_s n8708 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03587 c_8_8_a c_6_10_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03586 c_6_10_s1_s p_6_10_pi2j c_6_10_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03585 c_6_10_s2_s n8708 c_5_11_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03584 n8708 c_5_11_cout c_6_10_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03583 vss p_6_10_pi2j n8705 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03582 n8705 c_6_10_a n8703 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03581 n8703 c_5_11_cout n8704 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03580 vss p_6_10_pi2j n8704 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03579 n8704 c_6_10_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03578 vss n8703 c_8_9_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03577 p_6_10_pi2j c_6_10_a c_6_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03576 vss n9080 c_6_9_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03575 n8830 p_6_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03574 vss c_6_9_a n8830 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_03573 n9080 c_6_9_cin n8830 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03572 n8829 p_6_9_pi2j n9080 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03571 vss c_6_9_a n8829 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_03570 n9076 c_6_9_cin c_6_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03569 c_6_9_s2_s n9076 c_6_9_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03568 c_6_9_a p_6_9_pi2j c_6_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03567 c_6_9_s1_s c_6_9_a p_6_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03566 c_8_7_a c_6_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03565 vss c_6_9_s1_s n9076 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03564 n9088 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03563 vss a_7 n8832 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03562 n8832 p_6_2_d2j n9090 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03561 n9090 p_6_2_d2jbar n8831 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03560 n8831 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03559 vss p_6_9_t_s p_6_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03558 p_6_9_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03557 n9090 n9088 p_6_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03556 p_6_9_t_s n9090 n9088 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03555 n9457 p_6_2_d2j n9458 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03554 n9456 p_6_2_d2jbar n9457 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03553 p_6_8_t_s n9457 n9455 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03552 n9457 n9455 p_6_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03551 p_6_8_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03550 vss p_6_8_t_s p_6_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03549 n9455 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03548 vss a_7 n9456 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03547 n9458 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03546 vss c_6_8_s1_s n9450 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03545 c_8_6_a c_6_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03544 c_6_8_s1_s p_6_8_pi2j c_6_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03543 c_6_8_s2_s n9450 c_5_9_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03542 n9450 c_5_9_cout c_6_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03541 vss p_6_8_pi2j n9446 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03540 n9446 c_6_8_a n9445 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03539 n9445 c_5_9_cout n9447 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03538 vss p_6_8_pi2j n9447 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03537 n9447 c_6_8_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_03536 vss n9445 c_8_7_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03535 p_6_8_pi2j c_6_8_a c_6_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03534 vss n9869 c_6_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03533 n9585 p_6_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03532 vss c_6_7_a n9585 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_03531 n9869 c_6_7_cin n9585 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03530 n9444 p_6_7_pi2j n9869 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03529 vss c_6_7_a n9444 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_03528 n9864 c_6_7_cin c_6_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03527 c_6_7_s2_s n9864 c_6_7_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03526 c_6_7_a p_6_7_pi2j c_6_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03525 c_6_7_s1_s c_6_7_a p_6_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03524 c_8_5_a c_6_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03523 vss c_6_7_s1_s n9864 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03522 n9876 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03521 vss a_5 n9588 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03520 n9588 p_6_2_d2j n9871 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03519 n9871 p_6_2_d2jbar n9589 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03518 n9589 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03517 vss p_6_7_t_s p_6_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03516 p_6_7_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03515 n9871 n9876 p_6_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03514 p_6_7_t_s n9871 n9876 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03513 n10230 p_6_2_d2j n10039 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03512 n10038 p_6_2_d2jbar n10230 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03511 p_6_6_t_s n10230 n10231 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03510 n10230 n10231 p_6_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03509 p_6_6_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03508 vss p_6_6_t_s p_6_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03507 n10231 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03506 vss a_5 n10038 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03505 n10039 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03504 vss c_6_6_s1_s n10037 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03503 c_8_4_a c_6_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03502 c_6_6_s1_s p_6_6_pi2j c_6_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03501 c_6_6_s2_s n10037 c_5_7_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03500 n10037 c_5_7_cout c_6_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03499 vss p_6_6_pi2j n10224 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03498 n10224 c_6_6_a n10223 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03497 n10223 c_5_7_cout n10222 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03496 vss p_6_6_pi2j n10222 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03495 n10222 c_6_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03494 vss n10223 c_8_5_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03493 p_6_6_pi2j c_6_6_a c_6_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03492 vss n10643 c_6_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03491 n10402 c_6_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03490 vss c_6_5_a n10402 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03489 n10643 c_6_5_cin n10402 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03488 n10221 c_6_5_b n10643 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03487 vss c_6_5_a n10221 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03486 n10404 c_6_5_cin c_6_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03485 c_6_5_s2_s n10404 c_6_5_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03484 c_6_5_a c_6_5_b c_6_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03483 c_6_5_s1_s c_6_5_a c_6_5_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03482 c_8_3_a c_6_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03481 vss c_6_5_s1_s n10404 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03480 n10651 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03479 vss a_3 n10233 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03478 n10233 p_6_2_d2j n10646 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03477 n10646 p_6_2_d2jbar n10232 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03476 n10232 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03475 vss p_6_5_t_s c_6_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03474 c_6_5_b p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03473 n10646 n10651 p_6_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03472 p_6_5_t_s n10646 n10651 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03471 n10844 p_6_2_d2j n10842 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03470 n10843 p_6_2_d2jbar n10844 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03469 p_6_4_t_s n10844 n10841 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03468 n10844 n10841 p_6_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03467 p_6_4_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03466 vss p_6_4_t_s p_6_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03465 n10841 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03464 vss a_3 n10843 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03463 n10842 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03462 vss c_6_4_s1_s n10838 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03461 c_8_2_a c_6_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03460 c_6_4_s1_s p_6_4_pi2j c_6_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03459 c_6_4_s2_s n10838 c_5_5_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03458 n10838 c_5_5_cout c_6_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03457 vss p_6_4_pi2j n10993 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03456 n10993 c_6_4_a n10835 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03455 n10835 c_5_5_cout n10992 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03454 vss p_6_4_pi2j n10992 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03453 n10992 c_6_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03452 vss n10835 c_8_3_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03451 p_6_4_pi2j c_6_4_a c_6_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03450 vss n11191 c_6_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03449 n10991 c_6_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03448 vss c_6_3_a n10991 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03447 n11191 c_6_3_cin n10991 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03446 n10990 c_6_3_b n11191 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03445 vss c_6_3_a n10990 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03444 n11193 c_6_3_cin c_6_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03443 c_6_3_s2_s n11193 c_6_3_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03442 c_6_3_a c_6_3_b c_6_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03441 c_6_3_s1_s c_6_3_a c_6_3_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03440 c_8_1_a c_6_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03439 vss c_6_3_s1_s n11193 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03438 n11199 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03437 vss a_1 n10998 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03436 n10998 p_6_2_d2j n11201 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03435 n11201 p_6_2_d2jbar n10997 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03434 n10997 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03433 vss p_6_3_t_s c_6_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03432 c_6_3_b p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03431 n11201 n11199 p_6_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03430 p_6_3_t_s n11201 n11199 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03429 n11627 p_6_2_d2j n11626 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03428 n11625 p_6_2_d2jbar n11627 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03427 p_6_2_t_s n11627 n11624 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03426 n11627 n11624 p_6_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03425 c_6_2_b p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03424 vss p_6_2_t_s c_6_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03423 n11624 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03422 vss a_1 n11625 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03421 n11626 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03420 vss c_6_2_s1_s n11620 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03419 c_6_2_sum c_6_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03418 c_6_2_s1_s c_6_2_b c_6_2_a vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03417 c_6_2_s2_s n11620 c_5_3_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03416 n11620 c_5_3_cout c_6_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03415 vss c_6_2_b n11616 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03414 n11616 c_6_2_a n11617 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03413 n11617 c_5_3_cout n11615 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03412 vss c_6_2_b n11615 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03411 n11615 c_6_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03410 vss n11617 c_8_1_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03409 c_6_2_b c_6_2_a c_6_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03408 vss n11985 c_6_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03407 n11745 p_6_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03406 vss c_6_1_a n11745 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03405 n11985 c_6_1_cin n11745 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03404 n11744 p_6_1_pi2j n11985 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03403 vss c_6_1_a n11744 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03402 n11981 c_6_1_cin c_6_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03401 c_6_1_s2_s n11981 c_6_1_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03400 c_6_1_a p_6_1_pi2j c_6_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03399 c_6_1_s1_s c_6_1_a p_6_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03398 c_6_1_sum c_6_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03397 vss c_6_1_s1_s n11981 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03396 n11995 p_6_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03395 n11997 p_6_2_d2jbar n11748 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03394 n11748 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03393 vss p_6_1_t_s p_6_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03392 p_6_1_pi2j p_6_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03391 n11997 n11995 p_6_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03390 p_6_1_t_s n11997 n11995 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03389 cl4_6_s1_s n12357 c_5_1_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03388 n12357 c_5_1_sum cl4_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03387 vss cl4_6_s1_s p_8 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03386 vss c_5_1_sum n12347 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03385 n12347 n12357 n12348 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03384 n12345 n12348 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_03383 n12346 c_5_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_03382 vss c_5_2_sum n12346 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_03381 n12343 c_5_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03380 n12342 c_5_1_cout n12343 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03379 n12341 c_5_1_sum n12342 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03378 n12346 n12357 n12341 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03377 n12339 n12342 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_03376 cl4_6_s2_s c_5_1_cout c_5_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03375 c_5_1_cout c_5_2_sum cl4_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03374 vss cl4_6_s2_s n12338 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03373 cl4_6_s3_s n12338 n12345 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03372 n12338 n12345 cl4_6_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03371 vss cl4_6_s3_s p_9 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03370 vss c_5_33_s1_s n205 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03369 c_6_31_a c_5_33_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03368 c_5_33_s1_s c_5_31_a p_5_33_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03367 c_5_31_a p_5_33_pi2j c_5_33_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03366 c_5_33_s2_s n205 c_5_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03365 n205 c_5_32_cin c_5_33_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03364 vss c_5_31_a n28 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_03363 n28 p_5_33_pi2j n204 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03362 n204 c_5_32_cin n27 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03361 vss c_5_31_a n27 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_03360 n27 p_5_33_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03359 vss n204 c_6_32_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03358 n213 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03357 n215 a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03356 vss p_5_33_t_s p_5_33_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03355 p_5_33_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03354 n215 n213 p_5_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03353 p_5_33_t_s n215 n213 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03352 n554 p_5_2_d2j n555 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03351 n553 p_5_2_d2jbar n554 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03350 p_5_32_t_s n554 n552 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03349 n554 n552 p_5_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03348 p_5_32_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03347 vss p_5_32_t_s p_5_32_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03346 n552 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03345 vss a_31 n553 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03344 n555 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03343 vss c_5_32_s1_s n549 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03342 c_6_30_a c_5_32_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03341 c_5_32_s1_s p_5_32_pi2j c_5_31_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03340 c_5_32_s2_s n549 c_5_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03339 n549 c_5_32_cin c_5_32_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03338 vss p_5_32_pi2j n543 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03337 n543 c_5_31_a n544 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03336 n544 c_5_32_cin n545 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03335 vss p_5_32_pi2j n545 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03334 n545 c_5_31_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_03333 vss n544 c_6_31_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03332 p_5_32_pi2j c_5_31_a c_5_32_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03331 vss n906 c_5_31_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03330 n650 p_5_31_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03329 vss c_5_31_a n650 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_03328 n906 c_5_31_cin n650 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03327 n649 p_5_31_pi2j n906 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03326 vss c_5_31_a n649 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_03325 n902 c_5_31_cin c_5_31_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03324 c_5_31_s2_s n902 c_5_31_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03323 c_5_31_a p_5_31_pi2j c_5_31_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03322 c_5_31_s1_s c_5_31_a p_5_31_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03321 c_6_29_a c_5_31_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03320 vss c_5_31_s1_s n902 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03319 n912 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03318 vss a_29 n651 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03317 n651 p_5_2_d2j n911 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03316 n911 p_5_2_d2jbar n652 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03315 n652 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03314 vss p_5_31_t_s p_5_31_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03313 p_5_31_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03312 n911 n912 p_5_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03311 p_5_31_t_s n911 n912 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03310 n1314 p_5_2_d2j n1316 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03309 n1315 p_5_2_d2jbar n1314 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03308 p_5_30_t_s n1314 n1312 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03307 n1314 n1312 p_5_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03306 p_5_30_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03305 vss p_5_30_t_s p_5_30_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03304 n1312 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03303 vss a_29 n1315 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03302 n1316 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03301 vss c_5_30_s1_s n1308 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03300 c_6_28_a c_5_30_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03299 c_5_30_s1_s p_5_30_pi2j c_5_30_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03298 c_5_30_s2_s n1308 c_4_31_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03297 n1308 c_4_31_cout c_5_30_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03296 vss p_5_30_pi2j n1304 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03295 n1304 c_5_30_a n1305 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03294 n1305 c_4_31_cout n1303 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03293 vss p_5_30_pi2j n1303 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03292 n1303 c_5_30_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03291 vss n1305 c_6_29_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03290 p_5_30_pi2j c_5_30_a c_5_30_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03289 vss n1687 c_5_29_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03288 n1412 p_5_29_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03287 vss c_5_29_a n1412 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03286 n1687 c_5_29_cin n1412 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03285 n1302 p_5_29_pi2j n1687 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03284 vss c_5_29_a n1302 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03283 n1684 c_5_29_cin c_5_29_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03282 c_5_29_s2_s n1684 c_5_29_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03281 c_5_29_a p_5_29_pi2j c_5_29_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03280 c_5_29_s1_s c_5_29_a p_5_29_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03279 c_6_27_a c_5_29_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03278 vss c_5_29_s1_s n1684 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03277 n1695 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03276 vss a_27 n1413 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03275 n1413 p_5_2_d2j n1693 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03274 n1693 p_5_2_d2jbar n1414 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03273 n1414 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03272 vss p_5_29_t_s p_5_29_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03271 p_5_29_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03270 n1693 n1695 p_5_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03269 p_5_29_t_s n1693 n1695 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03268 n2067 p_5_2_d2j n2068 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03267 n2066 p_5_2_d2jbar n2067 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03266 p_5_28_t_s n2067 n2065 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03265 n2067 n2065 p_5_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03264 p_5_28_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03263 vss p_5_28_t_s p_5_28_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03262 n2065 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03261 vss a_27 n2066 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03260 n2068 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03259 vss c_5_28_s1_s n1851 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03258 c_6_26_a c_5_28_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03257 c_5_28_s1_s p_5_28_pi2j c_5_28_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03256 c_5_28_s2_s n1851 c_4_29_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03255 n1851 c_4_29_cout c_5_28_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03254 vss p_5_28_pi2j n2058 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03253 n2058 c_5_28_a n2057 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03252 n2057 c_4_29_cout n2056 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03251 vss p_5_28_pi2j n2056 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03250 n2056 c_5_28_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03249 vss n2057 c_6_27_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03248 p_5_28_pi2j c_5_28_a c_5_28_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03247 vss n2498 c_5_27_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03246 n2211 c_5_27_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03245 vss c_5_27_a n2211 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03244 n2498 c_5_27_cin n2211 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03243 n2055 c_5_27_b n2498 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03242 vss c_5_27_a n2055 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03241 n2491 c_5_27_cin c_5_27_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03240 c_5_27_s2_s n2491 c_5_27_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03239 c_5_27_a c_5_27_b c_5_27_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03238 c_5_27_s1_s c_5_27_a c_5_27_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03237 c_6_25_a c_5_27_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03236 vss c_5_27_s1_s n2491 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03235 n2505 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03234 vss a_25 n2215 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03233 n2215 p_5_2_d2j n2501 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03232 n2501 p_5_2_d2jbar n2217 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03231 n2217 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03230 vss p_5_27_t_s c_5_27_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03229 c_5_27_b p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03228 n2501 n2505 p_5_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03227 p_5_27_t_s n2501 n2505 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03226 n2681 p_5_2_d2j n2683 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03225 n2682 p_5_2_d2jbar n2681 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03224 p_5_26_t_s n2681 n2680 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03223 n2681 n2680 p_5_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03222 p_5_26_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03221 vss p_5_26_t_s p_5_26_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03220 n2680 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03219 vss a_25 n2682 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03218 n2683 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03217 vss c_5_26_s1_s n2679 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03216 c_6_24_a c_5_26_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03215 c_5_26_s1_s p_5_26_pi2j c_5_26_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03214 c_5_26_s2_s n2679 c_4_27_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03213 n2679 c_4_27_cout c_5_26_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03212 vss p_5_26_pi2j n2869 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03211 n2869 c_5_26_a n2868 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03210 n2868 c_4_27_cout n2870 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03209 vss p_5_26_pi2j n2870 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03208 n2870 c_5_26_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03207 vss n2868 c_6_25_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03206 p_5_26_pi2j c_5_26_a c_5_26_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03205 vss n3284 c_5_25_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03204 n2867 c_5_25_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03203 vss c_5_25_a n2867 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03202 n3284 c_5_25_cin n2867 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03201 n2866 c_5_25_b n3284 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03200 vss c_5_25_a n2866 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03199 n3039 c_5_25_cin c_5_25_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03198 c_5_25_s2_s n3039 c_5_25_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03197 c_5_25_a c_5_25_b c_5_25_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03196 c_5_25_s1_s c_5_25_a c_5_25_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03195 c_6_23_a c_5_25_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03194 vss c_5_25_s1_s n3039 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03193 n3288 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03192 vss a_23 n2876 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03191 n2876 p_5_2_d2j n3042 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03190 n3042 p_5_2_d2jbar n2877 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03189 n2877 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03188 vss p_5_25_t_s c_5_25_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03187 c_5_25_b p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03186 n3042 n3288 p_5_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03185 p_5_25_t_s n3042 n3288 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03184 n3482 p_5_2_d2j n3484 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03183 n3483 p_5_2_d2jbar n3482 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03182 p_5_24_t_s n3482 n3481 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03181 n3482 n3481 p_5_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03180 c_5_24_b p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03179 vss p_5_24_t_s c_5_24_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03178 n3481 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03177 vss a_23 n3483 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03176 n3484 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03175 vss c_5_24_s1_s n3480 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03174 c_6_22_a c_5_24_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03173 c_5_24_s1_s c_5_24_b c_5_24_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03172 c_5_24_s2_s n3480 c_4_25_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03171 n3480 c_4_25_cout c_5_24_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03170 vss c_5_24_b n3626 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03169 n3626 c_5_24_a n3474 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03168 n3474 c_4_25_cout n3627 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03167 vss c_5_24_b n3627 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03166 n3627 c_5_24_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03165 vss n3474 c_6_23_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03164 c_5_24_b c_5_24_a c_5_24_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03163 vss n3873 c_5_23_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03162 n3625 c_5_23_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03161 vss c_5_23_a n3625 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03160 n3873 c_5_23_cin n3625 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03159 n3624 c_5_23_b n3873 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03158 vss c_5_23_a n3624 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03157 n3875 c_5_23_cin c_5_23_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03156 c_5_23_s2_s n3875 c_5_23_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03155 c_5_23_a c_5_23_b c_5_23_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03154 c_5_23_s1_s c_5_23_a c_5_23_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03153 c_6_21_a c_5_23_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03152 vss c_5_23_s1_s n3875 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03151 n3880 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03150 vss a_21 n3630 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03149 n3630 p_5_2_d2j n3879 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03148 n3879 p_5_2_d2jbar n3632 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03147 n3632 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03146 vss p_5_23_t_s c_5_23_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03145 c_5_23_b p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_03144 n3879 n3880 p_5_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03143 p_5_23_t_s n3879 n3880 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03142 n4293 p_5_2_d2j n4295 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03141 n4294 p_5_2_d2jbar n4293 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03140 p_5_22_t_s n4293 n4291 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03139 n4293 n4291 p_5_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03138 p_5_22_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03137 vss p_5_22_t_s p_5_22_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03136 n4291 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03135 vss a_21 n4294 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03134 n4295 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03133 vss c_5_22_s1_s n4289 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03132 c_6_20_a c_5_22_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03131 c_5_22_s1_s p_5_22_pi2j c_5_22_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03130 c_5_22_s2_s n4289 c_4_23_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03129 n4289 c_4_23_cout c_5_22_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03128 vss p_5_22_pi2j n4282 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03127 n4282 c_5_22_a n4283 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03126 n4283 c_4_23_cout n4284 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03125 vss p_5_22_pi2j n4284 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03124 n4284 c_5_22_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03123 vss n4283 c_6_21_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03122 p_5_22_pi2j c_5_22_a c_5_22_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03121 vss n4650 c_5_21_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03120 n4401 p_5_21_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03119 vss c_5_21_a n4401 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03118 n4650 c_5_21_cin n4401 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03117 n4400 p_5_21_pi2j n4650 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03116 vss c_5_21_a n4400 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03115 n4647 c_5_21_cin c_5_21_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03114 c_5_21_s2_s n4647 c_5_21_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03113 c_5_21_a p_5_21_pi2j c_5_21_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03112 c_5_21_s1_s c_5_21_a p_5_21_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03111 c_6_19_a c_5_21_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03110 vss c_5_21_s1_s n4647 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03109 n4659 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03108 vss a_19 n4402 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03107 n4402 p_5_2_d2j n4658 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03106 n4658 p_5_2_d2jbar n4403 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03105 n4403 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03104 vss p_5_21_t_s p_5_21_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03103 p_5_21_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03102 n4658 n4659 p_5_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03101 p_5_21_t_s n4658 n4659 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03100 n5039 p_5_2_d2j n5041 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03099 n5040 p_5_2_d2jbar n5039 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03098 p_5_20_t_s n5039 n5037 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03097 n5039 n5037 p_5_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03096 p_5_20_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03095 vss p_5_20_t_s p_5_20_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03094 n5037 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03093 vss a_19 n5040 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03092 n5041 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03091 vss c_5_20_s1_s n5035 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03090 c_6_18_a c_5_20_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03089 c_5_20_s1_s p_5_20_pi2j c_5_20_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03088 c_5_20_s2_s n5035 c_4_21_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03087 n5035 c_4_21_cout c_5_20_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03086 vss p_5_20_pi2j n5030 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03085 n5030 c_5_20_a n5029 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03084 n5029 c_4_21_cout n5028 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03083 vss p_5_20_pi2j n5028 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03082 n5028 c_5_20_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03081 vss n5029 c_6_19_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03080 p_5_20_pi2j c_5_20_a c_5_20_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03079 vss n5415 c_5_19_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03078 n5142 p_5_19_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03077 vss c_5_19_a n5142 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03076 n5415 c_5_19_cin n5142 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03075 n5141 p_5_19_pi2j n5415 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03074 vss c_5_19_a n5141 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03073 n5411 c_5_19_cin c_5_19_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03072 c_5_19_s2_s n5411 c_5_19_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03071 c_5_19_a p_5_19_pi2j c_5_19_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03070 c_5_19_s1_s c_5_19_a p_5_19_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03069 c_6_17_a c_5_19_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03068 vss c_5_19_s1_s n5411 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03067 n5422 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03066 vss a_17 n5143 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03065 n5143 p_5_2_d2j n5420 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03064 n5420 p_5_2_d2jbar n5144 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03063 n5144 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03062 vss p_5_19_t_s p_5_19_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03061 p_5_19_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03060 n5420 n5422 p_5_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03059 p_5_19_t_s n5420 n5422 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03058 n5791 p_5_2_d2j n5794 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03057 n5790 p_5_2_d2jbar n5791 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03056 p_5_18_t_s n5791 n5792 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03055 n5791 n5792 p_5_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03054 p_5_18_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03053 vss p_5_18_t_s p_5_18_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03052 n5792 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03051 vss a_17 n5790 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03050 n5794 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03049 vss c_5_18_s1_s n5577 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03048 c_6_16_a c_5_18_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03047 c_5_18_s1_s p_5_18_pi2j c_5_18_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03046 c_5_18_s2_s n5577 c_4_19_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03045 n5577 c_4_19_cout c_5_18_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03044 vss p_5_18_pi2j n5783 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03043 n5783 c_5_18_a n5782 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03042 n5782 c_4_19_cout n5784 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03041 vss p_5_18_pi2j n5784 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03040 n5784 c_5_18_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03039 vss n5782 c_6_17_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03038 p_5_18_pi2j c_5_18_a c_5_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03037 vss n6209 c_5_17_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_03036 n5912 p_5_17_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03035 vss c_5_17_a n5912 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03034 n6209 c_5_17_cin n5912 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03033 n5781 p_5_17_pi2j n6209 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03032 vss c_5_17_a n5781 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03031 n6199 c_5_17_cin c_5_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03030 c_5_17_s2_s n6199 c_5_17_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03029 c_5_17_a p_5_17_pi2j c_5_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03028 c_5_17_s1_s c_5_17_a p_5_17_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03027 c_6_15_a c_5_17_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03026 vss c_5_17_s1_s n6199 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03025 n6216 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03024 vss a_15 n5914 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03023 n5914 p_5_2_d2j n6210 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03022 n6210 p_5_2_d2jbar n5916 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03021 n5916 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03020 vss p_5_17_t_s p_5_17_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03019 p_5_17_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03018 n6210 n6216 p_5_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03017 p_5_17_t_s n6210 n6216 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03016 n6380 p_5_2_d2j n6382 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03015 n6381 p_5_2_d2jbar n6380 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_03014 p_5_16_t_s n6380 n6572 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03013 n6380 n6572 p_5_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03012 p_5_16_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03011 vss p_5_16_t_s p_5_16_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_03010 n6572 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_03009 vss a_15 n6381 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03008 n6382 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_03007 vss c_5_16_s1_s n6379 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_03006 c_6_14_a c_5_16_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_03005 c_5_16_s1_s p_5_16_pi2j c_5_16_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03004 c_5_16_s2_s n6379 c_4_17_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03003 n6379 c_4_17_cout c_5_16_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_03002 vss p_5_16_pi2j n6564 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03001 n6564 c_5_16_a n6565 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_03000 n6565 c_4_17_cout n6566 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02999 vss p_5_16_pi2j n6566 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02998 n6566 c_5_16_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02997 vss n6565 c_6_15_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02996 p_5_16_pi2j c_5_16_a c_5_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02995 vss n6987 c_5_15_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02994 n6563 c_5_15_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02993 vss c_5_15_a n6563 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02992 n6987 c_5_15_cin n6563 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02991 n6562 c_5_15_b n6987 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02990 vss c_5_15_a n6562 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02989 n6740 c_5_15_cin c_5_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02988 c_5_15_s2_s n6740 c_5_15_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02987 c_5_15_a c_5_15_b c_5_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02986 c_5_15_s1_s c_5_15_a c_5_15_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02985 c_6_13_a c_5_15_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02984 vss c_5_15_s1_s n6740 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02983 n6990 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02982 vss a_13 n6573 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02981 n6573 p_5_2_d2j n6743 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02980 n6743 p_5_2_d2jbar n6574 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02979 n6574 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02978 vss p_5_15_t_s c_5_15_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02977 c_5_15_b p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02976 n6743 n6990 p_5_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02975 p_5_15_t_s n6743 n6990 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02974 n7178 p_5_2_d2j n7180 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02973 n7179 p_5_2_d2jbar n7178 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02972 p_5_14_t_s n7178 n7177 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02971 n7178 n7177 p_5_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02970 p_5_14_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02969 vss p_5_14_t_s p_5_14_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02968 n7177 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02967 vss a_13 n7179 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02966 n7180 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02965 vss c_5_14_s1_s n7176 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02964 c_6_12_a c_5_14_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02963 c_5_14_s1_s p_5_14_pi2j c_5_14_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02962 c_5_14_s2_s n7176 c_4_15_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02961 n7176 c_4_15_cout c_5_14_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02960 vss p_5_14_pi2j n7333 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02959 n7333 c_5_14_a n7171 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02958 n7171 c_4_15_cout n7334 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02957 vss p_5_14_pi2j n7334 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02956 n7334 c_5_14_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02955 vss n7171 c_6_13_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02954 p_5_14_pi2j c_5_14_a c_5_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02953 vss n7542 c_5_13_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02952 n7332 c_5_13_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02951 vss c_5_13_a n7332 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02950 n7542 c_5_13_cin n7332 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02949 n7331 c_5_13_b n7542 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02948 vss c_5_13_a n7331 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02947 n7544 c_5_13_cin c_5_13_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02946 c_5_13_s2_s n7544 c_5_13_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02945 c_5_13_a c_5_13_b c_5_13_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02944 c_5_13_s1_s c_5_13_a c_5_13_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02943 c_6_11_a c_5_13_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02942 vss c_5_13_s1_s n7544 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02941 n7548 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02940 vss a_11 n7338 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02939 n7338 p_5_2_d2j n7547 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02938 n7547 p_5_2_d2jbar n7339 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02937 n7339 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02936 vss p_5_13_t_s c_5_13_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02935 c_5_13_b p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02934 n7547 n7548 p_5_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02933 p_5_13_t_s n7547 n7548 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02932 n7975 p_5_2_d2j n7977 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02931 n7976 p_5_2_d2jbar n7975 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02930 p_5_12_t_s n7975 n7973 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02929 n7975 n7973 p_5_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02928 c_5_12_b p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02927 vss p_5_12_t_s c_5_12_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02926 n7973 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02925 vss a_11 n7976 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02924 n7977 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02923 vss c_5_12_s1_s n7972 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02922 c_6_10_a c_5_12_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02921 c_5_12_s1_s c_5_12_b c_5_12_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02920 c_5_12_s2_s n7972 c_4_13_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02919 n7972 c_4_13_cout c_5_12_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02918 vss c_5_12_b n7965 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02917 n7965 c_5_12_a n7967 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02916 n7967 c_4_13_cout n7966 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02915 vss c_5_12_b n7966 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02914 n7966 c_5_12_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02913 vss n7967 c_6_11_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02912 c_5_12_b c_5_12_a c_5_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02911 vss n8340 c_5_11_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02910 n8088 p_5_11_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02909 vss c_5_11_a n8088 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02908 n8340 c_5_11_cin n8088 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02907 n8087 p_5_11_pi2j n8340 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02906 vss c_5_11_a n8087 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02905 n8335 c_5_11_cin c_5_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02904 c_5_11_s2_s n8335 c_5_11_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02903 c_5_11_a p_5_11_pi2j c_5_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02902 c_5_11_s1_s c_5_11_a p_5_11_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02901 c_6_9_a c_5_11_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02900 vss c_5_11_s1_s n8335 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02899 n8347 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02898 vss a_9 n8090 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02897 n8090 p_5_2_d2j n8346 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02896 n8346 p_5_2_d2jbar n8091 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02895 n8091 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02894 vss p_5_11_t_s p_5_11_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02893 p_5_11_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02892 n8346 n8347 p_5_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02891 p_5_11_t_s n8346 n8347 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02890 n8728 p_5_2_d2j n8730 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02889 n8729 p_5_2_d2jbar n8728 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02888 p_5_10_t_s n8728 n8726 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02887 n8728 n8726 p_5_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02886 p_5_10_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02885 vss p_5_10_t_s p_5_10_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02884 n8726 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02883 vss a_9 n8729 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02882 n8730 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02881 vss c_5_10_s1_s n8722 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02880 c_6_8_a c_5_10_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02879 c_5_10_s1_s p_5_10_pi2j c_5_10_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02878 c_5_10_s2_s n8722 c_4_11_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02877 n8722 c_4_11_cout c_5_10_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02876 vss p_5_10_pi2j n8719 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02875 n8719 c_5_10_a n8718 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02874 n8718 c_4_11_cout n8717 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02873 vss p_5_10_pi2j n8717 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02872 n8717 c_5_10_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02871 vss n8718 c_6_9_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02870 p_5_10_pi2j c_5_10_a c_5_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02869 vss n9103 c_5_9_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02868 n8834 p_5_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02867 vss c_5_9_a n8834 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02866 n9103 c_5_9_cin n8834 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02865 n8833 p_5_9_pi2j n9103 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02864 vss c_5_9_a n8833 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02863 n9099 c_5_9_cin c_5_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02862 c_5_9_s2_s n9099 c_5_9_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02861 c_5_9_a p_5_9_pi2j c_5_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02860 c_5_9_s1_s c_5_9_a p_5_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02859 c_6_7_a c_5_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02858 vss c_5_9_s1_s n9099 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02857 n9110 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02856 vss a_7 n8835 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02855 n8835 p_5_2_d2j n9108 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02854 n9108 p_5_2_d2jbar n8836 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02853 n8836 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02852 vss p_5_9_t_s p_5_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02851 p_5_9_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02850 n9108 n9110 p_5_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02849 p_5_9_t_s n9108 n9110 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02848 n9470 p_5_2_d2j n9473 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02847 n9469 p_5_2_d2jbar n9470 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02846 p_5_8_t_s n9470 n9471 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02845 n9470 n9471 p_5_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02844 p_5_8_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02843 vss p_5_8_t_s p_5_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02842 n9471 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02841 vss a_7 n9469 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02840 n9473 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02839 vss c_5_8_s1_s n9459 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02838 c_6_6_a c_5_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02837 c_5_8_s1_s p_5_8_pi2j c_5_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02836 c_5_8_s2_s n9459 c_4_9_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02835 n9459 c_4_9_cout c_5_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02834 vss p_5_8_pi2j n9462 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02833 n9462 c_5_8_a n9461 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02832 n9461 c_4_9_cout n9463 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02831 vss p_5_8_pi2j n9463 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02830 n9463 c_5_8_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02829 vss n9461 c_6_7_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02828 p_5_8_pi2j c_5_8_a c_5_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02827 vss n9892 c_5_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02826 n9590 p_5_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02825 vss c_5_7_a n9590 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02824 n9892 c_5_7_cin n9590 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02823 n9460 p_5_7_pi2j n9892 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02822 vss c_5_7_a n9460 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02821 n9887 c_5_7_cin c_5_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02820 c_5_7_s2_s n9887 c_5_7_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02819 c_5_7_a p_5_7_pi2j c_5_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02818 c_5_7_s1_s c_5_7_a p_5_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02817 c_6_5_a c_5_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02816 vss c_5_7_s1_s n9887 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02815 n9900 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02814 vss a_5 n9592 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02813 n9592 p_5_2_d2j n9894 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02812 n9894 p_5_2_d2jbar n9594 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02811 n9594 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02810 vss p_5_7_t_s p_5_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02809 p_5_7_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02808 n9894 n9900 p_5_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02807 p_5_7_t_s n9894 n9900 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02806 n10244 p_5_2_d2j n10044 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02805 n10043 p_5_2_d2jbar n10244 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02804 p_5_6_t_s n10244 n10245 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02803 n10244 n10245 p_5_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02802 p_5_6_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02801 vss p_5_6_t_s p_5_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02800 n10245 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02799 vss a_5 n10043 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02798 n10044 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02797 vss c_5_6_s1_s n10042 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02796 c_6_4_a c_5_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02795 c_5_6_s1_s p_5_6_pi2j c_5_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02794 c_5_6_s2_s n10042 c_4_7_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02793 n10042 c_4_7_cout c_5_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02792 vss p_5_6_pi2j n10236 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02791 n10236 c_5_6_a n10237 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02790 n10237 c_4_7_cout n10238 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02789 vss p_5_6_pi2j n10238 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02788 n10238 c_5_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02787 vss n10237 c_6_5_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02786 p_5_6_pi2j c_5_6_a c_5_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02785 vss n10662 c_5_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02784 n10411 c_5_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02783 vss c_5_5_a n10411 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02782 n10662 c_5_5_cin n10411 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02781 n10235 c_5_5_b n10662 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02780 vss c_5_5_a n10235 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02779 n10415 c_5_5_cin c_5_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02778 c_5_5_s2_s n10415 c_5_5_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02777 c_5_5_a c_5_5_b c_5_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02776 c_5_5_s1_s c_5_5_a c_5_5_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02775 c_6_3_a c_5_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02774 vss c_5_5_s1_s n10415 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02773 n10668 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02772 vss a_3 n10246 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02771 n10246 p_5_2_d2j n10665 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02770 n10665 p_5_2_d2jbar n10247 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02769 n10247 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02768 vss p_5_5_t_s c_5_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02767 c_5_5_b p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02766 n10665 n10668 p_5_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02765 p_5_5_t_s n10665 n10668 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02764 n10852 p_5_2_d2j n10854 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02763 n10853 p_5_2_d2jbar n10852 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02762 p_5_4_t_s n10852 n10851 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02761 n10852 n10851 p_5_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02760 p_5_4_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02759 vss p_5_4_t_s p_5_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02758 n10851 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02757 vss a_3 n10853 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02756 n10854 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02755 vss c_5_4_s1_s n10850 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02754 c_6_2_a c_5_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02753 c_5_4_s1_s p_5_4_pi2j c_5_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02752 c_5_4_s2_s n10850 c_4_5_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02751 n10850 c_4_5_cout c_5_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02750 vss p_5_4_pi2j n11001 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02749 n11001 c_5_4_a n10845 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02748 n10845 c_4_5_cout n11002 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02747 vss p_5_4_pi2j n11002 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02746 n11002 c_5_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02745 vss n10845 c_6_3_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02744 p_5_4_pi2j c_5_4_a c_5_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02743 vss n11207 c_5_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02742 n11000 c_5_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02741 vss c_5_3_a n11000 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02740 n11207 c_5_3_cin n11000 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02739 n10999 c_5_3_b n11207 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02738 vss c_5_3_a n10999 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02737 n11209 c_5_3_cin c_5_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02736 c_5_3_s2_s n11209 c_5_3_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02735 c_5_3_a c_5_3_b c_5_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02734 c_5_3_s1_s c_5_3_a c_5_3_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02733 c_6_1_a c_5_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02732 vss c_5_3_s1_s n11209 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02731 n11213 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02730 vss a_1 n11006 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02729 n11006 p_5_2_d2j n11212 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02728 n11212 p_5_2_d2jbar n11007 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02727 n11007 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02726 vss p_5_3_t_s c_5_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02725 c_5_3_b p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02724 n11212 n11213 p_5_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02723 p_5_3_t_s n11212 n11213 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02722 n11638 p_5_2_d2j n11640 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02721 n11639 p_5_2_d2jbar n11638 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02720 p_5_2_t_s n11638 n11636 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02719 n11638 n11636 p_5_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02718 c_5_2_b p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02717 vss p_5_2_t_s c_5_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02716 n11636 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02715 vss a_1 n11639 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02714 n11640 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02713 vss c_5_2_s1_s n11635 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02712 c_5_2_sum c_5_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02711 c_5_2_s1_s c_5_2_b c_5_2_a vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02710 c_5_2_s2_s n11635 c_4_3_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02709 n11635 c_4_3_cout c_5_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02708 vss c_5_2_b n11628 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02707 n11628 c_5_2_a n11629 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02706 n11629 c_4_3_cout n11630 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02705 vss c_5_2_b n11630 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02704 n11630 c_5_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02703 vss n11629 c_6_1_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02702 c_5_2_b c_5_2_a c_5_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02701 vss n12004 c_5_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02700 n11750 p_5_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02699 vss c_5_1_a n11750 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02698 n12004 c_5_1_cin n11750 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02697 n11749 p_5_1_pi2j n12004 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02696 vss c_5_1_a n11749 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02695 n12001 c_5_1_cin c_5_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02694 c_5_1_s2_s n12001 c_5_1_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02693 c_5_1_a p_5_1_pi2j c_5_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02692 c_5_1_s1_s c_5_1_a p_5_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02691 c_5_1_sum c_5_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02690 vss c_5_1_s1_s n12001 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02689 n12015 p_5_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02688 n12014 p_5_2_d2jbar n11753 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02687 n11753 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02686 vss p_5_1_t_s p_5_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02685 p_5_1_pi2j p_5_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02684 n12014 n12015 p_5_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02683 p_5_1_t_s n12014 n12015 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02682 cl4_5_s1_s n12375 c_4_1_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02681 n12375 c_4_1_sum cl4_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02680 vss cl4_5_s1_s p_6 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02679 vss c_4_1_sum n12365 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02678 n12365 n12375 n12364 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02677 n12363 n12364 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02676 n12362 c_4_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_02675 vss c_4_2_sum n12362 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_02674 n12359 c_4_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02673 n12361 c_4_1_cout n12359 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02672 n12360 c_4_1_sum n12361 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02671 n12362 n12375 n12360 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02670 n12357 n12361 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02669 cl4_5_s2_s c_4_1_cout c_4_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02668 c_4_1_cout c_4_2_sum cl4_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02667 vss cl4_5_s2_s n12356 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02666 cl4_5_s3_s n12356 n12363 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02665 n12356 n12363 cl4_5_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02664 vss cl4_5_s3_s p_7 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02663 vss c_4_33_s1_s n223 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02662 c_5_31_a c_4_33_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02661 c_4_33_s1_s c_4_31_a p_4_33_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02660 c_4_31_a p_4_33_pi2j c_4_33_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02659 c_4_33_s2_s n223 c_4_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02658 n223 c_4_32_cin c_4_33_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02657 vss c_4_31_a n29 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02656 n29 p_4_33_pi2j n220 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02655 n220 c_4_32_cin n30 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02654 vss c_4_31_a n30 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02653 n30 p_4_33_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02652 vss n220 c_5_32_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02651 n228 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02650 n229 a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02649 vss p_4_33_t_s p_4_33_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02648 p_4_33_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02647 n229 n228 p_4_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02646 p_4_33_t_s n229 n228 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02645 n568 p_4_2_d2j n566 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02644 n567 p_4_2_d2jbar n568 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02643 p_4_32_t_s n568 n565 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02642 n568 n565 p_4_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02641 p_4_32_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02640 vss p_4_32_t_s p_4_32_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02639 n565 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02638 vss a_31 n567 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02637 n566 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02636 vss c_4_32_s1_s n561 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02635 c_5_30_a c_4_32_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02634 c_4_32_s1_s p_4_32_pi2j c_4_31_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02633 c_4_32_s2_s n561 c_4_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02632 n561 c_4_32_cin c_4_32_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02631 vss p_4_32_pi2j n557 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02630 n557 c_4_31_a n558 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02629 n558 c_4_32_cin n556 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02628 vss p_4_32_pi2j n556 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02627 n556 c_4_31_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02626 vss n558 c_5_31_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02625 p_4_32_pi2j c_4_31_a c_4_32_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02624 vss n925 c_4_31_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02623 n654 p_4_31_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02622 vss c_4_31_a n654 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02621 n925 c_4_31_cin n654 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02620 n653 p_4_31_pi2j n925 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02619 vss c_4_31_a n653 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02618 n922 c_4_31_cin c_4_31_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02617 c_4_31_s2_s n922 c_4_31_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02616 c_4_31_a p_4_31_pi2j c_4_31_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02615 c_4_31_s1_s c_4_31_a p_4_31_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02614 c_5_29_a c_4_31_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02613 vss c_4_31_s1_s n922 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02612 n932 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02611 vss a_29 n656 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02610 n656 p_4_2_d2j n929 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02609 n929 p_4_2_d2jbar n655 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02608 n655 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02607 vss p_4_31_t_s p_4_31_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02606 p_4_31_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02605 n929 n932 p_4_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02604 p_4_31_t_s n929 n932 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02603 n1331 p_4_2_d2j n1329 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02602 n1330 p_4_2_d2jbar n1331 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02601 p_4_30_t_s n1331 n1328 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02600 n1331 n1328 p_4_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02599 p_4_30_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02598 vss p_4_30_t_s p_4_30_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02597 n1328 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02596 vss a_29 n1330 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02595 n1329 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02594 vss c_4_30_s1_s n1325 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02593 c_5_28_a c_4_30_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02592 c_4_30_s1_s p_4_30_pi2j c_4_30_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02591 c_4_30_s2_s n1325 c_3_31_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02590 n1325 c_3_31_cout c_4_30_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02589 vss p_4_30_pi2j n1319 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02588 n1319 c_4_30_a n1318 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02587 n1318 c_3_31_cout n1320 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02586 vss p_4_30_pi2j n1320 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02585 n1320 c_4_30_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02584 vss n1318 c_5_29_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02583 p_4_30_pi2j c_4_30_a c_4_30_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02582 vss n1709 c_4_29_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02581 n1415 p_4_29_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02580 vss c_4_29_a n1415 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02579 n1709 c_4_29_cin n1415 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02578 n1317 p_4_29_pi2j n1709 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02577 vss c_4_29_a n1317 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02576 n1704 c_4_29_cin c_4_29_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02575 c_4_29_s2_s n1704 c_4_29_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02574 c_4_29_a p_4_29_pi2j c_4_29_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02573 c_4_29_s1_s c_4_29_a p_4_29_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02572 c_5_27_a c_4_29_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02571 vss c_4_29_s1_s n1704 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02570 n1716 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02569 vss a_27 n1417 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02568 n1417 p_4_2_d2j n1714 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02567 n1714 p_4_2_d2jbar n1416 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02566 n1416 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02565 vss p_4_29_t_s p_4_29_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02564 p_4_29_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02563 n1714 n1716 p_4_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02562 p_4_29_t_s n1714 n1716 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02561 n2081 p_4_2_d2j n2079 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02560 n2080 p_4_2_d2jbar n2081 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02559 p_4_28_t_s n2081 n2082 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02558 n2081 n2082 p_4_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02557 p_4_28_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02556 vss p_4_28_t_s p_4_28_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02555 n2082 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02554 vss a_27 n2080 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02553 n2079 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02552 vss c_4_28_s1_s n1859 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02551 c_5_26_a c_4_28_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02550 c_4_28_s1_s p_4_28_pi2j c_4_28_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02549 c_4_28_s2_s n1859 c_3_29_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02548 n1859 c_3_29_cout c_4_28_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02547 vss p_4_28_pi2j n2073 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02546 n2073 c_4_28_a n2071 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02545 n2071 c_3_29_cout n2072 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02544 vss p_4_28_pi2j n2072 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02543 n2072 c_4_28_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02542 vss n2071 c_5_27_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02541 p_4_28_pi2j c_4_28_a c_4_28_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02540 vss n2521 c_4_27_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02539 n2218 c_4_27_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02538 vss c_4_27_a n2218 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02537 n2521 c_4_27_cin n2218 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02536 n2070 c_4_27_b n2521 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02535 vss c_4_27_a n2070 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02534 n2511 c_4_27_cin c_4_27_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02533 c_4_27_s2_s n2511 c_4_27_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02532 c_4_27_a c_4_27_b c_4_27_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02531 c_4_27_s1_s c_4_27_a c_4_27_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02530 c_5_25_a c_4_27_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02529 vss c_4_27_s1_s n2511 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02528 n2526 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02527 vss a_25 n2223 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02526 n2223 p_4_2_d2j n2522 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02525 n2522 p_4_2_d2jbar n2224 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02524 n2224 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02523 vss p_4_27_t_s c_4_27_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02522 c_4_27_b p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02521 n2522 n2526 p_4_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02520 p_4_27_t_s n2522 n2526 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02519 n2691 p_4_2_d2j n2689 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02518 n2690 p_4_2_d2jbar n2691 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02517 p_4_26_t_s n2691 n2688 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02516 n2691 n2688 p_4_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02515 p_4_26_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02514 vss p_4_26_t_s p_4_26_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02513 n2688 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02512 vss a_25 n2690 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02511 n2689 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02510 vss c_4_26_s1_s n2687 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02509 c_5_24_a c_4_26_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02508 c_4_26_s1_s p_4_26_pi2j c_4_26_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02507 c_4_26_s2_s n2687 c_3_27_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02506 n2687 c_3_27_cout c_4_26_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02505 vss p_4_26_pi2j n2882 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02504 n2882 c_4_26_a n2883 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02503 n2883 c_3_27_cout n2878 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02502 vss p_4_26_pi2j n2878 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02501 n2878 c_4_26_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02500 vss n2883 c_5_25_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02499 p_4_26_pi2j c_4_26_a c_4_26_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02498 vss n3302 c_4_25_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02497 n2881 c_4_25_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02496 vss c_4_25_a n2881 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02495 n3302 c_4_25_cin n2881 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02494 n2880 c_4_25_b n3302 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02493 vss c_4_25_a n2880 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02492 n3049 c_4_25_cin c_4_25_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02491 c_4_25_s2_s n3049 c_4_25_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02490 c_4_25_a c_4_25_b c_4_25_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02489 c_4_25_s1_s c_4_25_a c_4_25_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02488 c_5_23_a c_4_25_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02487 vss c_4_25_s1_s n3049 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02486 n3305 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02485 vss a_23 n2889 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02484 n2889 p_4_2_d2j n3051 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02483 n3051 p_4_2_d2jbar n2888 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02482 n2888 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02481 vss p_4_25_t_s c_4_25_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02480 c_4_25_b p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02479 n3051 n3305 p_4_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02478 p_4_25_t_s n3051 n3305 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02477 n3495 p_4_2_d2j n3493 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02476 n3494 p_4_2_d2jbar n3495 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02475 p_4_24_t_s n3495 n3492 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02474 n3495 n3492 p_4_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02473 c_4_24_b p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02472 vss p_4_24_t_s c_4_24_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02471 n3492 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02470 vss a_23 n3494 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02469 n3493 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02468 vss c_4_24_s1_s n3489 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02467 c_5_22_a c_4_24_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02466 c_4_24_s1_s c_4_24_b c_4_24_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02465 c_4_24_s2_s n3489 c_3_25_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02464 n3489 c_3_25_cout c_4_24_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02463 vss c_4_24_b n3635 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02462 n3635 c_4_24_a n3485 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02461 n3485 c_3_25_cout n3631 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02460 vss c_4_24_b n3631 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02459 n3631 c_4_24_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02458 vss n3485 c_5_23_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02457 c_4_24_b c_4_24_a c_4_24_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02456 vss n3891 c_4_23_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02455 n3634 c_4_23_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02454 vss c_4_23_a n3634 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02453 n3891 c_4_23_cin n3634 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02452 n3633 c_4_23_b n3891 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02451 vss c_4_23_a n3633 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02450 n3892 c_4_23_cin c_4_23_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02449 c_4_23_s2_s n3892 c_4_23_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02448 c_4_23_a c_4_23_b c_4_23_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02447 c_4_23_s1_s c_4_23_a c_4_23_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02446 c_5_21_a c_4_23_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02445 vss c_4_23_s1_s n3892 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02444 n3898 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02443 vss a_21 n3639 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02442 n3639 p_4_2_d2j n3895 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02441 n3895 p_4_2_d2jbar n3638 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02440 n3638 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02439 vss p_4_23_t_s c_4_23_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02438 c_4_23_b p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02437 n3895 n3898 p_4_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02436 p_4_23_t_s n3895 n3898 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02435 n4309 p_4_2_d2j n4307 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02434 n4308 p_4_2_d2jbar n4309 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02433 p_4_22_t_s n4309 n4306 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02432 n4309 n4306 p_4_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02431 p_4_22_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02430 vss p_4_22_t_s p_4_22_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02429 n4306 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02428 vss a_21 n4308 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02427 n4307 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02426 vss c_4_22_s1_s n4301 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02425 c_5_20_a c_4_22_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02424 c_4_22_s1_s p_4_22_pi2j c_4_22_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02423 c_4_22_s2_s n4301 c_3_23_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02422 n4301 c_3_23_cout c_4_22_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02421 vss p_4_22_pi2j n4297 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02420 n4297 c_4_22_a n4298 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02419 n4298 c_3_23_cout n4296 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02418 vss p_4_22_pi2j n4296 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02417 n4296 c_4_22_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02416 vss n4298 c_5_21_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02415 p_4_22_pi2j c_4_22_a c_4_22_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02414 vss n4671 c_4_21_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02413 n4405 p_4_21_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02412 vss c_4_21_a n4405 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02411 n4671 c_4_21_cin n4405 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02410 n4404 p_4_21_pi2j n4671 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02409 vss c_4_21_a n4404 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02408 n4667 c_4_21_cin c_4_21_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02407 c_4_21_s2_s n4667 c_4_21_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02406 c_4_21_a p_4_21_pi2j c_4_21_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02405 c_4_21_s1_s c_4_21_a p_4_21_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02404 c_5_19_a c_4_21_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02403 vss c_4_21_s1_s n4667 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02402 n4679 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02401 vss a_19 n4407 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02400 n4407 p_4_2_d2j n4676 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02399 n4676 p_4_2_d2jbar n4406 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02398 n4406 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02397 vss p_4_21_t_s p_4_21_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02396 p_4_21_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02395 n4676 n4679 p_4_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02394 p_4_21_t_s n4676 n4679 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02393 n5055 p_4_2_d2j n5053 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02392 n5054 p_4_2_d2jbar n5055 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02391 p_4_20_t_s n5055 n5052 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02390 n5055 n5052 p_4_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02389 p_4_20_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02388 vss p_4_20_t_s p_4_20_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02387 n5052 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02386 vss a_19 n5054 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02385 n5053 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02384 vss c_4_20_s1_s n5048 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02383 c_5_18_a c_4_20_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02382 c_4_20_s1_s p_4_20_pi2j c_4_20_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02381 c_4_20_s2_s n5048 c_3_21_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02380 n5048 c_3_21_cout c_4_20_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02379 vss p_4_20_pi2j n5043 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02378 n5043 c_4_20_a n5042 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02377 n5042 c_3_21_cout n5044 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02376 vss p_4_20_pi2j n5044 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02375 n5044 c_4_20_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02374 vss n5042 c_5_19_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02373 p_4_20_pi2j c_4_20_a c_4_20_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02372 vss n5436 c_4_19_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02371 n5145 p_4_19_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02370 vss c_4_19_a n5145 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02369 n5436 c_4_19_cin n5145 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02368 n5146 p_4_19_pi2j n5436 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02367 vss c_4_19_a n5146 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02366 n5431 c_4_19_cin c_4_19_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02365 c_4_19_s2_s n5431 c_4_19_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02364 c_4_19_a p_4_19_pi2j c_4_19_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02363 c_4_19_s1_s c_4_19_a p_4_19_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02362 c_5_17_a c_4_19_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02361 vss c_4_19_s1_s n5431 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02360 n5443 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02359 vss a_17 n5148 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02358 n5148 p_4_2_d2j n5441 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02357 n5441 p_4_2_d2jbar n5147 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02356 n5147 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02355 vss p_4_19_t_s p_4_19_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02354 p_4_19_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02353 n5441 n5443 p_4_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02352 p_4_19_t_s n5441 n5443 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02351 n5808 p_4_2_d2j n5807 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02350 n5805 p_4_2_d2jbar n5808 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02349 p_4_18_t_s n5808 n5806 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02348 n5808 n5806 p_4_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02347 p_4_18_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02346 vss p_4_18_t_s p_4_18_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02345 n5806 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02344 vss a_17 n5805 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02343 n5807 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02342 vss c_4_18_s1_s n5585 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02341 c_5_16_a c_4_18_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02340 c_4_18_s1_s p_4_18_pi2j c_4_18_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02339 c_4_18_s2_s n5585 c_3_19_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02338 n5585 c_3_19_cout c_4_18_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02337 vss p_4_18_pi2j n5797 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02336 n5797 c_4_18_a n5799 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02335 n5799 c_3_19_cout n5798 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02334 vss p_4_18_pi2j n5798 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02333 n5798 c_4_18_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02332 vss n5799 c_5_17_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02331 p_4_18_pi2j c_4_18_a c_4_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02330 vss n6233 c_4_17_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02329 n5917 p_4_17_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02328 vss c_4_17_a n5917 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02327 n6233 c_4_17_cin n5917 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02326 n5796 p_4_17_pi2j n6233 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02325 vss c_4_17_a n5796 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02324 n6222 c_4_17_cin c_4_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02323 c_4_17_s2_s n6222 c_4_17_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02322 c_4_17_a p_4_17_pi2j c_4_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02321 c_4_17_s1_s c_4_17_a p_4_17_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02320 c_5_15_a c_4_17_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02319 vss c_4_17_s1_s n6222 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02318 n6239 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02317 vss a_15 n5920 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02316 n5920 p_4_2_d2j n6234 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02315 n6234 p_4_2_d2jbar n5921 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02314 n5921 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02313 vss p_4_17_t_s p_4_17_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02312 p_4_17_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02311 n6234 n6239 p_4_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02310 p_4_17_t_s n6234 n6239 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02309 n6389 p_4_2_d2j n6387 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02308 n6388 p_4_2_d2jbar n6389 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02307 p_4_16_t_s n6389 n6585 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02306 n6389 n6585 p_4_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02305 p_4_16_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02304 vss p_4_16_t_s p_4_16_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02303 n6585 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02302 vss a_15 n6388 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02301 n6387 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02300 vss c_4_16_s1_s n6386 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02299 c_5_14_a c_4_16_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02298 c_4_16_s1_s p_4_16_pi2j c_4_16_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02297 c_4_16_s2_s n6386 c_3_17_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02296 n6386 c_3_17_cout c_4_16_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02295 vss p_4_16_pi2j n6579 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02294 n6579 c_4_16_a n6580 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02293 n6580 c_3_17_cout n6575 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02292 vss p_4_16_pi2j n6575 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02291 n6575 c_4_16_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02290 vss n6580 c_5_15_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02289 p_4_16_pi2j c_4_16_a c_4_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02288 vss n7003 c_4_15_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02287 n6578 c_4_15_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02286 vss c_4_15_a n6578 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02285 n7003 c_4_15_cin n6578 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02284 n6577 c_4_15_b n7003 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02283 vss c_4_15_a n6577 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02282 n6750 c_4_15_cin c_4_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02281 c_4_15_s2_s n6750 c_4_15_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02280 c_4_15_a c_4_15_b c_4_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02279 c_4_15_s1_s c_4_15_a c_4_15_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02278 c_5_13_a c_4_15_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02277 vss c_4_15_s1_s n6750 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02276 n7007 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02275 vss a_13 n6587 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02274 n6587 p_4_2_d2j n6752 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02273 n6752 p_4_2_d2jbar n6586 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02272 n6586 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02271 vss p_4_15_t_s c_4_15_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02270 c_4_15_b p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02269 n6752 n7007 p_4_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02268 p_4_15_t_s n6752 n7007 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02267 n7190 p_4_2_d2j n7188 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02266 n7189 p_4_2_d2jbar n7190 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02265 p_4_14_t_s n7190 n7187 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02264 n7190 n7187 p_4_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02263 p_4_14_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02262 vss p_4_14_t_s p_4_14_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02261 n7187 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02260 vss a_13 n7189 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02259 n7188 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02258 vss c_4_14_s1_s n7184 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02257 c_5_12_a c_4_14_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02256 c_4_14_s1_s p_4_14_pi2j c_4_14_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02255 c_4_14_s2_s n7184 c_3_15_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02254 n7184 c_3_15_cout c_4_14_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02253 vss p_4_14_pi2j n7344 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02252 n7344 c_4_14_a n7181 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02251 n7181 c_3_15_cout n7340 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02250 vss p_4_14_pi2j n7340 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02249 n7340 c_4_14_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02248 vss n7181 c_5_13_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02247 p_4_14_pi2j c_4_14_a c_4_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02246 vss n7556 c_4_13_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02245 n7343 c_4_13_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02244 vss c_4_13_a n7343 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02243 n7556 c_4_13_cin n7343 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02242 n7342 c_4_13_b n7556 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02241 vss c_4_13_a n7342 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02240 n7558 c_4_13_cin c_4_13_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02239 c_4_13_s2_s n7558 c_4_13_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02238 c_4_13_a c_4_13_b c_4_13_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02237 c_4_13_s1_s c_4_13_a c_4_13_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02236 c_5_11_a c_4_13_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02235 vss c_4_13_s1_s n7558 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02234 n7563 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02233 vss a_11 n7348 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02232 n7348 p_4_2_d2j n7560 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02231 n7560 p_4_2_d2jbar n7347 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02230 n7347 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02229 vss p_4_13_t_s c_4_13_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02228 c_4_13_b p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02227 n7560 n7563 p_4_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02226 p_4_13_t_s n7560 n7563 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02225 n7990 p_4_2_d2j n7988 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02224 n7989 p_4_2_d2jbar n7990 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02223 p_4_12_t_s n7990 n7987 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02222 n7990 n7987 p_4_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02221 c_4_12_b p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02220 vss p_4_12_t_s c_4_12_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02219 n7987 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02218 vss a_11 n7989 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02217 n7988 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02216 vss c_4_12_s1_s n7983 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02215 c_5_10_a c_4_12_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02214 c_4_12_s1_s c_4_12_b c_4_12_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02213 c_4_12_s2_s n7983 c_3_13_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02212 n7983 c_3_13_cout c_4_12_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02211 vss c_4_12_b n7980 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02210 n7980 c_4_12_a n7978 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02209 n7978 c_3_13_cout n7979 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02208 vss c_4_12_b n7979 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02207 n7979 c_4_12_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02206 vss n7978 c_5_11_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02205 c_4_12_b c_4_12_a c_4_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02204 vss n8360 c_4_11_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02203 n8093 p_4_11_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02202 vss c_4_11_a n8093 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02201 n8360 c_4_11_cin n8093 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02200 n8092 p_4_11_pi2j n8360 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02199 vss c_4_11_a n8092 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02198 n8355 c_4_11_cin c_4_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02197 c_4_11_s2_s n8355 c_4_11_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02196 c_4_11_a p_4_11_pi2j c_4_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02195 c_4_11_s1_s c_4_11_a p_4_11_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02194 c_5_9_a c_4_11_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02193 vss c_4_11_s1_s n8355 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02192 n8367 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02191 vss a_9 n8096 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02190 n8096 p_4_2_d2j n8364 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02189 n8364 p_4_2_d2jbar n8095 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02188 n8095 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02187 vss p_4_11_t_s p_4_11_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02186 p_4_11_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02185 n8364 n8367 p_4_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02184 p_4_11_t_s n8364 n8367 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02183 n8744 p_4_2_d2j n8742 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02182 n8743 p_4_2_d2jbar n8744 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02181 p_4_10_t_s n8744 n8741 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02180 n8744 n8741 p_4_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02179 p_4_10_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02178 vss p_4_10_t_s p_4_10_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02177 n8741 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02176 vss a_9 n8743 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02175 n8742 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02174 vss c_4_10_s1_s n8738 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02173 c_5_8_a c_4_10_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02172 c_4_10_s1_s p_4_10_pi2j c_4_10_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02171 c_4_10_s2_s n8738 c_3_11_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02170 n8738 c_3_11_cout c_4_10_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02169 vss p_4_10_pi2j n8732 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02168 n8732 c_4_10_a n8731 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02167 n8731 c_3_11_cout n8733 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02166 vss p_4_10_pi2j n8733 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02165 n8733 c_4_10_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02164 vss n8731 c_5_9_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02163 p_4_10_pi2j c_4_10_a c_4_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02162 vss n9124 c_4_9_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02161 n8838 p_4_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02160 vss c_4_9_a n8838 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02159 n9124 c_4_9_cin n8838 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02158 n8837 p_4_9_pi2j n9124 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02157 vss c_4_9_a n8837 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02156 n9119 c_4_9_cin c_4_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02155 c_4_9_s2_s n9119 c_4_9_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02154 c_4_9_a p_4_9_pi2j c_4_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02153 c_4_9_s1_s c_4_9_a p_4_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02152 c_5_7_a c_4_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02151 vss c_4_9_s1_s n9119 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02150 n9131 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02149 vss a_7 n8840 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02148 n8840 p_4_2_d2j n9129 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02147 n9129 p_4_2_d2jbar n8839 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02146 n8839 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02145 vss p_4_9_t_s p_4_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02144 p_4_9_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02143 n9129 n9131 p_4_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02142 p_4_9_t_s n9129 n9131 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02141 n9488 p_4_2_d2j n9487 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02140 n9485 p_4_2_d2jbar n9488 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02139 p_4_8_t_s n9488 n9486 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02138 n9488 n9486 p_4_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02137 p_4_8_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02136 vss p_4_8_t_s p_4_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02135 n9486 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02134 vss a_7 n9485 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02133 n9487 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02132 vss c_4_8_s1_s n9474 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02131 c_5_6_a c_4_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02130 c_4_8_s1_s p_4_8_pi2j c_4_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02129 c_4_8_s2_s n9474 c_3_9_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02128 n9474 c_3_9_cout c_4_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02127 vss p_4_8_pi2j n9477 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02126 n9477 c_4_8_a n9479 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02125 n9479 c_3_9_cout n9478 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02124 vss p_4_8_pi2j n9478 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02123 n9478 c_4_8_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02122 vss n9479 c_5_7_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02121 p_4_8_pi2j c_4_8_a c_4_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02120 vss n9917 c_4_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02119 n9595 p_4_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02118 vss c_4_7_a n9595 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02117 n9917 c_4_7_cin n9595 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02116 n9476 p_4_7_pi2j n9917 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02115 vss c_4_7_a n9476 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_02114 n9912 c_4_7_cin c_4_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02113 c_4_7_s2_s n9912 c_4_7_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02112 c_4_7_a p_4_7_pi2j c_4_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02111 c_4_7_s1_s c_4_7_a p_4_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02110 c_5_5_a c_4_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02109 vss c_4_7_s1_s n9912 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02108 n9923 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02107 vss a_5 n9599 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02106 n9599 p_4_2_d2j n9918 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02105 n9918 p_4_2_d2jbar n9598 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02104 n9598 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02103 vss p_4_7_t_s p_4_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02102 p_4_7_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02101 n9918 n9923 p_4_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02100 p_4_7_t_s n9918 n9923 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02099 n10257 p_4_2_d2j n10048 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02098 n10049 p_4_2_d2jbar n10257 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02097 p_4_6_t_s n10257 n10259 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02096 n10257 n10259 p_4_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02095 p_4_6_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02094 vss p_4_6_t_s p_4_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02093 n10259 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02092 vss a_5 n10049 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02091 n10048 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02090 vss c_4_6_s1_s n10047 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02089 c_5_4_a c_4_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02088 c_4_6_s1_s p_4_6_pi2j c_4_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02087 c_4_6_s2_s n10047 c_3_7_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02086 n10047 c_3_7_cout c_4_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02085 vss p_4_6_pi2j n10253 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02084 n10253 c_4_6_a n10252 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02083 n10252 c_3_7_cout n10248 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02082 vss p_4_6_pi2j n10248 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02081 n10248 c_4_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02080 vss n10252 c_5_5_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02079 p_4_6_pi2j c_4_6_a c_4_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02078 vss n10682 c_4_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02077 n10420 c_4_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02076 vss c_4_5_a n10420 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02075 n10682 c_4_5_cin n10420 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02074 n10251 c_4_5_b n10682 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02073 vss c_4_5_a n10251 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02072 n10425 c_4_5_cin c_4_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02071 c_4_5_s2_s n10425 c_4_5_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02070 c_4_5_a c_4_5_b c_4_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02069 c_4_5_s1_s c_4_5_a c_4_5_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02068 c_5_3_a c_4_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02067 vss c_4_5_s1_s n10425 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02066 n10686 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02065 vss a_3 n10261 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02064 n10261 p_4_2_d2j n10683 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02063 n10683 p_4_2_d2jbar n10260 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02062 n10260 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02061 vss p_4_5_t_s c_4_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02060 c_4_5_b p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02059 n10683 n10686 p_4_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02058 p_4_5_t_s n10683 n10686 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02057 n10864 p_4_2_d2j n10862 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02056 n10863 p_4_2_d2jbar n10864 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02055 p_4_4_t_s n10864 n10861 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02054 n10864 n10861 p_4_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02053 p_4_4_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02052 vss p_4_4_t_s p_4_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_02051 n10861 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02050 vss a_3 n10863 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02049 n10862 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02048 vss c_4_4_s1_s n10860 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02047 c_5_2_a c_4_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02046 c_4_4_s1_s p_4_4_pi2j c_4_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02045 c_4_4_s2_s n10860 c_3_5_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02044 n10860 c_3_5_cout c_4_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02043 vss p_4_4_pi2j n11012 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02042 n11012 c_4_4_a n10855 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02041 n10855 c_3_5_cout n11008 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02040 vss p_4_4_pi2j n11008 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02039 n11008 c_4_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02038 vss n10855 c_5_3_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02037 p_4_4_pi2j c_4_4_a c_4_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02036 vss n11221 c_4_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_02035 n11011 c_4_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02034 vss c_4_3_a n11011 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02033 n11221 c_4_3_cin n11011 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02032 n11010 c_4_3_b n11221 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02031 vss c_4_3_a n11010 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02030 n11223 c_4_3_cin c_4_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02029 c_4_3_s2_s n11223 c_4_3_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02028 c_4_3_a c_4_3_b c_4_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02027 c_4_3_s1_s c_4_3_a c_4_3_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02026 c_5_1_a c_4_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02025 vss c_4_3_s1_s n11223 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02024 n11228 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02023 vss a_1 n11016 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02022 n11016 p_4_2_d2j n11225 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02021 n11225 p_4_2_d2jbar n11015 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02020 n11015 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02019 vss p_4_3_t_s c_4_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02018 c_4_3_b p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02017 n11225 n11228 p_4_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02016 p_4_3_t_s n11225 n11228 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02015 n11653 p_4_2_d2j n11651 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02014 n11652 p_4_2_d2jbar n11653 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_02013 p_4_2_t_s n11653 n11650 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02012 n11653 n11650 p_4_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02011 c_4_2_b p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02010 vss p_4_2_t_s c_4_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_02009 n11650 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02008 vss a_1 n11652 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02007 n11651 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02006 vss c_4_2_s1_s n11646 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_02005 c_4_2_sum c_4_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02004 c_4_2_s1_s c_4_2_b c_4_2_a vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02003 c_4_2_s2_s n11646 c_3_3_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02002 n11646 c_3_3_cout c_4_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_02001 vss c_4_2_b n11641 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_02000 n11641 c_4_2_a n11643 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01999 n11643 c_3_3_cout n11642 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01998 vss c_4_2_b n11642 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01997 n11642 c_4_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01996 vss n11643 c_5_1_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01995 c_4_2_b c_4_2_a c_4_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01994 vss n12025 c_4_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01993 n11755 p_4_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01992 vss c_4_1_a n11755 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01991 n12025 c_4_1_cin n11755 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01990 n11754 p_4_1_pi2j n12025 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01989 vss c_4_1_a n11754 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01988 n12024 c_4_1_cin c_4_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01987 c_4_1_s2_s n12024 c_4_1_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01986 c_4_1_a p_4_1_pi2j c_4_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01985 c_4_1_s1_s c_4_1_a p_4_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01984 c_4_1_sum c_4_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01983 vss c_4_1_s1_s n12024 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01982 n12034 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01981 n12035 p_4_2_d2jbar n11758 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01980 n11758 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01979 vss p_4_1_t_s p_4_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01978 p_4_1_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01977 n12035 n12034 p_4_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01976 p_4_1_t_s n12035 n12034 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01975 cl4_4_s1_s n12392 c_3_1_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01974 n12392 c_3_1_sum cl4_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01973 vss cl4_4_s1_s p_4 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01972 vss c_3_1_sum n12382 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01971 n12382 n12392 n12381 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01970 n12380 n12381 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01969 n12378 c_3_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01968 vss c_3_2_sum n12378 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01967 n12379 c_3_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01966 n12377 c_3_1_cout n12379 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01965 n12374 c_3_1_sum n12377 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01964 n12378 n12392 n12374 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01963 n12375 n12377 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01962 cl4_4_s2_s c_3_1_cout c_3_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01961 c_3_1_cout c_3_2_sum cl4_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01960 vss cl4_4_s2_s n12372 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01959 cl4_4_s3_s n12372 n12380 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01958 n12372 n12380 cl4_4_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01957 vss cl4_4_s3_s p_5 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01956 vss c_3_33_s1_s n238 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01955 c_4_31_a c_3_33_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01954 c_3_33_s1_s c_3_31_a p_3_33_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01953 c_3_31_a p_3_33_pi2j c_3_33_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01952 c_3_33_s2_s n238 c_3_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01951 n238 c_3_32_cin c_3_33_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01950 vss c_3_31_a n31 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01949 n31 p_3_33_pi2j n230 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01948 n230 c_3_32_cin n32 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01947 vss c_3_31_a n32 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01946 n32 p_3_33_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01945 vss n230 c_4_32_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01944 n240 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01943 n243 a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01942 vss p_3_33_t_s p_3_33_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01941 p_3_33_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01940 n243 n240 p_3_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01939 p_3_33_t_s n243 n240 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01938 n580 p_3_2_d2j n581 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01937 n579 p_3_2_d2jbar n580 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01936 p_3_32_t_s n580 n578 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01935 n580 n578 p_3_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01934 p_3_32_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01933 vss p_3_32_t_s p_3_32_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01932 n578 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01931 vss a_31 n579 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01930 n581 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01929 vss c_3_32_s1_s n574 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01928 c_4_30_a c_3_32_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01927 c_3_32_s1_s p_3_32_pi2j c_3_31_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01926 c_3_32_s2_s n574 c_3_32_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01925 n574 c_3_32_cin c_3_32_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01924 vss p_3_32_pi2j n570 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01923 n570 c_3_31_a n569 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01922 n569 c_3_32_cin n571 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01921 vss p_3_32_pi2j n571 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01920 n571 c_3_31_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01919 vss n569 c_4_31_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01918 p_3_32_pi2j c_3_31_a c_3_32_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01917 vss n936 c_3_31_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01916 n658 p_3_31_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01915 vss c_3_31_a n658 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01914 n936 c_3_31_cin n658 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01913 n657 p_3_31_pi2j n936 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01912 vss c_3_31_a n657 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01911 n944 c_3_31_cin c_3_31_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01910 c_3_31_s2_s n944 c_3_31_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01909 c_3_31_a p_3_31_pi2j c_3_31_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01908 c_3_31_s1_s c_3_31_a p_3_31_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01907 c_4_29_a c_3_31_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01906 vss c_3_31_s1_s n944 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01905 n945 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01904 vss a_29 n659 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01903 n659 p_3_2_d2j n948 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01902 n948 p_3_2_d2jbar n660 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01901 n660 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01900 vss p_3_31_t_s p_3_31_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01899 p_3_31_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01898 n948 n945 p_3_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01897 p_3_31_t_s n948 n945 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01896 n1346 p_3_2_d2j n1344 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01895 n1345 p_3_2_d2jbar n1346 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01894 p_3_30_t_s n1346 n1343 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01893 n1346 n1343 p_3_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01892 p_3_30_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01891 vss p_3_30_t_s p_3_30_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01890 n1343 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01889 vss a_29 n1345 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01888 n1344 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01887 vss c_3_30_s1_s n1338 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01886 c_4_28_a c_3_30_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01885 c_3_30_s1_s p_3_30_pi2j c_3_30_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01884 c_3_30_s2_s n1338 c_2_31_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01883 n1338 c_2_31_cout c_3_30_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01882 vss p_3_30_pi2j n1335 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01881 n1335 c_3_30_a n1333 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01880 n1333 c_2_31_cout n1334 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01879 vss p_3_30_pi2j n1334 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01878 n1334 c_3_30_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01877 vss n1333 c_4_29_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01876 p_3_30_pi2j c_3_30_a c_3_30_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01875 vss n1721 c_3_29_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01874 n1418 p_3_29_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01873 vss c_3_29_a n1418 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01872 n1721 c_3_29_cin n1418 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01871 n1332 p_3_29_pi2j n1721 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01870 vss c_3_29_a n1332 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01869 n1728 c_3_29_cin c_3_29_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01868 c_3_29_s2_s n1728 c_3_29_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01867 c_3_29_a p_3_29_pi2j c_3_29_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01866 c_3_29_s1_s c_3_29_a p_3_29_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01865 c_4_27_a c_3_29_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01864 vss c_3_29_s1_s n1728 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01863 n1731 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01862 vss a_27 n1419 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01861 n1419 p_3_2_d2j n1734 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01860 n1734 p_3_2_d2jbar n1420 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01859 n1420 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01858 vss p_3_29_t_s p_3_29_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01857 p_3_29_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01856 n1734 n1731 p_3_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01855 p_3_29_t_s n1734 n1731 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01854 n2095 p_3_2_d2j n2096 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01853 n2094 p_3_2_d2jbar n2095 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01852 p_3_28_t_s n2095 n2093 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01851 n2095 n2093 p_3_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01850 p_3_28_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01849 vss p_3_28_t_s p_3_28_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01848 n2093 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01847 vss a_27 n2094 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01846 n2096 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01845 vss c_3_28_s1_s n1866 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01844 c_4_26_a c_3_28_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01843 c_3_28_s1_s p_3_28_pi2j c_3_28_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01842 c_3_28_s2_s n1866 c_2_29_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01841 n1866 c_2_29_cout c_3_28_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01840 vss p_3_28_pi2j n2086 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01839 n2086 c_3_28_a n2085 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01838 n2085 c_2_29_cout n2084 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01837 vss p_3_28_pi2j n2084 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01836 n2084 c_3_28_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01835 vss n2085 c_4_27_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01834 p_3_28_pi2j c_3_28_a c_3_28_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01833 vss n2534 c_3_27_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01832 n2225 c_3_27_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01831 vss c_3_27_a n2225 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01830 n2534 c_3_27_cin n2225 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01829 n2083 c_3_27_b n2534 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01828 vss c_3_27_a n2083 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01827 n2531 c_3_27_cin c_3_27_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01826 c_3_27_s2_s n2531 c_3_27_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01825 c_3_27_a c_3_27_b c_3_27_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01824 c_3_27_s1_s c_3_27_a c_3_27_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01823 c_4_25_a c_3_27_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01822 vss c_3_27_s1_s n2531 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01821 n2543 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01820 vss a_25 n2231 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01819 n2231 p_3_2_d2j n2542 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01818 n2542 p_3_2_d2jbar n2230 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01817 n2230 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01816 vss p_3_27_t_s c_3_27_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01815 c_3_27_b p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01814 n2542 n2543 p_3_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01813 p_3_27_t_s n2542 n2543 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01812 n2698 p_3_2_d2j n2699 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01811 n2697 p_3_2_d2jbar n2698 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01810 p_3_26_t_s n2698 n2696 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01809 n2698 n2696 p_3_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01808 p_3_26_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01807 vss p_3_26_t_s p_3_26_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01806 n2696 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01805 vss a_25 n2697 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01804 n2699 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01803 vss c_3_26_s1_s n2695 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01802 c_4_24_a c_3_26_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01801 c_3_26_s1_s p_3_26_pi2j c_3_26_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01800 c_3_26_s2_s n2695 c_2_27_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01799 n2695 c_2_27_cout c_3_26_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01798 vss p_3_26_pi2j n2893 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01797 n2893 c_3_26_a n2892 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01796 n2892 c_2_27_cout n2894 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01795 vss p_3_26_pi2j n2894 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01794 n2894 c_3_26_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01793 vss n2892 c_4_25_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01792 p_3_26_pi2j c_3_26_a c_3_26_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01791 vss n3310 c_3_25_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01790 n2891 c_3_25_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01789 vss c_3_25_a n2891 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01788 n3310 c_3_25_cin n2891 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01787 n2890 c_3_25_b n3310 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01786 vss c_3_25_a n2890 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01785 n3058 c_3_25_cin c_3_25_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01784 c_3_25_s2_s n3058 c_3_25_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01783 c_3_25_a c_3_25_b c_3_25_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01782 c_3_25_s1_s c_3_25_a c_3_25_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01781 c_4_23_a c_3_25_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01780 vss c_3_25_s1_s n3058 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01779 n3320 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01778 vss a_23 n2900 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01777 n2900 p_3_2_d2j n3060 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01776 n3060 p_3_2_d2jbar n2901 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01775 n2901 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01774 vss p_3_25_t_s c_3_25_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01773 c_3_25_b p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01772 n3060 n3320 p_3_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01771 p_3_25_t_s n3060 n3320 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01770 n3505 p_3_2_d2j n3506 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01769 n3504 p_3_2_d2jbar n3505 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01768 p_3_24_t_s n3505 n3503 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01767 n3505 n3503 p_3_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01766 c_3_24_b p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01765 vss p_3_24_t_s c_3_24_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01764 n3503 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01763 vss a_23 n3504 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01762 n3506 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01761 vss c_3_24_s1_s n3500 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01760 c_4_22_a c_3_24_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01759 c_3_24_s1_s c_3_24_b c_3_24_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01758 c_3_24_s2_s n3500 c_2_25_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01757 n3500 c_2_25_cout c_3_24_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01756 vss c_3_24_b n3643 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01755 n3643 c_3_24_a n3496 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01754 n3496 c_2_25_cout n3642 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01753 vss c_3_24_b n3642 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01752 n3642 c_3_24_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01751 vss n3496 c_4_23_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01750 c_3_24_b c_3_24_a c_3_24_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01749 vss n3901 c_3_23_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01748 n3641 c_3_23_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01747 vss c_3_23_a n3641 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01746 n3901 c_3_23_cin n3641 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01745 n3640 c_3_23_b n3901 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01744 vss c_3_23_a n3640 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01743 n3908 c_3_23_cin c_3_23_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01742 c_3_23_s2_s n3908 c_3_23_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01741 c_3_23_a c_3_23_b c_3_23_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01740 c_3_23_s1_s c_3_23_a c_3_23_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01739 c_4_21_a c_3_23_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01738 vss c_3_23_s1_s n3908 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01737 n3909 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01736 vss a_21 n3646 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01735 n3646 p_3_2_d2j n3912 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01734 n3912 p_3_2_d2jbar n3647 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01733 n3647 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01732 vss p_3_23_t_s c_3_23_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01731 c_3_23_b p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01730 n3912 n3909 p_3_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01729 p_3_23_t_s n3912 n3909 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01728 n4322 p_3_2_d2j n4323 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01727 n4321 p_3_2_d2jbar n4322 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01726 p_3_22_t_s n4322 n4320 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01725 n4322 n4320 p_3_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01724 p_3_22_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01723 vss p_3_22_t_s p_3_22_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01722 n4320 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01721 vss a_21 n4321 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01720 n4323 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01719 vss c_3_22_s1_s n4315 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01718 c_4_20_a c_3_22_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01717 c_3_22_s1_s p_3_22_pi2j c_3_22_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01716 c_3_22_s2_s n4315 c_2_23_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01715 n4315 c_2_23_cout c_3_22_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01714 vss p_3_22_pi2j n4311 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01713 n4311 c_3_22_a n4310 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01712 n4310 c_2_23_cout n4312 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01711 vss p_3_22_pi2j n4312 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01710 n4312 c_3_22_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01709 vss n4310 c_4_21_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01708 p_3_22_pi2j c_3_22_a c_3_22_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01707 vss n4683 c_3_21_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01706 n4409 p_3_21_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01705 vss c_3_21_a n4409 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01704 n4683 c_3_21_cin n4409 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01703 n4408 p_3_21_pi2j n4683 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01702 vss c_3_21_a n4408 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01701 n4688 c_3_21_cin c_3_21_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01700 c_3_21_s2_s n4688 c_3_21_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01699 c_3_21_a p_3_21_pi2j c_3_21_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01698 c_3_21_s1_s c_3_21_a p_3_21_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01697 c_4_19_a c_3_21_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01696 vss c_3_21_s1_s n4688 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01695 n4692 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01694 vss a_19 n4410 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01693 n4410 p_3_2_d2j n4695 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01692 n4695 p_3_2_d2jbar n4411 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01691 n4411 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01690 vss p_3_21_t_s p_3_21_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01689 p_3_21_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01688 n4695 n4692 p_3_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01687 p_3_21_t_s n4695 n4692 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01686 n5068 p_3_2_d2j n5069 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01685 n5067 p_3_2_d2jbar n5068 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01684 p_3_20_t_s n5068 n5066 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01683 n5068 n5066 p_3_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01682 p_3_20_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01681 vss p_3_20_t_s p_3_20_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01680 n5066 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01679 vss a_19 n5067 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01678 n5069 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01677 vss c_3_20_s1_s n5061 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01676 c_4_18_a c_3_20_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01675 c_3_20_s1_s p_3_20_pi2j c_3_20_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01674 c_3_20_s2_s n5061 c_2_21_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01673 n5061 c_2_21_cout c_3_20_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01672 vss p_3_20_pi2j n5057 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01671 n5057 c_3_20_a n5058 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01670 n5058 c_2_21_cout n5056 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01669 vss p_3_20_pi2j n5056 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01668 n5056 c_3_20_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01667 vss n5058 c_4_19_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01666 p_3_20_pi2j c_3_20_a c_3_20_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01665 vss n5448 c_3_19_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01664 n5150 p_3_19_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01663 vss c_3_19_a n5150 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01662 n5448 c_3_19_cin n5150 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01661 n5149 p_3_19_pi2j n5448 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01660 vss c_3_19_a n5149 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01659 n5455 c_3_19_cin c_3_19_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01658 c_3_19_s2_s n5455 c_3_19_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01657 c_3_19_a p_3_19_pi2j c_3_19_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01656 c_3_19_s1_s c_3_19_a p_3_19_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01655 c_4_17_a c_3_19_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01654 vss c_3_19_s1_s n5455 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01653 n5458 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01652 vss a_17 n5151 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01651 n5151 p_3_2_d2j n5461 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01650 n5461 p_3_2_d2jbar n5152 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01649 n5152 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01648 vss p_3_19_t_s p_3_19_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01647 p_3_19_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01646 n5461 n5458 p_3_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01645 p_3_19_t_s n5461 n5458 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01644 n5822 p_3_2_d2j n5821 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01643 n5819 p_3_2_d2jbar n5822 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01642 p_3_18_t_s n5822 n5820 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01641 n5822 n5820 p_3_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01640 p_3_18_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01639 vss p_3_18_t_s p_3_18_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01638 n5820 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01637 vss a_17 n5819 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01636 n5821 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01635 vss c_3_18_s1_s n5592 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01634 c_4_16_a c_3_18_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01633 c_3_18_s1_s p_3_18_pi2j c_3_18_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01632 c_3_18_s2_s n5592 c_2_19_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01631 n5592 c_2_19_cout c_3_18_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01630 vss p_3_18_pi2j n5810 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01629 n5810 c_3_18_a n5812 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01628 n5812 c_2_19_cout n5811 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01627 vss p_3_18_pi2j n5811 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01626 n5811 c_3_18_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01625 vss n5812 c_4_17_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01624 p_3_18_pi2j c_3_18_a c_3_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01623 vss n6247 c_3_17_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01622 n5922 p_3_17_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01621 vss c_3_17_a n5922 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01620 n6247 c_3_17_cin n5922 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01619 n5809 p_3_17_pi2j n6247 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01618 vss c_3_17_a n5809 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01617 n6243 c_3_17_cin c_3_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01616 c_3_17_s2_s n6243 c_3_17_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01615 c_3_17_a p_3_17_pi2j c_3_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01614 c_3_17_s1_s c_3_17_a p_3_17_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01613 c_4_15_a c_3_17_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01612 vss c_3_17_s1_s n6243 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01611 n6258 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01610 vss a_15 n5925 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01609 n5925 p_3_2_d2j n6257 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01608 n6257 p_3_2_d2jbar n5926 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01607 n5926 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01606 vss p_3_17_t_s p_3_17_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01605 p_3_17_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01604 n6257 n6258 p_3_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01603 p_3_17_t_s n6257 n6258 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01602 n6395 p_3_2_d2j n6396 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01601 n6394 p_3_2_d2jbar n6395 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01600 p_3_16_t_s n6395 n6597 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01599 n6395 n6597 p_3_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01598 p_3_16_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01597 vss p_3_16_t_s p_3_16_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01596 n6597 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01595 vss a_15 n6394 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01594 n6396 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01593 vss c_3_16_s1_s n6393 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01592 c_4_14_a c_3_16_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01591 c_3_16_s1_s p_3_16_pi2j c_3_16_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01590 c_3_16_s2_s n6393 c_2_17_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01589 n6393 c_2_17_cout c_3_16_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01588 vss p_3_16_pi2j n6591 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01587 n6591 c_3_16_a n6592 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01586 n6592 c_2_17_cout n6590 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01585 vss p_3_16_pi2j n6590 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01584 n6590 c_3_16_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01583 vss n6592 c_4_15_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01582 p_3_16_pi2j c_3_16_a c_3_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01581 vss n7012 c_3_15_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01580 n6589 c_3_15_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01579 vss c_3_15_a n6589 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01578 n7012 c_3_15_cin n6589 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01577 n6588 c_3_15_b n7012 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01576 vss c_3_15_a n6588 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01575 n6759 c_3_15_cin c_3_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01574 c_3_15_s2_s n6759 c_3_15_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01573 c_3_15_a c_3_15_b c_3_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01572 c_3_15_s1_s c_3_15_a c_3_15_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01571 c_4_13_a c_3_15_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01570 vss c_3_15_s1_s n6759 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01569 n7021 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01568 vss a_13 n6599 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01567 n6599 p_3_2_d2j n6761 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01566 n6761 p_3_2_d2jbar n6600 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01565 n6600 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01564 vss p_3_15_t_s c_3_15_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01563 c_3_15_b p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01562 n6761 n7021 p_3_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01561 p_3_15_t_s n6761 n7021 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01560 n7199 p_3_2_d2j n7200 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01559 n7198 p_3_2_d2jbar n7199 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01558 p_3_14_t_s n7199 n7197 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01557 n7199 n7197 p_3_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01556 p_3_14_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01555 vss p_3_14_t_s p_3_14_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01554 n7197 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01553 vss a_13 n7198 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01552 n7200 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01551 vss c_3_14_s1_s n7194 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01550 c_4_12_a c_3_14_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01549 c_3_14_s1_s p_3_14_pi2j c_3_14_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01548 c_3_14_s2_s n7194 c_2_15_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01547 n7194 c_2_15_cout c_3_14_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01546 vss p_3_14_pi2j n7351 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01545 n7351 c_3_14_a n7191 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01544 n7191 c_2_15_cout n7352 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01543 vss p_3_14_pi2j n7352 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01542 n7352 c_3_14_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01541 vss n7191 c_4_13_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01540 p_3_14_pi2j c_3_14_a c_3_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01539 vss n7565 c_3_13_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01538 n7350 c_3_13_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01537 vss c_3_13_a n7350 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01536 n7565 c_3_13_cin n7350 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01535 n7349 c_3_13_b n7565 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01534 vss c_3_13_a n7349 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01533 n7571 c_3_13_cin c_3_13_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01532 c_3_13_s2_s n7571 c_3_13_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01531 c_3_13_a c_3_13_b c_3_13_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01530 c_3_13_s1_s c_3_13_a c_3_13_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01529 c_4_11_a c_3_13_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01528 vss c_3_13_s1_s n7571 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01527 n7572 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01526 vss a_11 n7356 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01525 n7356 p_3_2_d2j n7574 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01524 n7574 p_3_2_d2jbar n7357 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01523 n7357 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01522 vss p_3_13_t_s c_3_13_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01521 c_3_13_b p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01520 n7574 n7572 p_3_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01519 p_3_13_t_s n7574 n7572 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01518 n8002 p_3_2_d2j n8003 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01517 n8001 p_3_2_d2jbar n8002 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01516 p_3_12_t_s n8002 n8000 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01515 n8002 n8000 p_3_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01514 c_3_12_b p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01513 vss p_3_12_t_s c_3_12_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01512 n8000 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01511 vss a_11 n8001 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01510 n8003 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01509 vss c_3_12_s1_s n7996 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01508 c_4_10_a c_3_12_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01507 c_3_12_s1_s c_3_12_b c_3_12_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01506 c_3_12_s2_s n7996 c_2_13_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01505 n7996 c_2_13_cout c_3_12_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01504 vss c_3_12_b n7992 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01503 n7992 c_3_12_a n7993 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01502 n7993 c_2_13_cout n7991 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01501 vss c_3_12_b n7991 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01500 n7991 c_3_12_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01499 vss n7993 c_4_11_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01498 c_3_12_b c_3_12_a c_3_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01497 vss n8372 c_3_11_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01496 n8098 p_3_11_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01495 vss c_3_11_a n8098 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01494 n8372 c_3_11_cin n8098 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01493 n8097 p_3_11_pi2j n8372 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01492 vss c_3_11_a n8097 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01491 n8377 c_3_11_cin c_3_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01490 c_3_11_s2_s n8377 c_3_11_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01489 c_3_11_a p_3_11_pi2j c_3_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01488 c_3_11_s1_s c_3_11_a p_3_11_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01487 c_4_9_a c_3_11_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01486 vss c_3_11_s1_s n8377 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01485 n8380 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01484 vss a_9 n8100 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01483 n8100 p_3_2_d2j n8383 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01482 n8383 p_3_2_d2jbar n8101 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01481 n8101 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01480 vss p_3_11_t_s p_3_11_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01479 p_3_11_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01478 n8383 n8380 p_3_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01477 p_3_11_t_s n8383 n8380 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01476 n8757 p_3_2_d2j n8758 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01475 n8756 p_3_2_d2jbar n8757 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01474 p_3_10_t_s n8757 n8755 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01473 n8757 n8755 p_3_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01472 p_3_10_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01471 vss p_3_10_t_s p_3_10_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01470 n8755 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01469 vss a_9 n8756 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01468 n8758 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01467 vss c_3_10_s1_s n8750 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01466 c_4_8_a c_3_10_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01465 c_3_10_s1_s p_3_10_pi2j c_3_10_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01464 c_3_10_s2_s n8750 c_2_11_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01463 n8750 c_2_11_cout c_3_10_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01462 vss p_3_10_pi2j n8747 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01461 n8747 c_3_10_a n8745 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01460 n8745 c_2_11_cout n8746 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01459 vss p_3_10_pi2j n8746 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01458 n8746 c_3_10_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01457 vss n8745 c_4_9_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01456 p_3_10_pi2j c_3_10_a c_3_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01455 vss n9136 c_3_9_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01454 n8842 p_3_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01453 vss c_3_9_a n8842 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01452 n9136 c_3_9_cin n8842 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01451 n8841 p_3_9_pi2j n9136 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01450 vss c_3_9_a n8841 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01449 n9143 c_3_9_cin c_3_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01448 c_3_9_s2_s n9143 c_3_9_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01447 c_3_9_a p_3_9_pi2j c_3_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01446 c_3_9_s1_s c_3_9_a p_3_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01445 c_4_7_a c_3_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01444 vss c_3_9_s1_s n9143 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01443 n9146 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01442 vss a_7 n8843 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01441 n8843 p_3_2_d2j n9149 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01440 n9149 p_3_2_d2jbar n8844 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01439 n8844 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01438 vss p_3_9_t_s p_3_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01437 p_3_9_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01436 n9149 n9146 p_3_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01435 p_3_9_t_s n9149 n9146 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01434 n9503 p_3_2_d2j n9502 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01433 n9500 p_3_2_d2jbar n9503 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01432 p_3_8_t_s n9503 n9501 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01431 n9503 n9501 p_3_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01430 p_3_8_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01429 vss p_3_8_t_s p_3_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01428 n9501 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01427 vss a_7 n9500 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01426 n9502 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01425 vss c_3_8_s1_s n9493 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01424 c_4_6_a c_3_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01423 c_3_8_s1_s p_3_8_pi2j c_3_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01422 c_3_8_s2_s n9493 c_2_9_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01421 n9493 c_2_9_cout c_3_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01420 vss p_3_8_pi2j n9490 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01419 n9490 c_3_8_a n9491 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01418 n9491 c_2_9_cout n9492 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01417 vss p_3_8_pi2j n9492 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01416 n9492 c_3_8_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01415 vss n9491 c_4_7_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01414 p_3_8_pi2j c_3_8_a c_3_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01413 vss n9930 c_3_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01412 n9600 p_3_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01411 vss c_3_7_a n9600 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01410 n9930 c_3_7_cin n9600 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01409 n9489 p_3_7_pi2j n9930 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01408 vss c_3_7_a n9489 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01407 n9939 c_3_7_cin c_3_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01406 c_3_7_s2_s n9939 c_3_7_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01405 c_3_7_a p_3_7_pi2j c_3_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01404 c_3_7_s1_s c_3_7_a p_3_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01403 c_4_5_a c_3_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01402 vss c_3_7_s1_s n9939 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01401 n9942 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01400 vss a_5 n9603 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01399 n9603 p_3_2_d2j n9941 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01398 n9941 p_3_2_d2jbar n9604 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01397 n9604 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01396 vss p_3_7_t_s p_3_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01395 p_3_7_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01394 n9941 n9942 p_3_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01393 p_3_7_t_s n9941 n9942 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01392 n10271 p_3_2_d2j n10054 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01391 n10053 p_3_2_d2jbar n10271 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01390 p_3_6_t_s n10271 n10272 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01389 n10271 n10272 p_3_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01388 p_3_6_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01387 vss p_3_6_t_s p_3_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01386 n10272 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01385 vss a_5 n10053 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01384 n10054 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01383 vss c_3_6_s1_s n10052 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01382 c_4_4_a c_3_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01381 c_3_6_s1_s p_3_6_pi2j c_3_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01380 c_3_6_s2_s n10052 c_2_7_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01379 n10052 c_2_7_cout c_3_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01378 vss p_3_6_pi2j n10264 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01377 n10264 c_3_6_a n10265 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01376 n10265 c_2_7_cout n10263 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01375 vss p_3_6_pi2j n10263 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01374 n10263 c_3_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01373 vss n10265 c_4_5_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01372 p_3_6_pi2j c_3_6_a c_3_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01371 vss n10692 c_3_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01370 n10429 c_3_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01369 vss c_3_5_a n10429 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01368 n10692 c_3_5_cin n10429 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01367 n10262 c_3_5_b n10692 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01366 vss c_3_5_a n10262 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01365 n10434 c_3_5_cin c_3_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01364 c_3_5_s2_s n10434 c_3_5_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01363 c_3_5_a c_3_5_b c_3_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01362 c_3_5_s1_s c_3_5_a c_3_5_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01361 c_4_3_a c_3_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01360 vss c_3_5_s1_s n10434 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01359 n10701 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01358 vss a_3 n10274 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01357 n10274 p_3_2_d2j n10702 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01356 n10702 p_3_2_d2jbar n10275 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01355 n10275 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01354 vss p_3_5_t_s c_3_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01353 c_3_5_b p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01352 n10702 n10701 p_3_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01351 p_3_5_t_s n10702 n10701 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01350 n10873 p_3_2_d2j n10874 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01349 n10872 p_3_2_d2jbar n10873 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01348 p_3_4_t_s n10873 n10871 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01347 n10873 n10871 p_3_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01346 p_3_4_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01345 vss p_3_4_t_s p_3_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01344 n10871 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01343 vss a_3 n10872 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01342 n10874 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01341 vss c_3_4_s1_s n10870 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01340 c_4_2_a c_3_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01339 c_3_4_s1_s p_3_4_pi2j c_3_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01338 c_3_4_s2_s n10870 c_2_5_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01337 n10870 c_2_5_cout c_3_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01336 vss p_3_4_pi2j n11019 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01335 n11019 c_3_4_a n10865 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01334 n10865 c_2_5_cout n11020 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01333 vss p_3_4_pi2j n11020 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01332 n11020 c_3_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01331 vss n10865 c_4_3_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01330 p_3_4_pi2j c_3_4_a c_3_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01329 vss n11230 c_3_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01328 n11018 c_3_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01327 vss c_3_3_a n11018 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01326 n11230 c_3_3_cin n11018 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01325 n11017 c_3_3_b n11230 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01324 vss c_3_3_a n11017 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01323 n11236 c_3_3_cin c_3_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01322 c_3_3_s2_s n11236 c_3_3_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01321 c_3_3_a c_3_3_b c_3_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01320 c_3_3_s1_s c_3_3_a c_3_3_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01319 c_4_1_a c_3_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01318 vss c_3_3_s1_s n11236 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01317 n11237 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01316 vss a_1 n11024 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01315 n11024 p_3_2_d2j n11239 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01314 n11239 p_3_2_d2jbar n11025 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01313 n11025 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01312 vss p_3_3_t_s c_3_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01311 c_3_3_b p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01310 n11239 n11237 p_3_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01309 p_3_3_t_s n11239 n11237 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01308 n11665 p_3_2_d2j n11666 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01307 n11664 p_3_2_d2jbar n11665 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01306 p_3_2_t_s n11665 n11663 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01305 n11665 n11663 p_3_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01304 c_3_2_b p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01303 vss p_3_2_t_s c_3_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01302 n11663 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01301 vss a_1 n11664 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01300 n11666 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01299 vss c_3_2_s1_s n11659 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01298 c_3_2_sum c_3_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01297 c_3_2_s1_s c_3_2_b c_3_2_a vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01296 c_3_2_s2_s n11659 c_2_3_cout vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01295 n11659 c_2_3_cout c_3_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01294 vss c_3_2_b n11655 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01293 n11655 c_3_2_a n11656 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01292 n11656 c_2_3_cout n11654 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01291 vss c_3_2_b n11654 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01290 n11654 c_3_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01289 vss n11656 c_4_1_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01288 c_3_2_b c_3_2_a c_3_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01287 vss n12039 c_3_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01286 n11760 p_3_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01285 vss c_3_1_a n11760 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01284 n12039 c_3_1_cin n11760 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01283 n11759 p_3_1_pi2j n12039 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01282 vss c_3_1_a n11759 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01281 n12046 c_3_1_cin c_3_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01280 c_3_1_s2_s n12046 c_3_1_cin vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01279 c_3_1_a p_3_1_pi2j c_3_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01278 c_3_1_s1_s c_3_1_a p_3_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01277 c_3_1_sum c_3_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01276 vss c_3_1_s1_s n12046 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01275 n12050 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01274 n12054 p_3_2_d2jbar n11763 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01273 n11763 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01272 vss p_3_1_t_s p_3_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01271 p_3_1_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01270 n12054 n12050 p_3_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01269 p_3_1_t_s n12054 n12050 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01268 cl4_3_s1_s n12406 c_2_1_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01267 n12406 c_2_1_sum cl4_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01266 vss cl4_3_s1_s p_2 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01265 vss c_2_1_sum n12399 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01264 n12399 n12406 n12397 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01263 n12398 n12397 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01262 n12396 c_2_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01261 vss c_2_2_sum n12396 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01260 n12393 c_2_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01259 n12394 c_2_1_cout n12393 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01258 n12391 c_2_1_sum n12394 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01257 n12396 n12406 n12391 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01256 n12392 n12394 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01255 cl4_3_s2_s c_2_1_cout c_2_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01254 c_2_1_cout c_2_2_sum cl4_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01253 vss cl4_3_s2_s n12390 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01252 cl4_3_s3_s n12390 n12398 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01251 n12390 n12398 cl4_3_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01250 vss cl4_3_s3_s p_3 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01249 vss n248 c_3_32_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01248 n34 p_2_33_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01247 vss c_2_31_a n34 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01246 n248 vss n34 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01245 n33 p_2_33_pi2j n248 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01244 vss c_2_31_a n33 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01243 n251 vss c_2_33_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01242 c_2_33_s2_s n251 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01241 c_2_31_a p_2_33_pi2j c_2_33_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01240 c_2_33_s1_s c_2_31_a p_2_33_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01239 c_3_31_a c_2_33_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01238 vss c_2_33_s1_s n251 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01237 n255 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01236 n258 a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01235 vss p_2_33_t_s p_2_33_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01234 p_2_33_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01233 n258 n255 p_2_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01232 p_2_33_t_s n258 n255 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01231 n590 p_2_2_d2j n589 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01230 n588 p_2_2_d2jbar n590 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01229 p_2_32_t_s n590 n586 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01228 n590 n586 p_2_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01227 c_2_32_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01226 vss p_2_32_t_s c_2_32_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01225 n586 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01224 vss a_31 n588 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01223 n589 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01222 c_3_31_cin n583 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01221 vss c_2_31_a n582 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01220 n582 c_2_32_b n583 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01219 c_2_32_b c_2_31_a c_2_32_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01218 c_2_32_s1_s c_2_32_b c_2_31_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01217 c_3_30_a c_2_32_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_01216 vss n955 c_2_31_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01215 n662 p_2_31_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01214 vss c_2_31_a n662 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01213 n955 vss n662 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01212 n661 p_2_31_pi2j n955 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01211 vss c_2_31_a n661 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01210 n958 vss c_2_31_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01209 c_2_31_s2_s n958 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01208 c_2_31_a p_2_31_pi2j c_2_31_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01207 c_2_31_s1_s c_2_31_a p_2_31_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01206 c_3_29_a c_2_31_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01205 vss c_2_31_s1_s n958 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01204 n963 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01203 vss a_29 n663 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01202 n663 p_2_2_d2j n968 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01201 n968 p_2_2_d2jbar n664 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01200 n664 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01199 vss p_2_31_t_s p_2_31_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01198 p_2_31_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01197 n968 n963 p_2_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01196 p_2_31_t_s n968 n963 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01195 n1355 p_2_2_d2j n1357 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01194 n1356 p_2_2_d2jbar n1355 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01193 p_2_30_t_s n1355 n1354 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01192 n1355 n1354 p_2_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01191 p_2_30_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01190 vss p_2_30_t_s p_2_30_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01189 n1354 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01188 vss a_29 n1356 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01187 n1357 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01186 c_3_29_cin n1349 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01185 vss c_2_30_a n1348 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01184 n1348 p_2_30_pi2j n1349 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01183 p_2_30_pi2j c_2_30_a c_2_30_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01182 c_2_30_s1_s p_2_30_pi2j c_2_30_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01181 c_3_28_a c_2_30_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_01180 vss n1739 c_2_29_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01179 n1421 p_2_29_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01178 vss c_2_29_a n1421 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01177 n1739 p_18_1_c2j n1421 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01176 n1347 p_2_29_pi2j n1739 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01175 vss c_2_29_a n1347 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01174 n1745 p_18_1_c2j c_2_29_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01173 c_2_29_s2_s n1745 p_18_1_c2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01172 c_2_29_a p_2_29_pi2j c_2_29_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01171 c_2_29_s1_s c_2_29_a p_2_29_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01170 c_3_27_a c_2_29_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01169 vss c_2_29_s1_s n1745 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01168 n1751 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01167 vss a_27 n1422 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01166 n1422 p_2_2_d2j n1754 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01165 n1754 p_2_2_d2jbar n1423 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01164 n1423 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01163 vss p_2_29_t_s p_2_29_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01162 p_2_29_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01161 n1754 n1751 p_2_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01160 p_2_29_t_s n1754 n1751 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01159 n2106 p_2_2_d2j n2105 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01158 n2107 p_2_2_d2jbar n2106 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01157 p_2_28_t_s n2106 n2104 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01156 n2106 n2104 p_2_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01155 p_2_28_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01154 vss p_2_28_t_s p_2_28_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01153 n2104 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01152 vss a_27 n2107 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01151 n2105 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01150 c_3_27_cin n2099 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01149 vss c_2_28_a n2098 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01148 n2098 p_2_28_pi2j n2099 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01147 p_2_28_pi2j c_2_28_a c_2_28_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01146 c_2_28_s1_s p_2_28_pi2j c_2_28_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01145 c_3_26_a c_2_28_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_01144 vss n2552 c_2_27_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01143 n2232 c_2_27_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01142 vss n2555 n2232 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01141 n2552 p_17_1_c2j n2232 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01140 n2097 c_2_27_b n2552 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01139 vss n2555 n2097 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_01138 n2551 p_17_1_c2j c_2_27_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01137 c_2_27_s2_s n2551 p_17_1_c2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01136 n2555 c_2_27_b c_2_27_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01135 c_2_27_s1_s n2555 c_2_27_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01134 c_3_25_a c_2_27_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01133 vss c_2_27_s1_s n2551 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01132 n2560 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01131 vss a_25 n2238 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01130 n2238 p_2_2_d2j n2561 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01129 n2561 p_2_2_d2jbar n2239 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01128 n2239 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01127 vss p_2_27_t_s c_2_27_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01126 c_2_27_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01125 n2561 n2560 p_2_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01124 p_2_27_t_s n2561 n2560 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01123 n2701 p_2_2_d2j n2703 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01122 n2702 p_2_2_d2jbar n2701 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01121 p_2_26_t_s n2701 n2700 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01120 n2701 n2700 p_2_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01119 c_2_26_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01118 vss p_2_26_t_s c_2_26_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01117 n2700 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01116 vss a_25 n2702 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01115 n2703 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01114 c_3_25_cin n2905 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01113 vss c_2_26_a n2903 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01112 n2903 c_2_26_b n2905 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01111 c_2_26_b c_2_26_a c_2_26_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01110 c_2_26_s1_s c_2_26_b c_2_26_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01109 c_3_24_a c_2_26_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_01108 vss n3325 c_2_25_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01107 n2904 c_2_25_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01106 vss c_2_25_a n2904 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01105 n3325 p_16_1_c2j n2904 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01104 n2902 c_2_25_b n3325 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01103 vss c_2_25_a n2902 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01102 n3065 p_16_1_c2j c_2_25_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01101 c_2_25_s2_s n3065 p_16_1_c2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01100 c_2_25_a c_2_25_b c_2_25_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01099 c_2_25_s1_s c_2_25_a c_2_25_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01098 c_3_23_a c_2_25_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01097 vss c_2_25_s1_s n3065 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01096 n3334 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01095 vss a_23 n2910 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01094 n2910 p_2_2_d2j n3071 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01093 n3071 p_2_2_d2jbar n2911 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01092 n2911 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01091 vss p_2_25_t_s c_2_25_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01090 c_2_25_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01089 n3071 n3334 p_2_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01088 p_2_25_t_s n3071 n3334 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01087 n3514 p_2_2_d2j n3513 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01086 n3512 p_2_2_d2jbar n3514 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01085 p_2_24_t_s n3514 n3511 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01084 n3514 n3511 p_2_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01083 c_2_24_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01082 vss p_2_24_t_s c_2_24_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01081 n3511 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01080 vss a_23 n3512 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01079 n3513 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01078 c_3_23_cin n3508 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01077 vss c_2_24_a n3507 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01076 n3507 c_2_24_b n3508 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01075 c_2_24_b c_2_24_a c_2_24_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01074 c_2_24_s1_s c_2_24_b c_2_24_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01073 c_3_22_a c_2_24_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_01072 vss n3917 c_2_23_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01071 n3649 c_2_23_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01070 vss c_2_23_a n3649 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01069 n3917 p_15_1_c2j n3649 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01068 n3648 c_2_23_b n3917 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01067 vss c_2_23_a n3648 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01066 n3921 p_15_1_c2j c_2_23_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01065 c_2_23_s2_s n3921 p_15_1_c2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01064 c_2_23_a c_2_23_b c_2_23_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01063 c_2_23_s1_s c_2_23_a c_2_23_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01062 c_3_21_a c_2_23_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01061 vss c_2_23_s1_s n3921 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01060 n3925 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01059 vss a_21 n3652 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01058 n3652 p_2_2_d2j n3930 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01057 n3930 p_2_2_d2jbar n3653 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01056 n3653 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01055 vss p_2_23_t_s c_2_23_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01054 c_2_23_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01053 n3930 n3925 p_2_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01052 p_2_23_t_s n3930 n3925 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01051 n4333 p_2_2_d2j n4332 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01050 n4331 p_2_2_d2jbar n4333 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01049 p_2_22_t_s n4333 n4329 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01048 n4333 n4329 p_2_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01047 c_2_22_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01046 vss p_2_22_t_s c_2_22_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01045 n4329 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01044 vss a_21 n4331 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01043 n4332 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01042 c_3_21_cin n4325 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01041 vss c_2_22_a n4324 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01040 n4324 c_2_22_b n4325 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01039 c_2_22_b c_2_22_a c_2_22_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01038 c_2_22_s1_s c_2_22_b c_2_22_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01037 c_3_20_a c_2_22_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_01036 vss n4702 c_2_21_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01035 n4413 p_2_21_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01034 vss c_2_21_a n4413 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01033 n4702 p_14_1_c2j n4413 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01032 n4412 p_2_21_pi2j n4702 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01031 vss c_2_21_a n4412 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01030 n4705 p_14_1_c2j c_2_21_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01029 c_2_21_s2_s n4705 p_14_1_c2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01028 c_2_21_a p_2_21_pi2j c_2_21_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01027 c_2_21_s1_s c_2_21_a p_2_21_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01026 c_3_19_a c_2_21_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01025 vss c_2_21_s1_s n4705 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01024 n4710 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01023 vss a_19 n4414 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01022 n4414 p_2_2_d2j n4715 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01021 n4715 p_2_2_d2jbar n4415 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01020 n4415 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01019 vss p_2_21_t_s p_2_21_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01018 p_2_21_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01017 n4715 n4710 p_2_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01016 p_2_21_t_s n4715 n4710 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01015 n5078 p_2_2_d2j n5079 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01014 n5077 p_2_2_d2jbar n5078 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01013 p_2_20_t_s n5078 n5075 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01012 n5078 n5075 p_2_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01011 p_2_20_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01010 vss p_2_20_t_s p_2_20_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_01009 n5075 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01008 vss a_19 n5077 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01007 n5079 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01006 c_3_19_cin n5071 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01005 vss c_2_20_a n5070 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01004 n5070 p_2_20_pi2j n5071 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01003 p_2_20_pi2j c_2_20_a c_2_20_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01002 c_2_20_s1_s p_2_20_pi2j c_2_20_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01001 c_3_18_a c_2_20_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_01000 vss n5467 c_2_19_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00999 n5154 p_2_19_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00998 vss c_2_19_a n5154 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00997 n5467 p_12_1_c2j n5154 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00996 n5153 p_2_19_pi2j n5467 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00995 vss c_2_19_a n5153 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00994 n5472 p_12_1_c2j c_2_19_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00993 c_2_19_s2_s n5472 p_12_1_c2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00992 c_2_19_a p_2_19_pi2j c_2_19_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00991 c_2_19_s1_s c_2_19_a p_2_19_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00990 c_3_17_a c_2_19_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00989 vss c_2_19_s1_s n5472 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00988 n5478 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00987 vss a_17 n5155 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00986 n5155 p_2_2_d2j n5481 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00985 n5481 p_2_2_d2jbar n5156 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00984 n5156 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00983 vss p_2_19_t_s p_2_19_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00982 p_2_19_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00981 n5481 n5478 p_2_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00980 p_2_19_t_s n5481 n5478 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00979 n5833 p_2_2_d2j n5831 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00978 n5832 p_2_2_d2jbar n5833 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00977 p_2_18_t_s n5833 n5830 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00976 n5833 n5830 p_2_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00975 p_2_18_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00974 vss p_2_18_t_s p_2_18_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00973 n5830 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00972 vss a_17 n5832 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00971 n5831 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00970 c_3_17_cin n5825 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00969 vss c_2_18_a n5824 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00968 n5824 p_2_18_pi2j n5825 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00967 p_2_18_pi2j c_2_18_a c_2_18_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00966 c_2_18_s1_s p_2_18_pi2j c_2_18_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00965 c_3_16_a c_2_18_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_00964 vss n6268 c_2_17_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00963 n5927 p_2_17_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00962 vss c_2_17_a n5927 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00961 n6268 p_11_1_c2j n5927 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00960 n5823 p_2_17_pi2j n6268 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00959 vss c_2_17_a n5823 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00958 n6265 p_11_1_c2j c_2_17_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00957 c_2_17_s2_s n6265 p_11_1_c2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00956 c_2_17_a p_2_17_pi2j c_2_17_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00955 c_2_17_s1_s c_2_17_a p_2_17_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00954 c_3_15_a c_2_17_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00953 vss c_2_17_s1_s n6265 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00952 n6277 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00951 vss a_15 n5931 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00950 n5931 p_2_2_d2j n6278 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00949 n6278 p_2_2_d2jbar n5930 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00948 n5930 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00947 vss p_2_17_t_s p_2_17_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00946 p_2_17_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00945 n6278 n6277 p_2_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00944 p_2_17_t_s n6278 n6277 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00943 n6397 p_2_2_d2j n6399 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00942 n6398 p_2_2_d2jbar n6397 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00941 p_2_16_t_s n6397 n6609 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00940 n6397 n6609 p_2_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00939 p_2_16_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00938 vss p_2_16_t_s p_2_16_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00937 n6609 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00936 vss a_15 n6398 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00935 n6399 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00934 c_3_15_cin n6604 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00933 vss c_2_16_a n6602 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00932 n6602 p_2_16_pi2j n6604 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00931 p_2_16_pi2j c_2_16_a c_2_16_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00930 c_2_16_s1_s p_2_16_pi2j c_2_16_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00929 c_3_14_a c_2_16_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_00928 vss n7028 c_2_15_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00927 n6603 c_2_15_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00926 vss c_2_15_a n6603 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00925 n7028 p_10_1_c2j n6603 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00924 n6601 c_2_15_b n7028 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00923 vss c_2_15_a n6601 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00922 n6766 p_10_1_c2j c_2_15_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00921 c_2_15_s2_s n6766 p_10_1_c2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00920 c_2_15_a c_2_15_b c_2_15_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00919 c_2_15_s1_s c_2_15_a c_2_15_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00918 c_3_13_a c_2_15_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00917 vss c_2_15_s1_s n6766 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00916 n7036 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00915 vss a_13 n6611 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00914 n6611 p_2_2_d2j n6772 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00913 n6772 p_2_2_d2jbar n6610 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00912 n6610 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00911 vss p_2_15_t_s c_2_15_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00910 c_2_15_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00909 n6772 n7036 p_2_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00908 p_2_15_t_s n6772 n7036 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00907 n7208 p_2_2_d2j n7207 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00906 n7206 p_2_2_d2jbar n7208 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00905 p_2_14_t_s n7208 n7205 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00904 n7208 n7205 p_2_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00903 p_2_14_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00902 vss p_2_14_t_s p_2_14_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00901 n7205 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00900 vss a_13 n7206 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00899 n7207 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00898 c_3_13_cin n7202 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00897 vss c_2_14_a n7201 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00896 n7201 p_2_14_pi2j n7202 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00895 p_2_14_pi2j c_2_14_a c_2_14_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00894 c_2_14_s1_s p_2_14_pi2j c_2_14_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00893 c_3_12_a c_2_14_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_00892 vss n7578 c_2_13_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00891 n7359 c_2_13_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00890 vss c_2_13_a n7359 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00889 n7578 p_9_1_c2j n7359 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00888 n7358 c_2_13_b n7578 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00887 vss c_2_13_a n7358 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00886 n7582 p_9_1_c2j c_2_13_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00885 c_2_13_s2_s n7582 p_9_1_c2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00884 c_2_13_a c_2_13_b c_2_13_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00883 c_2_13_s1_s c_2_13_a c_2_13_b vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00882 c_3_11_a c_2_13_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00881 vss c_2_13_s1_s n7582 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00880 n7585 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00879 vss a_11 n7362 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00878 n7362 p_2_2_d2j n7589 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00877 n7589 p_2_2_d2jbar n7363 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00876 n7363 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00875 vss p_2_13_t_s c_2_13_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00874 c_2_13_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00873 n7589 n7585 p_2_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00872 p_2_13_t_s n7589 n7585 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00871 n8012 p_2_2_d2j n8011 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00870 n8010 p_2_2_d2jbar n8012 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00869 p_2_12_t_s n8012 n8008 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00868 n8012 n8008 p_2_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00867 c_2_12_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00866 vss p_2_12_t_s c_2_12_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00865 n8008 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00864 vss a_11 n8010 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00863 n8011 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00862 c_3_11_cin n8005 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00861 vss c_2_12_a n8004 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00860 n8004 c_2_12_b n8005 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00859 c_2_12_b c_2_12_a c_2_12_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00858 c_2_12_s1_s c_2_12_b c_2_12_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00857 c_3_10_a c_2_12_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_00856 vss n8390 c_2_11_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00855 n8103 p_2_11_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00854 vss c_2_11_a n8103 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00853 n8390 p_8_1_c2j n8103 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00852 n8102 p_2_11_pi2j n8390 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00851 vss c_2_11_a n8102 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00850 n8394 p_8_1_c2j c_2_11_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00849 c_2_11_s2_s n8394 p_8_1_c2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00848 c_2_11_a p_2_11_pi2j c_2_11_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00847 c_2_11_s1_s c_2_11_a p_2_11_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00846 c_3_9_a c_2_11_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00845 vss c_2_11_s1_s n8394 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00844 n8398 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00843 vss a_9 n8105 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00842 n8105 p_2_2_d2j n8403 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00841 n8403 p_2_2_d2jbar n8106 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00840 n8106 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00839 vss p_2_11_t_s p_2_11_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00838 p_2_11_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00837 n8403 n8398 p_2_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00836 p_2_11_t_s n8403 n8398 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00835 n8767 p_2_2_d2j n8768 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00834 n8766 p_2_2_d2jbar n8767 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00833 p_2_10_t_s n8767 n8764 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00832 n8767 n8764 p_2_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00831 p_2_10_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00830 vss p_2_10_t_s p_2_10_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00829 n8764 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00828 vss a_9 n8766 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00827 n8768 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00826 c_3_9_cin n8760 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00825 vss c_2_10_a n8759 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00824 n8759 p_2_10_pi2j n8760 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00823 p_2_10_pi2j c_2_10_a c_2_10_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00822 c_2_10_s1_s p_2_10_pi2j c_2_10_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00821 c_3_8_a c_2_10_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00820 vss n9155 c_2_9_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00819 n8846 p_2_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00818 vss c_2_9_a n8846 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00817 n9155 p_6_1_c2j n8846 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00816 n8845 p_2_9_pi2j n9155 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00815 vss c_2_9_a n8845 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00814 n9160 p_6_1_c2j c_2_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00813 c_2_9_s2_s n9160 p_6_1_c2j vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00812 c_2_9_a p_2_9_pi2j c_2_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00811 c_2_9_s1_s c_2_9_a p_2_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00810 c_3_7_a c_2_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00809 vss c_2_9_s1_s n9160 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00808 n9166 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00807 vss a_7 n8847 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00806 n8847 p_2_2_d2j n9169 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00805 n9169 p_2_2_d2jbar n8848 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00804 n8848 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00803 vss p_2_9_t_s p_2_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00802 p_2_9_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00801 n9169 n9166 p_2_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00800 p_2_9_t_s n9169 n9166 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00799 n9514 p_2_2_d2j n9512 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00798 n9513 p_2_2_d2jbar n9514 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00797 p_2_8_t_s n9514 n9511 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00796 n9514 n9511 p_2_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00795 p_2_8_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00794 vss p_2_8_t_s p_2_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00793 n9511 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00792 vss a_7 n9513 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00791 n9512 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00790 c_3_7_cin n9506 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00789 vss c_2_8_a n9505 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00788 n9505 p_2_8_pi2j n9506 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00787 p_2_8_pi2j c_2_8_a c_2_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00786 c_2_8_s1_s p_2_8_pi2j c_2_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00785 c_3_6_a c_2_8_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00784 vss n9949 c_2_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00783 n9605 p_2_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00782 vss c_2_7_a n9605 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00781 n9949 p_5_1_c2j n9605 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00780 n9504 p_2_7_pi2j n9949 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00779 vss c_2_7_a n9504 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00778 n9957 p_5_1_c2j c_2_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00777 c_2_7_s2_s n9957 p_5_1_c2j vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00776 c_2_7_a p_2_7_pi2j c_2_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00775 c_2_7_s1_s c_2_7_a p_2_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00774 c_3_5_a c_2_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00773 vss c_2_7_s1_s n9957 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00772 n9962 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00771 vss a_5 n9609 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00770 n9609 p_2_2_d2j n9961 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00769 n9961 p_2_2_d2jbar n9608 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00768 n9608 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00767 vss p_2_7_t_s p_2_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00766 p_2_7_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00765 n9961 n9962 p_2_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00764 p_2_7_t_s n9961 n9962 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00763 n10283 p_2_2_d2j n10056 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00762 n10055 p_2_2_d2jbar n10283 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00761 p_2_6_t_s n10283 n10284 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00760 n10283 n10284 p_2_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00759 p_2_6_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00758 vss p_2_6_t_s p_2_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00757 n10284 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00756 vss a_5 n10055 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00755 n10056 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00754 c_3_5_cin n10278 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00753 vss c_2_6_a n10277 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00752 n10277 p_2_6_pi2j n10278 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00751 p_2_6_pi2j c_2_6_a c_2_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00750 c_2_6_s1_s p_2_6_pi2j c_2_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00749 c_3_4_a c_2_6_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00748 vss n10708 c_2_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00747 n10438 c_2_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00746 vss c_2_5_a n10438 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00745 n10708 p_4_1_c2j n10438 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00744 n10276 c_2_5_b n10708 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00743 vss c_2_5_a n10276 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00742 n10441 p_4_1_c2j c_2_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00741 c_2_5_s2_s n10441 p_4_1_c2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00740 c_2_5_a c_2_5_b c_2_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00739 c_2_5_s1_s c_2_5_a c_2_5_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00738 c_3_3_a c_2_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00737 vss c_2_5_s1_s n10441 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00736 n10716 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00735 vss a_3 n10286 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00734 n10286 p_2_2_d2j n10715 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00733 n10715 p_2_2_d2jbar n10285 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00732 n10285 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00731 vss p_2_5_t_s c_2_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00730 c_2_5_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00729 n10715 n10716 p_2_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00728 p_2_5_t_s n10715 n10716 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00727 n10879 p_2_2_d2j n10878 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00726 n10877 p_2_2_d2jbar n10879 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00725 p_2_4_t_s n10879 n10876 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00724 n10879 n10876 p_2_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00723 p_2_4_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00722 vss p_2_4_t_s p_2_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00721 n10876 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00720 vss a_3 n10877 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00719 n10878 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00718 c_3_3_cin n11026 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00717 vss c_2_4_a n10875 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00716 n10875 p_2_4_pi2j n11026 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00715 p_2_4_pi2j c_2_4_a c_2_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00714 c_2_4_s1_s p_2_4_pi2j c_2_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00713 c_3_2_a c_2_4_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00712 vss n11243 c_2_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00711 n11029 c_2_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00710 vss c_2_3_a n11029 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00709 n11243 p_3_1_c2j n11029 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00708 n11028 c_2_3_b n11243 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00707 vss c_2_3_a n11028 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00706 n11247 p_3_1_c2j c_2_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00705 c_2_3_s2_s n11247 p_3_1_c2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00704 c_2_3_a c_2_3_b c_2_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00703 c_2_3_s1_s c_2_3_a c_2_3_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00702 c_3_1_a c_2_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00701 vss c_2_3_s1_s n11247 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00700 n11250 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00699 vss a_1 n11033 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00698 n11033 p_2_2_d2j n11254 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00697 n11254 p_2_2_d2jbar n11034 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00696 n11034 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00695 vss p_2_3_t_s c_2_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00694 c_2_3_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00693 n11254 n11250 p_2_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00692 p_2_3_t_s n11254 n11250 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00691 n11675 p_2_2_d2j n11674 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00690 n11673 p_2_2_d2jbar n11675 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00689 p_2_2_t_s n11675 n11671 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00688 n11675 n11671 p_2_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00687 c_2_2_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00686 vss p_2_2_t_s c_2_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00685 n11671 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00684 vss a_1 n11673 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00683 n11674 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00682 c_3_1_cin n11668 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00681 vss c_2_2_a n11667 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00680 n11667 c_2_2_b n11668 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00679 c_2_2_b c_2_2_a c_2_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00678 c_2_2_s1_s c_2_2_b c_2_2_a vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00677 c_2_2_sum c_2_2_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_00676 vss n12056 c_2_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00675 n11765 p_2_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00674 vss c_2_1_a n11765 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00673 n12056 n12067 n11765 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00672 n11764 p_2_1_pi2j n12056 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00671 vss c_2_1_a n11764 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00670 n12064 n12067 c_2_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00669 c_2_1_s2_s n12064 n12067 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00668 c_2_1_a p_2_1_pi2j c_2_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00667 c_2_1_s1_s c_2_1_a p_2_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00666 c_2_1_sum c_2_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00665 vss c_2_1_s1_s n12064 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00664 p_2_1_t_s n12073 n12069 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00663 n12073 n12069 p_2_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00662 p_2_1_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00661 vss p_2_1_t_s p_2_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00660 n11768 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00659 n12073 p_2_2_d2jbar n11768 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00658 n12069 n12067 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00657 cl4_2_s1_s p_1_2_c2j n12416 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00656 p_1_2_c2j n12416 cl4_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00655 vss cl4_2_s1_s p_0 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00654 vss n12416 n12412 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00653 n12412 p_1_2_c2j n12410 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00652 n12411 n12410 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00651 vss p_1_2_pi2j n12409 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00650 n12408 n12416 n12407 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00649 n12409 p_1_2_c2j n12408 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00648 n12406 n12407 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00647 cl4_2_s3_s p_1_2_pi2j n12411 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00646 p_1_2_pi2j n12411 cl4_2_s3_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00645 vss cl4_2_s3_s p_1 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00644 vss p_1_33_t_s c_2_31_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00643 c_2_31_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00642 p_1_33_a n261 p_1_33_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00641 p_1_33_t_s p_1_33_a n261 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00640 n261 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00639 p_1_33_a a_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00638 vss d_0_n2j c_2_30_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00637 p_1_32_t_s n595 n592 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00636 vss a_31 n593 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00635 n595 d_0_d2j n594 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00634 n594 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00633 c_2_30_a p_1_32_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00632 n595 n592 p_1_32_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00631 n592 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00630 n593 d_0_d2jbar n595 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00629 p_1_31_a d_0_d2jbar n665 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00628 n666 d_0_d2j p_1_31_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00627 vss a_29 n666 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00626 n973 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00625 p_1_31_t_s p_1_31_a n973 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00624 p_1_31_a n973 p_1_31_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00623 c_2_29_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00622 vss p_1_31_t_s c_2_29_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00621 n665 a_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00620 vss d_0_n2j c_2_28_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00619 p_1_30_t_s n1362 n1359 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00618 vss a_29 n1360 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00617 n1362 d_0_d2j n1361 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00616 n1361 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00615 c_2_28_a p_1_30_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00614 n1362 n1359 p_1_30_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00613 n1359 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00612 n1360 d_0_d2jbar n1362 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00611 p_1_29_a d_0_d2jbar n1424 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00610 n1425 d_0_d2j p_1_29_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00609 vss a_27 n1425 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00608 n1759 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00607 p_1_29_t_s p_1_29_a n1759 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00606 p_1_29_a n1759 p_1_29_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00605 n2555 d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00604 vss p_1_29_t_s n2555 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00603 n1424 a_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00602 vss d_0_n2j c_2_26_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00601 p_1_28_t_s n2112 n2110 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00600 vss a_27 n2111 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00599 n2112 d_0_d2j n2113 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00598 n2113 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00597 c_2_26_a p_1_28_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00596 n2112 n2110 p_1_28_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00595 n2110 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00594 n2111 d_0_d2jbar n2112 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00593 p_1_27_a d_0_d2jbar n2242 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00592 n2243 d_0_d2j p_1_27_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00591 vss a_25 n2243 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00590 n2568 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00589 p_1_27_t_s p_1_27_a n2568 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00588 p_1_27_a n2568 p_1_27_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00587 c_2_25_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00586 vss p_1_27_t_s c_2_25_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00585 n2242 a_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00584 vss d_0_n2j c_2_24_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00583 p_1_26_t_s n2707 n2704 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00582 vss a_25 n2705 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00581 n2707 d_0_d2j n2706 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00580 n2706 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00579 c_2_24_a p_1_26_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00578 n2707 n2704 p_1_26_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00577 n2704 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00576 n2705 d_0_d2jbar n2707 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00575 p_1_25_a d_0_d2jbar n2913 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00574 n2914 d_0_d2j p_1_25_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00573 vss a_23 n2914 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00572 n3338 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00571 p_1_25_t_s p_1_25_a n3338 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00570 p_1_25_a n3338 p_1_25_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00569 c_2_23_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00568 vss p_1_25_t_s c_2_23_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00567 n2913 a_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00566 vss d_0_n2j c_2_22_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00565 p_1_24_t_s n3518 n3515 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00564 vss a_23 n3516 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00563 n3518 d_0_d2j n3517 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00562 n3517 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00561 c_2_22_a p_1_24_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00560 n3518 n3515 p_1_24_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00559 n3515 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00558 n3516 d_0_d2jbar n3518 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00557 p_1_23_a d_0_d2jbar n3655 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00556 n3656 d_0_d2j p_1_23_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00555 vss a_21 n3656 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00554 n3935 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00553 p_1_23_t_s p_1_23_a n3935 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00552 p_1_23_a n3935 p_1_23_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00551 c_2_21_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00550 vss p_1_23_t_s c_2_21_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00549 n3655 a_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00548 vss d_0_n2j c_2_20_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00547 p_1_22_t_s n4338 n4335 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00546 vss a_21 n4336 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00545 n4338 d_0_d2j n4337 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00544 n4337 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00543 c_2_20_a p_1_22_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00542 n4338 n4335 p_1_22_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00541 n4335 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00540 n4336 d_0_d2jbar n4338 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00539 p_1_21_a d_0_d2jbar n4416 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00538 n4417 d_0_d2j p_1_21_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00537 vss a_19 n4417 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00536 n4720 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00535 p_1_21_t_s p_1_21_a n4720 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00534 p_1_21_a n4720 p_1_21_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00533 c_2_19_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00532 vss p_1_21_t_s c_2_19_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00531 n4416 a_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00530 vss d_0_n2j c_2_18_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00529 p_1_20_t_s n5084 n5081 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00528 vss a_19 n5082 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00527 n5084 d_0_d2j n5083 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00526 n5083 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00525 c_2_18_a p_1_20_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00524 n5084 n5081 p_1_20_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00523 n5081 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00522 n5082 d_0_d2jbar n5084 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00521 p_1_19_a d_0_d2jbar n5157 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00520 n5158 d_0_d2j p_1_19_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00519 vss a_17 n5158 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00518 n5486 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00517 p_1_19_t_s p_1_19_a n5486 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00516 p_1_19_a n5486 p_1_19_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00515 c_2_17_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00514 vss p_1_19_t_s c_2_17_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00513 n5157 a_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00512 vss d_0_n2j c_2_16_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00511 p_1_18_t_s n5836 n5838 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00510 vss a_17 n5839 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00509 n5836 d_0_d2j n5837 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00508 n5837 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00507 c_2_16_a p_1_18_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00506 n5836 n5838 p_1_18_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00505 n5838 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00504 n5839 d_0_d2jbar n5836 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00503 p_1_17_a d_0_d2jbar n5935 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00502 n5934 d_0_d2j p_1_17_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00501 vss a_15 n5934 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00500 n6286 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00499 p_1_17_t_s p_1_17_a n6286 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00498 p_1_17_a n6286 p_1_17_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00497 c_2_15_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00496 vss p_1_17_t_s c_2_15_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00495 n5935 a_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00494 vss d_0_n2j c_2_14_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00493 p_1_16_t_s n6402 n6613 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00492 vss a_15 n6400 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00491 n6402 d_0_d2j n6401 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00490 n6401 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00489 c_2_14_a p_1_16_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00488 n6402 n6613 p_1_16_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00487 n6613 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00486 n6400 d_0_d2jbar n6402 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00485 p_1_15_a d_0_d2jbar n6614 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00484 n6615 d_0_d2j p_1_15_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00483 vss a_13 n6615 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00482 n7040 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00481 p_1_15_t_s p_1_15_a n7040 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00480 p_1_15_a n7040 p_1_15_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00479 c_2_13_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00478 vss p_1_15_t_s c_2_13_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00477 n6614 a_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00476 vss d_0_n2j c_2_12_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00475 p_1_14_t_s n7212 n7209 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00474 vss a_13 n7210 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00473 n7212 d_0_d2j n7211 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00472 n7211 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00471 c_2_12_a p_1_14_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00470 n7212 n7209 p_1_14_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00469 n7209 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00468 n7210 d_0_d2jbar n7212 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00467 p_1_13_a d_0_d2jbar n7365 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00466 n7366 d_0_d2j p_1_13_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00465 vss a_11 n7366 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00464 n7801 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00463 p_1_13_t_s p_1_13_a n7801 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00462 p_1_13_a n7801 p_1_13_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00461 c_2_11_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00460 vss p_1_13_t_s c_2_11_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00459 n7365 a_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00458 vss d_0_n2j c_2_10_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00457 p_1_12_t_s n8017 n8014 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00456 vss a_11 n8015 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00455 n8017 d_0_d2j n8016 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00454 n8016 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00453 c_2_10_a p_1_12_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00452 n8017 n8014 p_1_12_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00451 n8014 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00450 n8015 d_0_d2jbar n8017 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00449 p_1_11_a d_0_d2jbar n8107 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00448 n8108 d_0_d2j p_1_11_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00447 vss a_9 n8108 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00446 n8408 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00445 p_1_11_t_s p_1_11_a n8408 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00444 p_1_11_a n8408 p_1_11_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00443 c_2_9_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00442 vss p_1_11_t_s c_2_9_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00441 n8107 a_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00440 vss d_0_n2j c_2_8_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00439 p_1_10_t_s n8773 n8770 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00438 vss a_9 n8771 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00437 n8773 d_0_d2j n8772 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00436 n8772 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00435 c_2_8_a p_1_10_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00434 n8773 n8770 p_1_10_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00433 n8770 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00432 n8771 d_0_d2jbar n8773 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00431 p_1_9_a d_0_d2jbar n8849 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00430 n8850 d_0_d2j p_1_9_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00429 vss a_7 n8850 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00428 n9174 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00427 p_1_9_t_s p_1_9_a n9174 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00426 p_1_9_a n9174 p_1_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00425 c_2_7_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00424 vss p_1_9_t_s c_2_7_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00423 n8849 a_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00422 vss d_0_n2j c_2_6_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00421 p_1_8_t_s n9517 n9519 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00420 vss a_7 n9520 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00419 n9517 d_0_d2j n9518 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00418 n9518 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00417 c_2_6_a p_1_8_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00416 n9517 n9519 p_1_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00415 n9519 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00414 n9520 d_0_d2jbar n9517 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00413 p_1_7_a d_0_d2jbar n9612 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00412 n9613 d_0_d2j p_1_7_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00411 vss a_5 n9613 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00410 n9969 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00409 p_1_7_t_s p_1_7_a n9969 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00408 p_1_7_a n9969 p_1_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00407 c_2_5_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00406 vss p_1_7_t_s c_2_5_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00405 n9612 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00404 vss d_0_n2j c_2_4_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00403 p_1_6_t_s n10287 n10289 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00402 vss a_5 n10057 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00401 n10287 d_0_d2j n10058 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00400 n10058 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00399 c_2_4_a p_1_6_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00398 n10287 n10289 p_1_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00397 n10289 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00396 n10057 d_0_d2jbar n10287 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00395 p_1_5_a d_0_d2jbar n10291 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00394 n10292 d_0_d2j p_1_5_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00393 vss a_3 n10292 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00392 n10722 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00391 p_1_5_t_s p_1_5_a n10722 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00390 p_1_5_a n10722 p_1_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00389 c_2_3_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00388 vss p_1_5_t_s c_2_3_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00387 n10291 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00386 vss d_0_n2j c_2_2_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00385 p_1_4_t_s n10883 n10880 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00384 vss a_3 n10881 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00383 n10883 d_0_d2j n10882 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00382 n10882 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00381 c_2_2_a p_1_4_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00380 n10883 n10880 p_1_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00379 n10880 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00378 n10881 d_0_d2jbar n10883 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00377 p_1_3_a d_0_d2jbar n11036 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00376 n11037 d_0_d2j p_1_3_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00375 vss a_1 n11037 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00374 n11466 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00373 p_1_3_t_s p_1_3_a n11466 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00372 p_1_3_a n11466 p_1_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00371 c_2_1_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00370 vss p_1_3_t_s c_2_1_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00369 n11036 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00368 vss d_0_n2j p_1_2_pi2j vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00367 p_1_2_t_s n11680 n11677 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00366 vss a_1 n11678 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00365 n11680 d_0_d2j n11679 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00364 n11679 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00363 p_1_2_pi2j p_1_2_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00362 n11680 n11677 p_1_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00361 n11677 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00360 n11678 d_0_d2jbar n11680 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00359 n11769 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00358 vss p_1_1_t_s n12416 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00357 n12416 d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00356 n12077 n12076 p_1_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00355 p_1_1_t_s n12077 n12076 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00354 n12076 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00353 n12077 d_0_d2jbar n11769 vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00352 vss n978 p_18_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00351 p_18_1_c2j n976 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00350 vss n1367 n667 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00349 n667 n1373 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00348 n976 b_31 n667 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00347 vss n1366 n669 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00346 n669 n1373 n670 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00345 n670 n1367 n978 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00344 n978 b_29 n671 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00343 n671 b_30 n668 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00342 n668 b_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00341 p_18_2_d2j n1370 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00340 vss p_18_2_d2j p_18_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00339 n1364 n1366 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00338 n1366 b_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00337 vss b_31 n1365 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00336 n1365 n1367 n1371 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00335 n1367 b_29 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00334 n1364 b_29 n1372 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00333 n1373 b_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00332 n1371 n1373 n1370 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00331 n1370 b_30 n1372 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00330 vss n1766 p_17_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00329 p_17_1_c2j n1764 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00328 vss n2118 n1426 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00327 n1426 n2121 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00326 n1764 b_29 n1426 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00325 vss n2114 n1428 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00324 n1428 n2121 n1429 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00323 n1429 n2118 n1766 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00322 n1766 b_27 n1430 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00321 n1430 b_28 n1427 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00320 n1427 b_29 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00319 p_17_2_d2j n2128 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00318 vss p_17_2_d2j p_17_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00317 n2117 n2114 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00316 n2114 b_29 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00315 vss b_29 n2119 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00314 n2119 n2118 n2126 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00313 n2118 b_27 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00312 n2117 b_27 n2127 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00311 n2121 b_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00310 n2126 n2121 n2128 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00309 n2128 b_28 n2127 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00308 vss n2578 p_16_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00307 p_16_1_c2j n2576 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00306 vss n2917 n2116 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00305 n2116 n2921 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00304 n2576 b_27 n2116 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00303 vss n2915 n2125 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00302 n2125 n2921 n2124 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00301 n2124 n2917 n2578 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00300 n2578 b_25 n2122 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00299 n2122 b_26 n2123 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00298 n2123 b_27 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00297 p_16_2_d2j n2927 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00296 vss p_16_2_d2j p_16_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00295 n2919 n2915 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00294 n2915 b_27 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00293 vss b_27 n2920 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00292 n2920 n2917 n2928 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00291 n2917 b_25 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00290 n2919 b_25 n2929 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00289 n2921 b_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00288 n2928 n2921 n2927 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00287 n2927 b_26 n2929 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00286 vss n3080 p_15_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00285 p_15_1_c2j n3078 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00284 vss n3657 n2918 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00283 n2918 n3660 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00282 n3078 b_25 n2918 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00281 vss n3521 n2925 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00280 n2925 n3660 n2926 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00279 n2926 n3657 n3080 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00278 n3080 b_23 n2924 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00277 n2924 b_24 n2923 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00276 n2923 b_25 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00275 p_15_2_d2j n3668 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00274 vss p_15_2_d2j p_15_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00273 n3659 n3521 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00272 n3521 b_25 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00271 vss b_25 n3520 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00270 n3520 n3657 n3666 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00269 n3657 b_23 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00268 n3659 b_23 n3667 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00267 n3660 b_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00266 n3666 n3660 n3668 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00265 n3668 b_24 n3667 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00264 vss n3941 p_14_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00263 p_14_1_c2j n3938 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00262 vss n4344 n3658 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00261 n3658 n4349 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00260 n3938 b_23 n3658 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00259 vss n4342 n3663 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00258 n3663 n4349 n3664 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00257 n3664 n4344 n3941 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00256 n3941 b_21 n3665 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00255 n3665 b_22 n3662 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00254 n3662 b_23 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00253 p_14_2_d2j n4346 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00252 vss p_14_2_d2j p_14_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00251 n4340 n4342 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00250 n4342 b_23 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00249 vss b_23 n4341 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00248 n4341 n4344 n4347 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00247 n4344 b_21 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00246 n4340 b_21 n4348 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00245 n4349 b_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00244 n4347 n4349 n4346 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00243 n4346 b_22 n4348 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00242 vss n4725 p_12_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00241 p_12_1_c2j n4723 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00240 vss n5089 n4418 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00239 n4418 n5092 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00238 n4723 b_21 n4418 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00237 vss n5088 n4420 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00236 n4420 n5092 n4421 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00235 n4421 n5089 n4725 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00234 n4725 b_19 n4422 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00233 n4422 b_20 n4419 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00232 n4419 b_21 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00231 p_12_2_d2j n5093 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00230 vss p_12_2_d2j p_12_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00229 n5086 n5088 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00228 n5088 b_21 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00227 vss b_21 n5087 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00226 n5087 n5089 n5095 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00225 n5089 b_19 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00224 n5086 b_19 n5094 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00223 n5092 b_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00222 n5095 n5092 n5093 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00221 n5093 b_20 n5094 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00220 vss n5493 p_11_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00219 p_11_1_c2j n5491 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00218 vss n5844 n5159 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00217 n5159 n5846 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00216 n5491 b_19 n5159 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00215 vss n5840 n5161 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00214 n5161 n5846 n5162 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00213 n5162 n5844 n5493 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00212 n5493 b_17 n5163 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00211 n5163 b_18 n5160 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00210 n5160 b_19 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00209 p_11_2_d2j n5854 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00208 vss p_11_2_d2j p_11_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00207 n5843 n5840 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00206 n5840 b_19 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00205 vss b_19 n5845 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00204 n5845 n5844 n5852 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00203 n5844 b_17 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00202 n5843 b_17 n5853 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00201 n5846 b_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00200 n5852 n5846 n5854 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00199 n5854 b_18 n5853 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00198 vss n6296 p_10_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00197 p_10_1_c2j n6294 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00196 vss n6618 n5842 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00195 n5842 n6623 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00194 n6294 b_17 n5842 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00193 vss n6616 n5851 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00192 n5851 n6623 n5850 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00191 n5850 n6618 n6296 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00190 n6296 b_15 n5848 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00189 n5848 b_16 n5849 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00188 n5849 b_17 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00187 p_10_2_d2j n6628 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00186 vss p_10_2_d2j p_10_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00185 n6620 n6616 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00184 n6616 b_17 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00183 vss b_17 n6621 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00182 n6621 n6618 n6629 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00181 n6618 b_15 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00180 n6620 b_15 n6630 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00179 n6623 b_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00178 n6629 n6623 n6628 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00177 n6628 b_16 n6630 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00176 vss n7048 p_9_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00175 p_9_1_c2j n7046 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00174 vss n7367 n6619 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00173 n6619 n7371 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00172 n7046 b_15 n6619 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00171 vss n7214 n6626 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00170 n6626 n7371 n6627 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00169 n6627 n7367 n7048 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00168 n7048 b_13 n6625 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00167 n6625 b_14 n6624 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00166 n6624 b_15 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00165 p_9_2_d2j n7377 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00164 vss p_9_2_d2j p_9_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00163 n7369 n7214 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00162 n7214 b_15 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00161 vss b_15 n7370 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00160 n7370 n7367 n7378 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00159 n7367 b_13 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00158 n7369 b_13 n7379 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00157 n7371 b_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00156 n7378 n7371 n7377 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00155 n7377 b_14 n7379 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00154 vss n7598 p_8_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00153 p_8_1_c2j n7596 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00152 vss n8023 n7368 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00151 n7368 n8027 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00150 n7596 b_13 n7368 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00149 vss n8020 n7375 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00148 n7375 n8027 n7376 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00147 n7376 n8023 n7598 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00146 n7598 b_11 n7374 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00145 n7374 b_12 n7373 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00144 n7373 b_13 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00143 p_8_2_d2j n8024 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00142 vss p_8_2_d2j p_8_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00141 n8109 n8020 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00140 n8020 b_13 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00139 vss b_13 n8019 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00138 n8019 n8023 n8025 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00137 n8023 b_11 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00136 n8109 b_11 n8026 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00135 n8027 b_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00134 n8025 n8027 n8024 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00133 n8024 b_12 n8026 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00132 vss n8413 p_6_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00131 p_6_1_c2j n8411 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00130 vss n8775 n8110 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00129 n8110 n8781 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00128 n8411 b_11 n8110 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00127 vss n8778 n8112 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00126 n8112 n8781 n8113 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00125 n8113 n8775 n8413 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00124 n8413 b_9 n8114 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00123 n8114 b_10 n8111 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00122 n8111 b_11 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00121 p_6_2_d2j n8782 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00120 vss p_6_2_d2j p_6_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00119 n8776 n8778 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00118 n8778 b_11 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00117 vss b_11 n8777 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00116 n8777 n8775 n8784 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00115 n8775 b_9 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00114 n8776 b_9 n8783 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00113 n8781 b_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00112 n8784 n8781 n8782 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00111 n8782 b_10 n8783 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00110 vss n9180 p_5_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00109 p_5_1_c2j n9179 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00108 vss n9526 n8851 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00107 n8851 n9528 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00106 n9179 b_9 n8851 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00105 vss n9525 n8853 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00104 n8853 n9528 n8854 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00103 n8854 n9526 n9180 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00102 n9180 b_7 n8855 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00101 n8855 b_8 n8852 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00100 n8852 b_9 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00099 p_5_2_d2j n9529 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00098 vss p_5_2_d2j p_5_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00097 n9523 n9525 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00096 n9525 b_9 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00095 vss b_9 n9524 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00094 n9524 n9526 n9531 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00093 n9526 b_7 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00092 n9523 b_7 n9530 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00091 n9528 b_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00090 n9531 n9528 n9529 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00089 n9529 b_8 n9530 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00088 vss n9981 p_4_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00087 p_4_1_c2j n9979 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00086 vss n10298 n9522 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00085 n9522 n10300 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00084 n9979 b_7 n9522 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00083 vss n10293 n9617 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00082 n9617 n10300 n9616 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00081 n9616 n10298 n9981 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00080 n9981 b_5 n9614 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00079 n9614 b_6 n9615 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00078 n9615 b_7 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00077 p_4_2_d2j n10305 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00076 vss p_4_2_d2j p_4_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00075 n10296 n10293 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00074 n10293 b_7 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00073 vss b_7 n10297 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00072 n10297 n10298 n10306 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00071 n10298 b_5 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00070 n10296 b_5 n10307 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00069 n10300 b_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00068 n10306 n10300 n10305 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00067 n10305 b_6 n10307 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00066 vss n10730 p_3_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00065 p_3_1_c2j n10728 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00064 vss n11038 n10295 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00063 n10295 n11042 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00062 n10728 b_5 n10295 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00061 vss n10885 n10303 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00060 n10303 n11042 n10304 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00059 n10304 n11038 n10730 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00058 n10730 b_3 n10302 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00057 n10302 b_4 n10301 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00056 n10301 b_5 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00055 p_3_2_d2j n11048 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00054 vss p_3_2_d2j p_3_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00053 n11040 n10885 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00052 n10885 b_5 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00051 vss b_5 n11041 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00050 n11041 n11038 n11049 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00049 n11038 b_3 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00048 n11040 b_3 n11050 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00047 n11042 b_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00046 n11049 n11042 n11048 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00045 n11048 b_4 n11050 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00044 vss n11263 p_2_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00043 n12067 n11261 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00042 vss n11685 n11039 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00041 n11039 n11690 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00040 n11261 b_3 n11039 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00039 vss n11683 n11046 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00038 n11046 n11690 n11047 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00037 n11047 n11685 n11263 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00036 n11263 b_1 n11045 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00035 n11045 b_2 n11044 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00034 n11044 b_3 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00033 p_2_2_d2j n11687 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00032 vss p_2_2_d2j p_2_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00031 n11770 n11683 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00030 n11683 b_3 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00029 vss b_3 n11682 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00028 n11682 n11685 n11688 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00027 n11685 b_1 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00026 n11770 b_1 n11689 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00025 n11690 b_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00024 n11688 n11690 n11687 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00023 n11687 b_2 n11689 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00022 n12427 b_0 n12426 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00021 n12428 n12430 n12427 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00020 n12430 b_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00019 n12422 vss n12426 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00018 n12423 vss vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00017 n12424 n12423 n12428 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00016 vss b_1 n12424 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00015 n12421 b_1 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00014 n12422 n12421 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00013 vss d_0_d2j d_0_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00012 d_0_d2j n12427 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00011 n11774 b_1 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00010 n11775 b_0 n11774 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00009 n12083 vss n11775 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00008 n11772 n12423 n12083 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00007 n11773 n12430 n11772 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00006 vss n12421 n11773 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00005 n12080 b_1 n11771 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00004 n11771 n12430 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00003 vss n12423 n11771 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00002 p_1_2_c2j n12080 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00001 vss n12083 d_0_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
.ends ex_m32x32

