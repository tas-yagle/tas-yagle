
.subckt ex_shift32 ext in_d_0 in_d_1 in_d_2 in_d_3 in_d_4 in_d_5 in_d_6 
+ in_d_7 in_d_8 in_d_9 in_d_10 in_d_11 in_d_12 in_d_13 in_d_14 in_d_15 in_d_16 
+ in_d_17 in_d_18 in_d_19 in_d_20 in_d_21 in_d_22 in_d_23 in_d_24 in_d_25 
+ in_d_26 in_d_27 in_d_28 in_d_29 in_d_30 in_d_31 in_s_0 in_s_1 in_s_2 in_s_3 
+ in_s_4 left out_d_0 out_d_1 out_d_2 out_d_3 out_d_4 out_d_5 out_d_6 out_d_7 
+ out_d_8 out_d_9 out_d_10 out_d_11 out_d_12 out_d_13 out_d_14 out_d_15 
+ out_d_16 out_d_17 out_d_18 out_d_19 out_d_20 out_d_21 out_d_22 out_d_23 
+ out_d_24 out_d_25 out_d_26 out_d_27 out_d_28 out_d_29 out_d_30 out_d_31 rot 
+ vdd vss 
Mtr_02828 bsrmux_0_shr bshmat_0_nshr vdd vdd TP L=0.18U W=9.72U AS=3.4992P 
+ AD=3.4992P PS=20.16U PD=20.16U 
Mtr_02827 vdd n5 n3 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02826 n3 bshsel_0_nright vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02825 n12 n3 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02824 vdd n11 bshcmd_0_nasr vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02823 n11 n12 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02822 vdd in_d_31 n11 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02821 n11 ext vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02820 n5 rot vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02819 n9 bshlmx_0_nnleft vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02818 vdd n5 n9 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_02817 bshmat_0_nshr n9 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02816 bshlmx_0_asr bshcmd_0_nasr vdd vdd TP L=0.18U W=9.72U AS=3.4992P 
+ AD=3.4992P PS=20.16U PD=20.16U 
Mtr_02815 vdd n12 bshlmx_0_lsl vdd TP L=0.18U W=9.72U AS=3.4992P AD=3.4992P 
+ PS=20.16U PD=20.16U 
Mtr_02814 bshmatr_0_comr0 bssnbl_15_zero vdd vdd TP L=0.18U W=9.72U AS=3.4992P 
+ AD=3.4992P PS=20.16U PD=20.16U 
Mtr_02813 vdd bshsel_0_nright n699 vdd TP L=0.18U W=9.72U AS=3.4992P 
+ AD=3.4992P PS=20.16U PD=20.16U 
Mtr_02812 n693 bshlmx_0_nnleft vdd vdd TP L=0.18U W=9.72U AS=3.4992P 
+ AD=3.4992P PS=20.16U PD=20.16U 
Mtr_02811 bshsel_0_nright left vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02810 vdd bshsel_0_nright bshlmx_0_nnleft vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_02809 vdd bsm_0_15_out_2_s out_d_30 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02808 vdd bsoout_15_out_1_s out_d_31 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02807 vdd out_d_31 bsoout_15_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02806 vdd out_d_30 bsm_0_15_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02805 vdd bsoout_14_out_2_s out_d_28 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02804 vdd bsoout_14_out_1_s out_d_29 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02803 vdd out_d_29 bsoout_14_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02802 vdd out_d_28 bsoout_14_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02801 vdd bsoout_13_out_2_s out_d_26 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02800 vdd bsoout_13_out_1_s out_d_27 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02799 vdd out_d_27 bsoout_13_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02798 vdd out_d_26 bsoout_13_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02797 vdd bsm_0_12_out_2_s out_d_24 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02796 vdd bsoout_12_out_1_s out_d_25 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02795 vdd out_d_25 bsoout_12_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02794 vdd out_d_24 bsm_0_12_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02793 vdd bsm_0_11_out_2_s out_d_22 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02792 vdd bsoout_11_out_1_s out_d_23 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02791 vdd out_d_23 bsoout_11_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02790 vdd out_d_22 bsm_0_11_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02789 vdd bsm_0_10_out_2_s out_d_20 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02788 vdd bsoout_10_out_1_s out_d_21 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02787 vdd out_d_21 bsoout_10_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02786 vdd out_d_20 bsm_0_10_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02785 vdd bsm_0_9_out_2_s out_d_18 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02784 vdd bsoout_9_out_1_s out_d_19 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02783 vdd out_d_19 bsoout_9_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02782 vdd out_d_18 bsm_0_9_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02781 vdd bsoout_8_out_2_s out_d_16 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02780 vdd bsoout_8_out_1_s out_d_17 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02779 vdd out_d_17 bsoout_8_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02778 vdd out_d_16 bsoout_8_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02777 vdd bsm_0_7_out_2_s out_d_14 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02776 vdd bsoout_7_out_1_s out_d_15 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02775 vdd out_d_15 bsoout_7_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02774 vdd out_d_14 bsm_0_7_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02773 vdd bsm_0_6_out_2_s out_d_12 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02772 vdd bsoout_6_out_1_s out_d_13 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02771 vdd out_d_13 bsoout_6_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02770 vdd out_d_12 bsm_0_6_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02769 vdd bsm_0_5_out_2_s out_d_10 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02768 vdd bsoout_5_out_1_s out_d_11 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02767 vdd out_d_11 bsoout_5_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02766 vdd out_d_10 bsm_0_5_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02765 vdd bsm_0_4_out_2_s out_d_8 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02764 vdd bsoout_4_out_1_s out_d_9 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02763 vdd out_d_9 bsoout_4_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02762 vdd out_d_8 bsm_0_4_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02761 vdd bsoout_3_out_2_s out_d_6 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02760 vdd bsoout_3_out_1_s out_d_7 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02759 vdd out_d_7 bsoout_3_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02758 vdd out_d_6 bsoout_3_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02757 vdd bsm_0_2_out_2_s out_d_4 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02756 vdd bsoout_2_out_1_s out_d_5 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02755 vdd out_d_5 bsoout_2_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02754 vdd out_d_4 bsm_0_2_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02753 vdd bsm_0_1_out_2_s out_d_2 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02752 vdd bsoout_1_out_1_s out_d_3 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02751 vdd out_d_3 bsoout_1_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02750 vdd out_d_2 bsm_0_1_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02749 vdd bsm_0_0_out_2_s out_d_0 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02748 vdd bsoout_0_out_1_s out_d_1 vdd TP L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_02747 vdd out_d_1 bsoout_0_out_1_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02746 vdd out_d_0 bsm_0_0_out_2_s vdd TP L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02745 vdd n38 n681 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02744 n681 n38 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02743 vdd n28 bsrmux_15_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02742 bsrmux_15_f1 n28 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02741 vdd n38 n681 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02740 vdd n36 n38 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02739 n36 in_d_30 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02738 vdd bsrmux_0_shr n36 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02737 vdd n28 bsrmux_15_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02736 vdd n27 n28 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02735 n27 in_d_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02734 vdd bsrmux_0_shr n27 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02733 vdd n79 n676 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02732 n676 n79 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02731 vdd n66 bsrmux_14_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02730 bsrmux_14_f1 n66 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02729 vdd n79 n676 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02728 vdd n78 n79 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02727 n78 in_d_28 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02726 vdd bsrmux_0_shr n78 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02725 vdd n66 bsrmux_14_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02724 vdd n65 n66 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02723 n65 in_d_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02722 vdd bsrmux_0_shr n65 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02721 vdd n114 n673 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02720 n673 n114 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02719 vdd n105 bsrmux_13_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02718 bsrmux_13_f1 n105 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02717 vdd n114 n673 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02716 vdd n112 n114 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02715 n112 in_d_26 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02714 vdd bsrmux_0_shr n112 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02713 vdd n105 bsrmux_13_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02712 vdd n104 n105 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02711 n104 in_d_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02710 vdd bsrmux_0_shr n104 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02709 vdd n153 n671 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02708 n671 n153 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02707 vdd n145 bsrmux_12_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02706 bsrmux_12_f1 n145 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02705 vdd n153 n671 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02704 vdd n151 n153 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02703 n151 in_d_24 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02702 vdd bsrmux_0_shr n151 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02701 vdd n145 bsrmux_12_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02700 vdd n144 n145 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02699 n144 in_d_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02698 vdd bsrmux_0_shr n144 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02697 vdd n191 n666 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02696 n666 n191 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02695 vdd n180 bsrmux_11_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02694 bsrmux_11_f1 n180 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02693 vdd n191 n666 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02692 vdd n189 n191 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02691 n189 in_d_22 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02690 vdd bsrmux_0_shr n189 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02689 vdd n180 bsrmux_11_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02688 vdd n179 n180 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02687 n179 in_d_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02686 vdd bsrmux_0_shr n179 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02685 vdd n229 n662 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02684 n662 n229 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02683 vdd n218 bsrmux_10_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02682 bsrmux_10_f1 n218 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02681 vdd n229 n662 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02680 vdd n227 n229 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02679 n227 in_d_20 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02678 vdd bsrmux_0_shr n227 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02677 vdd n218 bsrmux_10_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02676 vdd n217 n218 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02675 n217 in_d_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02674 vdd bsrmux_0_shr n217 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02673 vdd n267 n656 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02672 n656 n267 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02671 vdd n256 bsrmux_9_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02670 bsrmux_9_f1 n256 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02669 vdd n267 n656 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02668 vdd n266 n267 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02667 n266 in_d_18 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02666 vdd bsrmux_0_shr n266 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02665 vdd n256 bsrmux_9_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02664 vdd n255 n256 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02663 n255 in_d_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02662 vdd bsrmux_0_shr n255 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02661 vdd n304 n653 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02660 n653 n304 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02659 vdd n294 bsrmux_8_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02658 bsrmux_8_f1 n294 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02657 vdd n304 n653 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02656 vdd n302 n304 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02655 n302 in_d_16 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02654 vdd bsrmux_0_shr n302 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02653 vdd n294 bsrmux_8_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02652 vdd n293 n294 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02651 n293 in_d_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02650 vdd bsrmux_0_shr n293 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02649 vdd n343 n652 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02648 n652 n343 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02647 vdd n334 bsrmux_7_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02646 bsrmux_7_f1 n334 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02645 vdd n343 n652 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02644 vdd n341 n343 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02643 n341 in_d_14 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02642 vdd bsrmux_0_shr n341 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02641 vdd n334 bsrmux_7_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02640 vdd n333 n334 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02639 n333 in_d_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02638 vdd bsrmux_0_shr n333 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02637 vdd n381 n646 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02636 n646 n381 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02635 vdd n370 bsrmux_6_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02634 bsrmux_6_f1 n370 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02633 vdd n381 n646 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02632 vdd n379 n381 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02631 n379 in_d_12 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02630 vdd bsrmux_0_shr n379 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02629 vdd n370 bsrmux_6_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02628 vdd n369 n370 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02627 n369 in_d_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02626 vdd bsrmux_0_shr n369 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02625 vdd n419 n641 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02624 n641 n419 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02623 vdd n408 bsrmux_5_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02622 bsrmux_5_f1 n408 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02621 vdd n419 n641 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02620 vdd n417 n419 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02619 n417 in_d_10 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02618 vdd bsrmux_0_shr n417 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02617 vdd n408 bsrmux_5_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02616 vdd n407 n408 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02615 n407 in_d_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02614 vdd bsrmux_0_shr n407 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02613 vdd n457 n636 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02612 n636 n457 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02611 vdd n446 bsrmux_4_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02610 bsrmux_4_f1 n446 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02609 vdd n457 n636 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02608 vdd n455 n457 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02607 n455 in_d_8 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02606 vdd bsrmux_0_shr n455 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02605 vdd n446 bsrmux_4_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02604 vdd n445 n446 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02603 n445 in_d_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02602 vdd bsrmux_0_shr n445 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02601 vdd n501 n633 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02600 n633 n501 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02599 vdd n487 bsrmux_3_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02598 bsrmux_3_f1 n487 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02597 vdd n501 n633 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02596 vdd n500 n501 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02595 n500 in_d_6 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02594 vdd bsrmux_0_shr n500 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02593 vdd n487 bsrmux_3_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02592 vdd n486 n487 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02591 n486 in_d_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02590 vdd bsrmux_0_shr n486 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02589 vdd n537 n632 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02588 n632 n537 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02587 vdd n528 bsrmux_2_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02586 bsrmux_2_f1 n528 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02585 vdd n537 n632 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02584 vdd n535 n537 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02583 n535 in_d_4 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02582 vdd bsrmux_0_shr n535 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02581 vdd n528 bsrmux_2_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02580 vdd n527 n528 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02579 n527 in_d_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02578 vdd bsrmux_0_shr n527 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02577 vdd n577 n627 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02576 n627 n577 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02575 vdd n566 bsrmux_1_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02574 bsrmux_1_f1 n566 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02573 vdd n577 n627 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02572 vdd n575 n577 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02571 n575 in_d_2 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02570 vdd bsrmux_0_shr n575 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02569 vdd n566 bsrmux_1_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02568 vdd n565 n566 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02567 n565 in_d_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02566 vdd bsrmux_0_shr n565 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02565 vdd n619 n622 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02564 n622 n619 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02563 vdd n606 bsrmux_0_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02562 bsrmux_0_f1 n606 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02561 vdd n619 n622 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02560 vdd n617 n619 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02559 n617 in_d_0 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02558 vdd bsrmux_0_shr n617 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02557 vdd n606 bsrmux_0_f1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02556 vdd n605 n606 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_02555 n605 in_d_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02554 vdd bsrmux_0_shr n605 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02553 bsm_0_15_in_2 n41 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02552 vdd n41 bsm_0_15_in_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02551 bsm_0_15_in_2 n41 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02550 vdd n43 n41 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02549 n41 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02548 vdd bshlmx_0_lsl n43 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02547 n43 in_d_30 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02546 bslmux_15_out_1 n30 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02545 vdd n30 bslmux_15_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02544 bslmux_15_out_1 n30 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02543 vdd n31 n30 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02542 n30 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02541 vdd bshlmx_0_lsl n31 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02540 n31 in_d_31 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02539 bslmux_14_out_2 n80 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02538 vdd n80 bslmux_14_out_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02537 bslmux_14_out_2 n80 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02536 vdd n84 n80 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02535 n80 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02534 vdd bshlmx_0_lsl n84 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02533 n84 in_d_28 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02532 bslmux_14_out_1 n69 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02531 vdd n69 bslmux_14_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02530 bslmux_14_out_1 n69 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02529 vdd n68 n69 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02528 n69 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02527 vdd bshlmx_0_lsl n68 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02526 n68 in_d_29 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02525 bslmux_13_out_2 n116 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02524 vdd n116 bslmux_13_out_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02523 bslmux_13_out_2 n116 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02522 vdd n118 n116 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02521 n116 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02520 vdd bshlmx_0_lsl n118 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02519 n118 in_d_26 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02518 bslmux_13_out_1 n106 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02517 vdd n106 bslmux_13_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02516 bslmux_13_out_1 n106 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02515 vdd n97 n106 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02514 n106 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02513 vdd bshlmx_0_lsl n97 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02512 n97 in_d_27 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02511 bslmux_12_out_2 n156 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02510 vdd n156 bslmux_12_out_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02509 bslmux_12_out_2 n156 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02508 vdd n158 n156 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02507 n156 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02506 vdd bshlmx_0_lsl n158 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02505 n158 in_d_24 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02504 bslmux_12_out_1 n146 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02503 vdd n146 bslmux_12_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02502 bslmux_12_out_1 n146 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02501 vdd n140 n146 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02500 n146 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02499 vdd bshlmx_0_lsl n140 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02498 n140 in_d_25 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02497 bslmux_11_out_2 n194 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02496 vdd n194 bslmux_11_out_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02495 bslmux_11_out_2 n194 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02494 vdd n196 n194 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02493 n194 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02492 vdd bshlmx_0_lsl n196 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02491 n196 in_d_22 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02490 bslmux_11_out_1 n182 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02489 vdd n182 bslmux_11_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02488 bslmux_11_out_1 n182 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02487 vdd n183 n182 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02486 n182 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02485 vdd bshlmx_0_lsl n183 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02484 n183 in_d_23 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02483 bsm_0_10_in_2 n232 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02482 vdd n232 bsm_0_10_in_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02481 bsm_0_10_in_2 n232 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02480 vdd n234 n232 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02479 n232 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02478 vdd bshlmx_0_lsl n234 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02477 n234 in_d_20 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02476 bslmux_10_out_1 n220 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02475 vdd n220 bslmux_10_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02474 bslmux_10_out_1 n220 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02473 vdd n221 n220 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02472 n220 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02471 vdd bshlmx_0_lsl n221 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02470 n221 in_d_21 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02469 bsm_0_9_in_2 n270 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02468 vdd n270 bsm_0_9_in_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02467 bsm_0_9_in_2 n270 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02466 vdd n273 n270 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02465 n270 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02464 vdd bshlmx_0_lsl n273 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02463 n273 in_d_18 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02462 bslmux_9_out_1 n259 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02461 vdd n259 bslmux_9_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02460 bslmux_9_out_1 n259 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02459 vdd n258 n259 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02458 n259 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02457 vdd bshlmx_0_lsl n258 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02456 n258 in_d_19 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02455 bslmux_8_out_2 n306 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02454 vdd n306 bslmux_8_out_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02453 bslmux_8_out_2 n306 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02452 vdd n309 n306 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02451 n306 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02450 vdd bshlmx_0_lsl n309 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02449 n309 in_d_16 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02448 bslmux_8_out_1 n295 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02447 vdd n295 bslmux_8_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02446 bslmux_8_out_1 n295 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02445 vdd n297 n295 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02444 n295 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02443 vdd bshlmx_0_lsl n297 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02442 n297 in_d_17 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02441 bslmux_7_out_2 n346 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02440 vdd n346 bslmux_7_out_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02439 bslmux_7_out_2 n346 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02438 vdd n348 n346 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02437 n346 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02436 vdd bshlmx_0_lsl n348 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02435 n348 in_d_14 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02434 bslmux_7_out_1 n335 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02433 vdd n335 bslmux_7_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02432 bslmux_7_out_1 n335 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02431 vdd n325 n335 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02430 n335 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02429 vdd bshlmx_0_lsl n325 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02428 n325 in_d_15 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02427 bslmux_6_out_2 n384 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02426 vdd n384 bslmux_6_out_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02425 bslmux_6_out_2 n384 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02424 vdd n386 n384 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02423 n384 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02422 vdd bshlmx_0_lsl n386 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02421 n386 in_d_12 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02420 bslmux_6_out_1 n372 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02419 vdd n372 bslmux_6_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02418 bslmux_6_out_1 n372 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02417 vdd n373 n372 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02416 n372 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02415 vdd bshlmx_0_lsl n373 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02414 n373 in_d_13 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02413 bslmux_5_out_2 n422 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02412 vdd n422 bslmux_5_out_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02411 bslmux_5_out_2 n422 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02410 vdd n424 n422 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02409 n422 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02408 vdd bshlmx_0_lsl n424 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02407 n424 in_d_10 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02406 bslmux_5_out_1 n410 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02405 vdd n410 bslmux_5_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02404 bslmux_5_out_1 n410 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02403 vdd n411 n410 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02402 n410 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02401 vdd bshlmx_0_lsl n411 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02400 n411 in_d_11 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02399 bslmux_4_out_2 n460 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02398 vdd n460 bslmux_4_out_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02397 bslmux_4_out_2 n460 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02396 vdd n462 n460 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02395 n460 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02394 vdd bshlmx_0_lsl n462 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02393 n462 in_d_8 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02392 bslmux_4_out_1 n448 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02391 vdd n448 bslmux_4_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02390 bslmux_4_out_1 n448 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02389 vdd n450 n448 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02388 n448 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02387 vdd bshlmx_0_lsl n450 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02386 n450 in_d_9 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02385 bslmux_3_out_2 n496 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02384 vdd n496 bslmux_3_out_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02383 bslmux_3_out_2 n496 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02382 vdd n502 n496 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02381 n496 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02380 vdd bshlmx_0_lsl n502 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02379 n502 in_d_6 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02378 bslmux_3_out_1 n490 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02377 vdd n490 bslmux_3_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02376 bslmux_3_out_1 n490 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02375 vdd n489 n490 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02374 n490 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02373 vdd bshlmx_0_lsl n489 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02372 n489 in_d_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02371 bslmux_2_out_2 n540 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02370 vdd n540 bslmux_2_out_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02369 bslmux_2_out_2 n540 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02368 vdd n542 n540 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02367 n540 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02366 vdd bshlmx_0_lsl n542 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02365 n542 in_d_4 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02364 bslmux_2_out_1 n529 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02363 vdd n529 bslmux_2_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02362 bslmux_2_out_1 n529 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02361 vdd n519 n529 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02360 n529 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02359 vdd bshlmx_0_lsl n519 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02358 n519 in_d_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02357 bslmux_1_out_2 n580 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02356 vdd n580 bslmux_1_out_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02355 bslmux_1_out_2 n580 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02354 vdd n582 n580 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02353 n580 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02352 vdd bshlmx_0_lsl n582 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02351 n582 in_d_2 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02350 bslmux_1_out_1 n568 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02349 vdd n568 bslmux_1_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02348 bslmux_1_out_1 n568 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02347 vdd n569 n568 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02346 n568 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02345 vdd bshlmx_0_lsl n569 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02344 n569 in_d_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02343 bslmux_0_out_2 n688 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02342 vdd n688 bslmux_0_out_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02341 bslmux_0_out_2 n688 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02340 vdd n691 n688 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02339 n688 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02338 vdd bshlmx_0_lsl n691 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02337 n691 in_d_0 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02336 bslmux_0_out_1 n608 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02335 vdd n608 bslmux_0_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02334 bslmux_0_out_1 n608 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02333 vdd n610 n608 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_02332 n608 bshlmx_0_asr vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_02331 vdd bshlmx_0_lsl n610 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02330 n610 in_d_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_02329 vdd bsdand_15_out_2 n48 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02328 bssnbl_15_out_1 bssnbl_15_in_2 vdd vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_02327 vdd bssnbl_15_in_2 bssnbl_15_out_1 vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_02326 bssnbl_15_out_1 bssnbl_15_in_2 vdd vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_02325 bslmux_15_com_2 n48 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02324 vdd n48 bslmux_15_com_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02323 bslmux_15_com_2 n48 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02322 vdd bsssel_14_out_2_s n86 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02321 vdd bssnbl_14_in_1 n71 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02320 bssnbl_14_out_1 n71 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02319 vdd n71 bssnbl_14_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02318 bssnbl_14_out_1 n71 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02317 bslmux_14_com_2 n86 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02316 vdd n86 bslmux_14_com_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02315 bslmux_14_com_2 n86 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02314 vdd bssnbl_13_in_2 n126 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02313 vdd bssnbl_13_in_1 n109 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02312 bssnbl_13_out_1 n109 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02311 vdd n109 bssnbl_13_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02310 bssnbl_13_out_1 n109 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02309 bslmux_13_com_2 n126 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02308 vdd n126 bslmux_13_com_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02307 bslmux_13_com_2 n126 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02306 vdd bssnbl_12_in_2 n161 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02305 vdd bssnbl_12_in_1 n148 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02304 bssnbl_12_out_1 n148 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02303 vdd n148 bssnbl_12_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02302 bssnbl_12_out_1 n148 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02301 bslmux_12_com_2 n161 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02300 vdd n161 bslmux_12_com_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02299 bslmux_12_com_2 n161 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02298 vdd bsssel_11_out_2_s n200 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02297 vdd bsssel_11_out_1_s n184 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02296 bssnbl_11_out_1 n184 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02295 vdd n184 bssnbl_11_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02294 bssnbl_11_out_1 n184 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02293 bslmux_11_com_2 n200 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02292 vdd n200 bslmux_11_com_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02291 bslmux_11_com_2 n200 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02290 vdd bsssel_10_out_2_s n238 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02289 vdd bsssel_10_out_1_s n222 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02288 bssnbl_10_out_1 n222 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02287 vdd n222 bssnbl_10_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02286 bssnbl_10_out_1 n222 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02285 bslmux_10_com_2 n238 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02284 vdd n238 bslmux_10_com_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02283 bslmux_10_com_2 n238 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02282 vdd bsssel_9_out_2_s n276 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02281 vdd bssnbl_9_in_1 n261 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02280 bssnbl_9_out_1 n261 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02279 vdd n261 bssnbl_9_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02278 bssnbl_9_out_1 n261 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02277 bslmux_9_com_2 n276 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02276 vdd n276 bslmux_9_com_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02275 bslmux_9_com_2 n276 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02274 vdd bssnbl_8_in_2 n316 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02273 vdd bssnbl_8_in_1 n299 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02272 bssnbl_8_out_1 n299 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02271 vdd n299 bssnbl_8_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02270 bssnbl_8_out_1 n299 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02269 bslmux_8_com_2 n316 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02268 vdd n316 bslmux_8_com_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02267 bslmux_8_com_2 n316 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02266 vdd bssnbl_7_in_2 n351 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02265 vdd bssnbl_7_in_1 n338 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02264 bssnbl_7_out_1 n338 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02263 vdd n338 bssnbl_7_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02262 bssnbl_7_out_1 n338 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02261 bslmux_7_com_2 n351 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02260 vdd n351 bslmux_7_com_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02259 bslmux_7_com_2 n351 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02258 vdd bsssel_6_out_2_s n390 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02257 vdd bsssel_6_out_1_s n374 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02256 bssnbl_6_out_1 n374 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02255 vdd n374 bssnbl_6_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02254 bssnbl_6_out_1 n374 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02253 bslmux_6_com_2 n390 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02252 vdd n390 bslmux_6_com_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02251 bslmux_6_com_2 n390 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02250 vdd bsssel_5_out_2_s n428 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02249 vdd bsssel_5_out_1_s n412 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02248 bssnbl_5_out_1 n412 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02247 vdd n412 bssnbl_5_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02246 bssnbl_5_out_1 n412 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02245 bslmux_5_com_2 n428 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02244 vdd n428 bslmux_5_com_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02243 bslmux_5_com_2 n428 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02242 vdd bsssel_4_out_2_s n464 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02241 vdd bssnbl_4_in_1 n452 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02240 bssnbl_4_out_1 n452 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02239 vdd n452 bssnbl_4_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02238 bssnbl_4_out_1 n452 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02237 bslmux_4_com_2 n464 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02236 vdd n464 bslmux_4_com_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02235 bslmux_4_com_2 n464 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02234 vdd bsssel_3_out_2_s n508 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02233 vdd bssnbl_3_in_1 n492 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02232 bssnbl_3_out_1 n492 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02231 vdd n492 bssnbl_3_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02230 bssnbl_3_out_1 n492 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02229 bslmux_3_com_2 n508 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02228 vdd n508 bslmux_3_com_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02227 bslmux_3_com_2 n508 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02226 vdd bssnbl_2_in_2 n558 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02225 vdd bssnbl_2_in_1 n532 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02224 bssnbl_2_out_1 n532 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02223 vdd n532 bssnbl_2_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02222 bssnbl_2_out_1 n532 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02221 bslmux_2_com_2 n558 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02220 vdd n558 bslmux_2_com_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02219 bslmux_2_com_2 n558 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02218 vdd bsssel_1_out_2_s n586 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02217 vdd bsssel_1_out_1_s n570 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02216 bssnbl_1_out_1 n570 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02215 vdd n570 bssnbl_1_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02214 bssnbl_1_out_1 n570 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02213 bslmux_1_com_2 n586 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02212 vdd n586 bslmux_1_com_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02211 bslmux_1_com_2 n586 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02210 vdd bsssel_0_out_2_s n696 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02209 vdd bsssel_0_out_1_s n611 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02208 bssnbl_0_out_1 n611 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02207 vdd n611 bssnbl_0_out_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02206 bssnbl_0_out_1 n611 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02205 bssnbl_0_out_2 n696 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02204 vdd n696 bssnbl_0_out_2 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02203 bssnbl_0_out_2 n696 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02202 vdd bsdand_15_out_1 bssnbl_15_in_2 vdd TP L=0.18U W=3.06U AS=1.1016P 
+ AD=1.1016P PS=6.84U PD=6.84U 
Mtr_02201 bssnbl_15_in_2 n699 vdd vdd TP L=0.18U W=3.06U AS=1.1016P AD=1.1016P 
+ PS=6.84U PD=6.84U 
Mtr_02200 vdd n693 bssnbl_15_zero vdd TP L=0.18U W=3.06U AS=1.1016P AD=1.1016P 
+ PS=6.84U PD=6.84U 
Mtr_02199 bssnbl_15_zero bsdand_15_out_1 vdd vdd TP L=0.18U W=3.06U AS=1.1016P 
+ AD=1.1016P PS=6.84U PD=6.84U 
Mtr_02198 vdd n71 bssnbl_14_in_1 vdd TP L=0.36U W=0.54U AS=0.1944P AD=0.1944P 
+ PS=1.8U PD=1.8U 
Mtr_02197 bsssel_14_out_2_s n86 vdd vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02196 vdd n109 bssnbl_13_in_1 vdd TP L=0.36U W=0.54U AS=0.1944P AD=0.1944P 
+ PS=1.8U PD=1.8U 
Mtr_02195 bssnbl_13_in_2 n126 vdd vdd TP L=0.36U W=0.54U AS=0.1944P AD=0.1944P 
+ PS=1.8U PD=1.8U 
Mtr_02194 vdd n148 bssnbl_12_in_1 vdd TP L=0.36U W=0.54U AS=0.1944P AD=0.1944P 
+ PS=1.8U PD=1.8U 
Mtr_02193 bssnbl_12_in_2 n161 vdd vdd TP L=0.36U W=0.54U AS=0.1944P AD=0.1944P 
+ PS=1.8U PD=1.8U 
Mtr_02192 vdd n184 bsssel_11_out_1_s vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02191 bsssel_11_out_2_s n200 vdd vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02190 vdd n222 bsssel_10_out_1_s vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02189 bsssel_10_out_2_s n238 vdd vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02188 vdd n261 bssnbl_9_in_1 vdd TP L=0.36U W=0.54U AS=0.1944P AD=0.1944P 
+ PS=1.8U PD=1.8U 
Mtr_02187 bsssel_9_out_2_s n276 vdd vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02186 vdd n299 bssnbl_8_in_1 vdd TP L=0.36U W=0.54U AS=0.1944P AD=0.1944P 
+ PS=1.8U PD=1.8U 
Mtr_02185 bssnbl_8_in_2 n316 vdd vdd TP L=0.36U W=0.54U AS=0.1944P AD=0.1944P 
+ PS=1.8U PD=1.8U 
Mtr_02184 vdd n338 bssnbl_7_in_1 vdd TP L=0.36U W=0.54U AS=0.1944P AD=0.1944P 
+ PS=1.8U PD=1.8U 
Mtr_02183 bssnbl_7_in_2 n351 vdd vdd TP L=0.36U W=0.54U AS=0.1944P AD=0.1944P 
+ PS=1.8U PD=1.8U 
Mtr_02182 vdd n374 bsssel_6_out_1_s vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02181 bsssel_6_out_2_s n390 vdd vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02180 vdd n412 bsssel_5_out_1_s vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02179 bsssel_5_out_2_s n428 vdd vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02178 vdd n452 bssnbl_4_in_1 vdd TP L=0.36U W=0.54U AS=0.1944P AD=0.1944P 
+ PS=1.8U PD=1.8U 
Mtr_02177 bsssel_4_out_2_s n464 vdd vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02176 vdd n492 bssnbl_3_in_1 vdd TP L=0.36U W=0.54U AS=0.1944P AD=0.1944P 
+ PS=1.8U PD=1.8U 
Mtr_02175 bsssel_3_out_2_s n508 vdd vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02174 vdd n532 bssnbl_2_in_1 vdd TP L=0.36U W=0.54U AS=0.1944P AD=0.1944P 
+ PS=1.8U PD=1.8U 
Mtr_02173 bssnbl_2_in_2 n558 vdd vdd TP L=0.36U W=0.54U AS=0.1944P AD=0.1944P 
+ PS=1.8U PD=1.8U 
Mtr_02172 vdd n570 bsssel_1_out_1_s vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02171 bsssel_1_out_2_s n586 vdd vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02170 vdd n611 bsssel_0_out_1_s vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02169 bsssel_0_out_2_s n696 vdd vdd TP L=0.36U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_02168 bsdand_15_out_1 n33 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02167 n33 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02166 vdd bsdand_0_v_4_2 n33 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02165 n33 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02164 vdd bsdand_1_v_0_1 n33 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02163 n33 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02162 n50 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02161 vdd bsdand_0_v_4_1 n50 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02160 n50 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02159 vdd bsdand_1_v_0_1 n50 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02158 n50 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02157 bsdand_15_out_2 n50 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02156 bsdand_14_out_1 n72 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02155 n72 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02154 vdd bsdand_0_v_4_1 n72 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02153 n72 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02152 vdd bsdand_0_v_0_1 n72 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02151 n72 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02150 n89 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02149 vdd bsdand_0_v_4_2 n89 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02148 n89 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02147 vdd bsdand_0_v_0_1 n89 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02146 n89 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02145 bsdand_14_out_2 n89 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02144 bsdand_13_out_1 n110 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02143 n110 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02142 vdd bsdand_0_v_4_1 n110 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02141 n110 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02140 vdd bsdand_1_v_0_1 n110 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02139 n110 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02138 n131 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02137 vdd bsdand_0_v_4_2 n131 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02136 n131 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02135 vdd bsdand_1_v_0_1 n131 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02134 n131 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02133 bsdand_13_out_2 n131 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02132 bsdand_12_out_1 n149 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02131 n149 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02130 vdd bsdand_0_v_4_1 n149 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02129 n149 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02128 vdd bsdand_0_v_0_1 n149 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02127 n149 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02126 n165 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02125 vdd bsdand_0_v_4_2 n165 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02124 n165 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02123 vdd bsdand_0_v_0_1 n165 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02122 n165 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02121 bsdand_12_out_2 n165 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02120 bsdand_11_out_1 n186 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02119 n186 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02118 vdd bsdand_0_v_4_1 n186 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02117 n186 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02116 vdd bsdand_1_v_0_1 n186 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02115 n186 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02114 n204 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02113 vdd bsdand_0_v_4_2 n204 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02112 n204 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02111 vdd bsdand_1_v_0_1 n204 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02110 n204 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02109 bsdand_11_out_2 n204 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02108 bsdand_10_out_1 n224 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02107 n224 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02106 vdd bsdand_0_v_4_1 n224 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02105 n224 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02104 vdd bsdand_0_v_0_1 n224 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02103 n224 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02102 n240 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02101 vdd bsdand_0_v_4_2 n240 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02100 n240 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02099 vdd bsdand_0_v_0_1 n240 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02098 n240 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02097 bsdand_10_out_2 n240 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02096 bsdand_9_out_1 n262 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02095 n262 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02094 vdd bsdand_0_v_4_1 n262 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02093 n262 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02092 vdd bsdand_1_v_0_1 n262 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02091 n262 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02090 n279 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02089 vdd bsdand_0_v_4_2 n279 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02088 n279 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02087 vdd bsdand_1_v_0_1 n279 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02086 n279 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02085 bsdand_9_out_2 n279 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02084 bsdand_8_out_1 n300 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02083 n300 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02082 vdd bsdand_0_v_4_1 n300 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02081 n300 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02080 vdd bsdand_0_v_0_1 n300 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02079 n300 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02078 n317 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02077 vdd bsdand_0_v_4_2 n317 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02076 n317 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02075 vdd bsdand_0_v_0_1 n317 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02074 n317 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02073 bsdand_8_out_2 n317 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02072 bsdand_7_out_1 n339 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02071 n339 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02070 vdd bsdand_0_v_4_1 n339 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02069 n339 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02068 vdd bsdand_1_v_0_1 n339 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02067 n339 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02066 n355 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02065 vdd bsdand_0_v_4_2 n355 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02064 n355 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02063 vdd bsdand_1_v_0_1 n355 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02062 n355 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02061 bsdand_7_out_2 n355 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02060 bsdand_6_out_1 n376 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02059 n376 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02058 vdd bsdand_0_v_4_1 n376 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02057 n376 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02056 vdd bsdand_0_v_0_1 n376 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02055 n376 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02054 n394 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02053 vdd bsdand_0_v_4_2 n394 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02052 n394 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02051 vdd bsdand_0_v_0_1 n394 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02050 n394 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02049 bsdand_6_out_2 n394 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02048 bsdand_5_out_1 n414 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02047 n414 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02046 vdd bsdand_0_v_4_1 n414 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02045 n414 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02044 vdd bsdand_1_v_0_1 n414 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02043 n414 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02042 n430 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02041 vdd bsdand_0_v_4_2 n430 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02040 n430 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02039 vdd bsdand_1_v_0_1 n430 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02038 n430 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02037 bsdand_5_out_2 n430 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02036 bsdand_4_out_1 n453 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02035 n453 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02034 vdd bsdand_0_v_4_1 n453 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02033 n453 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02032 vdd bsdand_0_v_0_1 n453 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02031 n453 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02030 n468 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02029 vdd bsdand_0_v_4_2 n468 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02028 n468 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02027 vdd bsdand_0_v_0_1 n468 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02026 n468 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02025 bsdand_4_out_2 n468 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02024 bsdand_3_out_1 n493 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02023 n493 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02022 vdd bsdand_0_v_4_1 n493 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02021 n493 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02020 vdd bsdand_1_v_0_1 n493 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02019 n493 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02018 n509 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02017 vdd bsdand_0_v_4_2 n509 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02016 n509 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02015 vdd bsdand_1_v_0_1 n509 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02014 n509 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02013 bsdand_3_out_2 n509 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02012 bsdand_2_out_1 n533 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02011 n533 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02010 vdd bsdand_0_v_4_1 n533 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02009 n533 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02008 vdd bsdand_0_v_0_1 n533 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02007 n533 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02006 n548 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02005 vdd bsdand_0_v_4_2 n548 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02004 n548 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02003 vdd bsdand_0_v_0_1 n548 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02002 n548 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_02001 bsdand_2_out_2 n548 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_02000 bsdand_1_out_1 n572 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01999 n572 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01998 vdd bsdand_0_v_4_1 n572 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01997 n572 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01996 vdd bsdand_1_v_0_1 n572 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01995 n572 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01994 n590 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01993 vdd bsdand_0_v_4_2 n590 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01992 n590 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01991 vdd bsdand_1_v_0_1 n590 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01990 n590 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01989 bsdand_1_out_2 n590 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01988 bsdand_0_out_1 n613 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01987 n613 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01986 vdd bsdand_0_v_4_1 n613 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01985 n613 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01984 vdd bsdand_0_v_0_1 n613 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01983 n613 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01982 n705 bsdand_0_v_3_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01981 vdd bsdand_0_v_4_2 n705 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01980 n705 bsdand_0_na1 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01979 vdd bsdand_0_v_0_1 n705 vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01978 n705 bsdand_0_v_2_2 vdd vdd TP L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_01977 bsdand_0_out_2 n705 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01976 bsdand_0_v_4_2 bsdand_0_v_4_1 vdd vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01975 vdd bsdand_0_v_4_1 bsdand_0_v_4_2 vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01974 bsdand_0_v_4_2 bsdand_0_v_4_1 vdd vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01973 bsdand_0_v_4_1 n475 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01972 vdd n475 bsdand_0_v_4_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01971 bsdand_0_v_4_1 n475 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01970 vdd in_s_4 n475 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_01969 bsdand_0_v_3_2 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01968 vdd bsdand_0_v_3_1 bsdand_0_v_3_2 vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01967 bsdand_0_v_3_2 bsdand_0_v_3_1 vdd vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01966 bsdand_0_v_3_1 n516 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01965 vdd n516 bsdand_0_v_3_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01964 bsdand_0_v_3_1 n516 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01963 vdd in_s_3 n516 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_01962 bsdand_0_v_2_2 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01961 vdd bsdand_0_v_2_1 bsdand_0_v_2_2 vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01960 bsdand_0_v_2_2 bsdand_0_v_2_1 vdd vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01959 bsdand_0_v_2_1 n553 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01958 vdd n553 bsdand_0_v_2_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01957 bsdand_0_v_2_1 n553 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01956 vdd in_s_2 n553 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_01955 bsdand_0_na1 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01954 vdd bsdand_0_v_1_1 bsdand_0_na1 vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01953 bsdand_0_na1 bsdand_0_v_1_1 vdd vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01952 bsdand_0_v_1_1 n595 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01951 vdd n595 bsdand_0_v_1_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01950 bsdand_0_v_1_1 n595 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01949 vdd in_s_1 n595 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_01948 bsdand_1_v_0_1 bsdand_0_v_0_1 vdd vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01947 vdd bsdand_0_v_0_1 bsdand_1_v_0_1 vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01946 bsdand_1_v_0_1 bsdand_0_v_0_1 vdd vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01945 bsdand_0_v_0_1 n715 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01944 vdd n715 bsdand_0_v_0_1 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01943 bsdand_0_v_0_1 n715 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01942 vdd in_s_0 n715 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_01941 bsrmux_0_shr bshmat_0_nshr vss vss TN L=0.18U W=4.86U AS=1.7496P 
+ AD=1.7496P PS=10.44U PD=10.44U 
Mtr_01940 n5 rot vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01939 vss n5 n1 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01938 n1 bshsel_0_nright n3 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01937 n12 n3 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01936 vss n11 bshcmd_0_nasr vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01935 n7 n12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01934 n8 in_d_31 n7 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01933 n11 ext n8 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01932 n10 bshlmx_0_nnleft n9 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01931 vss n5 n10 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01930 bshmat_0_nshr n9 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01929 vss n12 bshlmx_0_lsl vss TN L=0.18U W=4.86U AS=1.7496P AD=1.7496P 
+ PS=10.44U PD=10.44U 
Mtr_01928 bshlmx_0_asr bshcmd_0_nasr vss vss TN L=0.18U W=4.86U AS=1.7496P 
+ AD=1.7496P PS=10.44U PD=10.44U 
Mtr_01927 bshmatr_0_comr0 bssnbl_15_zero vss vss TN L=0.18U W=4.86U AS=1.7496P 
+ AD=1.7496P PS=10.44U PD=10.44U 
Mtr_01926 n693 bshlmx_0_nnleft vss vss TN L=0.18U W=4.86U AS=1.7496P 
+ AD=1.7496P PS=10.44U PD=10.44U 
Mtr_01925 vss bshsel_0_nright n699 vss TN L=0.18U W=4.86U AS=1.7496P 
+ AD=1.7496P PS=10.44U PD=10.44U 
Mtr_01924 vss bshsel_0_nright bshlmx_0_nnleft vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01923 bshsel_0_nright left vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01922 vss bsm_0_15_out_2_s out_d_30 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01921 vss bsoout_15_out_1_s out_d_31 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01920 vss bsoout_14_out_2_s out_d_28 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01919 vss bsoout_14_out_1_s out_d_29 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01918 vss bsoout_13_out_2_s out_d_26 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01917 vss bsoout_13_out_1_s out_d_27 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01916 vss bsm_0_12_out_2_s out_d_24 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01915 vss bsoout_12_out_1_s out_d_25 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01914 vss bsm_0_11_out_2_s out_d_22 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01913 vss bsoout_11_out_1_s out_d_23 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01912 vss bsm_0_10_out_2_s out_d_20 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01911 vss bsoout_10_out_1_s out_d_21 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01910 vss bsm_0_9_out_2_s out_d_18 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01909 vss bsoout_9_out_1_s out_d_19 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01908 vss bsoout_8_out_2_s out_d_16 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01907 vss bsoout_8_out_1_s out_d_17 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01906 vss bsm_0_7_out_2_s out_d_14 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01905 vss bsoout_7_out_1_s out_d_15 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01904 vss bsm_0_6_out_2_s out_d_12 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01903 vss bsoout_6_out_1_s out_d_13 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01902 vss bsm_0_5_out_2_s out_d_10 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01901 vss bsoout_5_out_1_s out_d_11 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01900 vss bsm_0_4_out_2_s out_d_8 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01899 vss bsoout_4_out_1_s out_d_9 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01898 vss bsoout_3_out_2_s out_d_6 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01897 vss bsoout_3_out_1_s out_d_7 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01896 vss bsm_0_2_out_2_s out_d_4 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01895 vss bsoout_2_out_1_s out_d_5 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01894 vss bsm_0_1_out_2_s out_d_2 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01893 vss bsoout_1_out_1_s out_d_3 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01892 vss bsm_0_0_out_2_s out_d_0 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01891 vss bsoout_0_out_1_s out_d_1 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_01890 vss n38 n681 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01889 n681 n38 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01888 vss n28 bsrmux_15_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01887 bsrmux_15_f1 n28 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01886 vss n38 n681 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01885 vss n36 n38 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01884 n37 in_d_30 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01883 n36 bsrmux_0_shr n37 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01882 vss n28 bsrmux_15_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01881 vss n27 n28 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01880 n27 bsrmux_0_shr n17 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01879 n17 in_d_31 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01878 vss n79 n676 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01877 n676 n79 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01876 vss n66 bsrmux_14_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01875 bsrmux_14_f1 n66 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01874 vss n79 n676 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01873 vss n78 n79 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01872 n74 in_d_28 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01871 n78 bsrmux_0_shr n74 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01870 vss n66 bsrmux_14_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01869 vss n65 n66 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01868 n65 bsrmux_0_shr n56 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01867 n56 in_d_29 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01866 vss n114 n673 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01865 n673 n114 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01864 vss n105 bsrmux_13_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01863 bsrmux_13_f1 n105 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01862 vss n114 n673 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01861 vss n112 n114 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01860 n113 in_d_26 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01859 n112 bsrmux_0_shr n113 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01858 vss n105 bsrmux_13_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01857 vss n104 n105 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01856 n104 bsrmux_0_shr n95 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01855 n95 in_d_27 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01854 vss n153 n671 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01853 n671 n153 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01852 vss n145 bsrmux_12_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01851 bsrmux_12_f1 n145 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01850 vss n153 n671 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01849 vss n151 n153 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01848 n152 in_d_24 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01847 n151 bsrmux_0_shr n152 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01846 vss n145 bsrmux_12_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01845 vss n144 n145 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01844 n144 bsrmux_0_shr n137 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01843 n137 in_d_25 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01842 vss n191 n666 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01841 n666 n191 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01840 vss n180 bsrmux_11_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01839 bsrmux_11_f1 n180 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01838 vss n191 n666 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01837 vss n189 n191 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01836 n190 in_d_22 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01835 n189 bsrmux_0_shr n190 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01834 vss n180 bsrmux_11_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01833 vss n179 n180 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01832 n179 bsrmux_0_shr n169 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01831 n169 in_d_23 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01830 vss n229 n662 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01829 n662 n229 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01828 vss n218 bsrmux_10_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01827 bsrmux_10_f1 n218 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01826 vss n229 n662 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01825 vss n227 n229 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01824 n228 in_d_20 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01823 n227 bsrmux_0_shr n228 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01822 vss n218 bsrmux_10_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01821 vss n217 n218 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01820 n217 bsrmux_0_shr n208 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01819 n208 in_d_21 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01818 vss n267 n656 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01817 n656 n267 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01816 vss n256 bsrmux_9_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01815 bsrmux_9_f1 n256 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01814 vss n267 n656 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01813 vss n266 n267 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01812 n264 in_d_18 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01811 n266 bsrmux_0_shr n264 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01810 vss n256 bsrmux_9_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01809 vss n255 n256 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01808 n255 bsrmux_0_shr n246 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01807 n246 in_d_19 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01806 vss n304 n653 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01805 n653 n304 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01804 vss n294 bsrmux_8_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01803 bsrmux_8_f1 n294 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01802 vss n304 n653 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01801 vss n302 n304 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01800 n303 in_d_16 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01799 n302 bsrmux_0_shr n303 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01798 vss n294 bsrmux_8_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01797 vss n293 n294 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01796 n293 bsrmux_0_shr n285 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01795 n285 in_d_17 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01794 vss n343 n652 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01793 n652 n343 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01792 vss n334 bsrmux_7_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01791 bsrmux_7_f1 n334 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01790 vss n343 n652 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01789 vss n341 n343 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01788 n342 in_d_14 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01787 n341 bsrmux_0_shr n342 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01786 vss n334 bsrmux_7_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01785 vss n333 n334 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01784 n333 bsrmux_0_shr n323 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01783 n323 in_d_15 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01782 vss n381 n646 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01781 n646 n381 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01780 vss n370 bsrmux_6_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01779 bsrmux_6_f1 n370 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01778 vss n381 n646 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01777 vss n379 n381 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01776 n380 in_d_12 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01775 n379 bsrmux_0_shr n380 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01774 vss n370 bsrmux_6_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01773 vss n369 n370 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01772 n369 bsrmux_0_shr n359 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01771 n359 in_d_13 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01770 vss n419 n641 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01769 n641 n419 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01768 vss n408 bsrmux_5_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01767 bsrmux_5_f1 n408 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01766 vss n419 n641 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01765 vss n417 n419 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01764 n418 in_d_10 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01763 n417 bsrmux_0_shr n418 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01762 vss n408 bsrmux_5_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01761 vss n407 n408 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01760 n407 bsrmux_0_shr n398 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01759 n398 in_d_11 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01758 vss n457 n636 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01757 n636 n457 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01756 vss n446 bsrmux_4_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01755 bsrmux_4_f1 n446 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01754 vss n457 n636 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01753 vss n455 n457 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01752 n456 in_d_8 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01751 n455 bsrmux_0_shr n456 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01750 vss n446 bsrmux_4_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01749 vss n445 n446 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01748 n445 bsrmux_0_shr n436 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01747 n436 in_d_9 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01746 vss n501 n633 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01745 n633 n501 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01744 vss n487 bsrmux_3_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01743 bsrmux_3_f1 n487 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01742 vss n501 n633 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01741 vss n500 n501 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01740 n494 in_d_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01739 n500 bsrmux_0_shr n494 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01738 vss n487 bsrmux_3_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01737 vss n486 n487 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01736 n486 bsrmux_0_shr n476 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01735 n476 in_d_7 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01734 vss n537 n632 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01733 n632 n537 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01732 vss n528 bsrmux_2_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01731 bsrmux_2_f1 n528 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01730 vss n537 n632 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01729 vss n535 n537 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01728 n536 in_d_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01727 n535 bsrmux_0_shr n536 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01726 vss n528 bsrmux_2_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01725 vss n527 n528 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01724 n527 bsrmux_0_shr n517 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01723 n517 in_d_5 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01722 vss n577 n627 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01721 n627 n577 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01720 vss n566 bsrmux_1_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01719 bsrmux_1_f1 n566 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01718 vss n577 n627 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01717 vss n575 n577 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01716 n576 in_d_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01715 n575 bsrmux_0_shr n576 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01714 vss n566 bsrmux_1_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01713 vss n565 n566 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01712 n565 bsrmux_0_shr n554 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01711 n554 in_d_3 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01710 vss n619 n622 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01709 n622 n619 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01708 vss n606 bsrmux_0_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01707 bsrmux_0_f1 n606 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01706 vss n619 n622 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01705 vss n617 n619 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01704 n618 in_d_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01703 n617 bsrmux_0_shr n618 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01702 vss n606 bsrmux_0_f1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01701 vss n605 n606 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01700 n605 bsrmux_0_shr n596 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01699 n596 in_d_1 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01698 n681 bshmatr_0_comr0 bsm_0_15_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01697 bsrmux_15_f1 bshmatr_0_comr0 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01696 n676 bshmatr_0_comr0 bsoout_14_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01695 bsrmux_14_f1 bshmatr_0_comr0 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01694 n673 bshmatr_0_comr0 bsoout_13_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01693 bsrmux_13_f1 bshmatr_0_comr0 bsoout_13_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01692 n671 bshmatr_0_comr0 bsm_0_12_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01691 bsrmux_12_f1 bshmatr_0_comr0 bsoout_12_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01690 n666 bshmatr_0_comr0 bsm_0_11_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01689 bsrmux_11_f1 bshmatr_0_comr0 bsoout_11_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01688 n662 bshmatr_0_comr0 bsm_0_10_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01687 bsrmux_10_f1 bshmatr_0_comr0 bsoout_10_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01686 n656 bshmatr_0_comr0 bsm_0_9_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01685 bsrmux_9_f1 bshmatr_0_comr0 bsoout_9_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01684 n653 bshmatr_0_comr0 bsoout_8_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01683 bsrmux_8_f1 bshmatr_0_comr0 bsoout_8_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01682 n652 bshmatr_0_comr0 bsm_0_7_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01681 bsrmux_7_f1 bshmatr_0_comr0 bsoout_7_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01680 n646 bshmatr_0_comr0 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01679 bsrmux_6_f1 bshmatr_0_comr0 bsoout_6_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01678 n641 bshmatr_0_comr0 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01677 bsrmux_5_f1 bshmatr_0_comr0 bsoout_5_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01676 n636 bshmatr_0_comr0 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01675 bsrmux_4_f1 bshmatr_0_comr0 bsoout_4_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01674 n633 bshmatr_0_comr0 bsoout_3_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01673 bsrmux_3_f1 bshmatr_0_comr0 bsoout_3_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01672 n632 bshmatr_0_comr0 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01671 bsrmux_2_f1 bshmatr_0_comr0 bsoout_2_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01670 n627 bshmatr_0_comr0 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01669 bsrmux_1_f1 bshmatr_0_comr0 bsoout_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01668 n622 bshmatr_0_comr0 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01667 bsrmux_0_f1 bshmatr_0_comr0 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01666 bsoout_15_out_1_s bssnbl_1_out_1 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01665 bslmux_0_out_2 bssnbl_0_out_1 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01664 bsm_0_15_out_2_s bssnbl_1_out_1 bslmux_0_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01663 bsrmux_15_f1 bssnbl_0_out_1 bsm_0_15_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01662 bsoout_14_out_1_s bssnbl_1_out_1 bsrmux_15_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01661 n681 bssnbl_0_out_1 bsoout_14_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01660 bsoout_14_out_2_s bssnbl_1_out_1 n681 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01659 bsrmux_14_f1 bssnbl_0_out_1 bsoout_14_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01658 bsoout_13_out_1_s bssnbl_1_out_1 bsrmux_14_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01657 n676 bssnbl_0_out_1 bsoout_13_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01656 bsoout_13_out_2_s bssnbl_1_out_1 n676 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01655 bsrmux_13_f1 bssnbl_0_out_1 bsoout_13_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01654 bsoout_12_out_1_s bssnbl_1_out_1 bsrmux_13_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01653 n673 bssnbl_0_out_1 bsoout_12_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01652 bsm_0_12_out_2_s bssnbl_1_out_1 n673 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01651 bsrmux_12_f1 bssnbl_0_out_1 bsm_0_12_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01650 bsoout_11_out_1_s bssnbl_1_out_1 bsrmux_12_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01649 n671 bssnbl_0_out_1 bsoout_11_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01648 bsm_0_11_out_2_s bssnbl_1_out_1 n671 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01647 bsrmux_11_f1 bssnbl_0_out_1 bsm_0_11_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01646 bsoout_10_out_1_s bssnbl_1_out_1 bsrmux_11_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01645 n666 bssnbl_0_out_1 bsoout_10_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01644 bsm_0_10_out_2_s bssnbl_1_out_1 n666 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01643 bsrmux_10_f1 bssnbl_0_out_1 bsm_0_10_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01642 bsoout_9_out_1_s bssnbl_1_out_1 bsrmux_10_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01641 n662 bssnbl_0_out_1 bsoout_9_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01640 bsm_0_9_out_2_s bssnbl_1_out_1 n662 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01639 bsrmux_9_f1 bssnbl_0_out_1 bsm_0_9_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01638 bsoout_8_out_1_s bssnbl_1_out_1 bsrmux_9_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01637 n656 bssnbl_0_out_1 bsoout_8_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01636 bsoout_8_out_2_s bssnbl_1_out_1 n656 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01635 bsrmux_8_f1 bssnbl_0_out_1 bsoout_8_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01634 bsoout_7_out_1_s bssnbl_1_out_1 bsrmux_8_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01633 n653 bssnbl_0_out_1 bsoout_7_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01632 bsm_0_7_out_2_s bssnbl_1_out_1 n653 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01631 bsrmux_7_f1 bssnbl_0_out_1 bsm_0_7_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01630 bsoout_6_out_1_s bssnbl_1_out_1 bsrmux_7_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01629 n652 bssnbl_0_out_1 bsoout_6_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01628 bsm_0_6_out_2_s bssnbl_1_out_1 n652 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01627 bsrmux_6_f1 bssnbl_0_out_1 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01626 bsoout_5_out_1_s bssnbl_1_out_1 bsrmux_6_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01625 n646 bssnbl_0_out_1 bsoout_5_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01624 bsm_0_5_out_2_s bssnbl_1_out_1 n646 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01623 bsrmux_5_f1 bssnbl_0_out_1 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01622 bsoout_4_out_1_s bssnbl_1_out_1 bsrmux_5_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01621 n641 bssnbl_0_out_1 bsoout_4_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01620 bsm_0_4_out_2_s bssnbl_1_out_1 n641 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01619 bsrmux_4_f1 bssnbl_0_out_1 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01618 bsoout_3_out_1_s bssnbl_1_out_1 bsrmux_4_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01617 n636 bssnbl_0_out_1 bsoout_3_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01616 bsoout_3_out_2_s bssnbl_1_out_1 n636 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01615 bsrmux_3_f1 bssnbl_0_out_1 bsoout_3_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01614 bsoout_2_out_1_s bssnbl_1_out_1 bsrmux_3_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01613 n633 bssnbl_0_out_1 bsoout_2_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01612 bsm_0_2_out_2_s bssnbl_1_out_1 n633 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01611 bsrmux_2_f1 bssnbl_0_out_1 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01610 bsoout_1_out_1_s bssnbl_1_out_1 bsrmux_2_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01609 n632 bssnbl_0_out_1 bsoout_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01608 bsm_0_1_out_2_s bssnbl_1_out_1 n632 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01607 bsrmux_1_f1 bssnbl_0_out_1 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01606 bsoout_0_out_1_s bssnbl_1_out_1 bsrmux_1_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01605 n627 bssnbl_0_out_1 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01604 bsm_0_0_out_2_s bssnbl_1_out_1 n627 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01603 bsrmux_0_f1 bssnbl_0_out_1 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01602 bsoout_15_out_1_s bssnbl_3_out_1 bslmux_1_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01601 bslmux_1_out_2 bssnbl_2_out_1 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01600 bsm_0_15_out_2_s bssnbl_3_out_1 bslmux_1_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01599 bslmux_0_out_1 bssnbl_2_out_1 bsm_0_15_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01598 bsoout_14_out_1_s bssnbl_3_out_1 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01597 bslmux_0_out_2 bssnbl_2_out_1 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01596 bsoout_14_out_2_s bssnbl_3_out_1 bslmux_0_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01595 bsrmux_15_f1 bssnbl_2_out_1 bsoout_14_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01594 bsoout_13_out_1_s bssnbl_3_out_1 bsrmux_15_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01593 n681 bssnbl_2_out_1 bsoout_13_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01592 bsoout_13_out_2_s bssnbl_3_out_1 n681 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01591 bsrmux_14_f1 bssnbl_2_out_1 bsoout_13_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01590 bsoout_12_out_1_s bssnbl_3_out_1 bsrmux_14_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01589 n676 bssnbl_2_out_1 bsoout_12_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01588 bsm_0_12_out_2_s bssnbl_3_out_1 n676 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01587 bsrmux_13_f1 bssnbl_2_out_1 bsm_0_12_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01586 bsoout_11_out_1_s bssnbl_3_out_1 bsrmux_13_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01585 n673 bssnbl_2_out_1 bsoout_11_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01584 bsm_0_11_out_2_s bssnbl_3_out_1 n673 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01583 bsrmux_12_f1 bssnbl_2_out_1 bsm_0_11_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01582 bsoout_10_out_1_s bssnbl_3_out_1 bsrmux_12_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01581 n671 bssnbl_2_out_1 bsoout_10_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01580 bsm_0_10_out_2_s bssnbl_3_out_1 n671 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01579 bsrmux_11_f1 bssnbl_2_out_1 bsm_0_10_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01578 bsoout_9_out_1_s bssnbl_3_out_1 bsrmux_11_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01577 n666 bssnbl_2_out_1 bsoout_9_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01576 bsm_0_9_out_2_s bssnbl_3_out_1 n666 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01575 bsrmux_10_f1 bssnbl_2_out_1 bsm_0_9_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01574 bsoout_8_out_1_s bssnbl_3_out_1 bsrmux_10_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01573 n662 bssnbl_2_out_1 bsoout_8_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01572 bsoout_8_out_2_s bssnbl_3_out_1 n662 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01571 bsrmux_9_f1 bssnbl_2_out_1 bsoout_8_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01570 bsoout_7_out_1_s bssnbl_3_out_1 bsrmux_9_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01569 n656 bssnbl_2_out_1 bsoout_7_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01568 bsm_0_7_out_2_s bssnbl_3_out_1 n656 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01567 bsrmux_8_f1 bssnbl_2_out_1 bsm_0_7_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01566 bsoout_6_out_1_s bssnbl_3_out_1 bsrmux_8_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01565 n653 bssnbl_2_out_1 bsoout_6_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01564 bsm_0_6_out_2_s bssnbl_3_out_1 n653 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01563 bsrmux_7_f1 bssnbl_2_out_1 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01562 bsoout_5_out_1_s bssnbl_3_out_1 bsrmux_7_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01561 n652 bssnbl_2_out_1 bsoout_5_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01560 bsm_0_5_out_2_s bssnbl_3_out_1 n652 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01559 bsrmux_6_f1 bssnbl_2_out_1 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01558 bsoout_4_out_1_s bssnbl_3_out_1 bsrmux_6_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01557 n646 bssnbl_2_out_1 bsoout_4_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01556 bsm_0_4_out_2_s bssnbl_3_out_1 n646 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01555 bsrmux_5_f1 bssnbl_2_out_1 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01554 bsoout_3_out_1_s bssnbl_3_out_1 bsrmux_5_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01553 n641 bssnbl_2_out_1 bsoout_3_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01552 bsoout_3_out_2_s bssnbl_3_out_1 n641 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01551 bsrmux_4_f1 bssnbl_2_out_1 bsoout_3_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01550 bsoout_2_out_1_s bssnbl_3_out_1 bsrmux_4_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01549 n636 bssnbl_2_out_1 bsoout_2_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01548 bsm_0_2_out_2_s bssnbl_3_out_1 n636 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01547 bsrmux_3_f1 bssnbl_2_out_1 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01546 bsoout_1_out_1_s bssnbl_3_out_1 bsrmux_3_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01545 n633 bssnbl_2_out_1 bsoout_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01544 bsm_0_1_out_2_s bssnbl_3_out_1 n633 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01543 bsrmux_2_f1 bssnbl_2_out_1 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01542 bsoout_0_out_1_s bssnbl_3_out_1 bsrmux_2_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01541 n632 bssnbl_2_out_1 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01540 bsm_0_0_out_2_s bssnbl_3_out_1 n632 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01539 bsrmux_1_f1 bssnbl_2_out_1 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01538 bsoout_15_out_1_s bssnbl_5_out_1 bslmux_2_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01537 bslmux_2_out_2 bssnbl_4_out_1 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01536 bsm_0_15_out_2_s bssnbl_5_out_1 bslmux_2_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01535 bslmux_1_out_1 bssnbl_4_out_1 bsm_0_15_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01534 bsoout_14_out_1_s bssnbl_5_out_1 bslmux_1_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01533 bslmux_1_out_2 bssnbl_4_out_1 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01532 bsoout_14_out_2_s bssnbl_5_out_1 bslmux_1_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01531 bslmux_0_out_1 bssnbl_4_out_1 bsoout_14_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01530 bsoout_13_out_1_s bssnbl_5_out_1 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01529 bslmux_0_out_2 bssnbl_4_out_1 bsoout_13_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01528 bsoout_13_out_2_s bssnbl_5_out_1 bslmux_0_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01527 bsrmux_15_f1 bssnbl_4_out_1 bsoout_13_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01526 bsoout_12_out_1_s bssnbl_5_out_1 bsrmux_15_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01525 n681 bssnbl_4_out_1 bsoout_12_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01524 bsm_0_12_out_2_s bssnbl_5_out_1 n681 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01523 bsrmux_14_f1 bssnbl_4_out_1 bsm_0_12_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01522 bsoout_11_out_1_s bssnbl_5_out_1 bsrmux_14_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01521 n676 bssnbl_4_out_1 bsoout_11_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01520 bsm_0_11_out_2_s bssnbl_5_out_1 n676 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01519 bsrmux_13_f1 bssnbl_4_out_1 bsm_0_11_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01518 bsoout_10_out_1_s bssnbl_5_out_1 bsrmux_13_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01517 n673 bssnbl_4_out_1 bsoout_10_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01516 bsm_0_10_out_2_s bssnbl_5_out_1 n673 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01515 bsrmux_12_f1 bssnbl_4_out_1 bsm_0_10_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01514 bsoout_9_out_1_s bssnbl_5_out_1 bsrmux_12_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01513 n671 bssnbl_4_out_1 bsoout_9_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01512 bsm_0_9_out_2_s bssnbl_5_out_1 n671 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01511 bsrmux_11_f1 bssnbl_4_out_1 bsm_0_9_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01510 bsoout_8_out_1_s bssnbl_5_out_1 bsrmux_11_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01509 n666 bssnbl_4_out_1 bsoout_8_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01508 bsoout_8_out_2_s bssnbl_5_out_1 n666 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01507 bsrmux_10_f1 bssnbl_4_out_1 bsoout_8_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01506 bsoout_7_out_1_s bssnbl_5_out_1 bsrmux_10_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01505 n662 bssnbl_4_out_1 bsoout_7_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01504 bsm_0_7_out_2_s bssnbl_5_out_1 n662 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01503 bsrmux_9_f1 bssnbl_4_out_1 bsm_0_7_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01502 bsoout_6_out_1_s bssnbl_5_out_1 bsrmux_9_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01501 n656 bssnbl_4_out_1 bsoout_6_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01500 bsm_0_6_out_2_s bssnbl_5_out_1 n656 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01499 bsrmux_8_f1 bssnbl_4_out_1 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01498 bsoout_5_out_1_s bssnbl_5_out_1 bsrmux_8_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01497 n653 bssnbl_4_out_1 bsoout_5_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01496 bsm_0_5_out_2_s bssnbl_5_out_1 n653 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01495 bsrmux_7_f1 bssnbl_4_out_1 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01494 bsoout_4_out_1_s bssnbl_5_out_1 bsrmux_7_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01493 n652 bssnbl_4_out_1 bsoout_4_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01492 bsm_0_4_out_2_s bssnbl_5_out_1 n652 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01491 bsrmux_6_f1 bssnbl_4_out_1 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01490 bsoout_3_out_1_s bssnbl_5_out_1 bsrmux_6_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01489 n646 bssnbl_4_out_1 bsoout_3_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01488 bsoout_3_out_2_s bssnbl_5_out_1 n646 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01487 bsrmux_5_f1 bssnbl_4_out_1 bsoout_3_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01486 bsoout_2_out_1_s bssnbl_5_out_1 bsrmux_5_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01485 n641 bssnbl_4_out_1 bsoout_2_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01484 bsm_0_2_out_2_s bssnbl_5_out_1 n641 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01483 bsrmux_4_f1 bssnbl_4_out_1 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01482 bsoout_1_out_1_s bssnbl_5_out_1 bsrmux_4_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01481 n636 bssnbl_4_out_1 bsoout_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01480 bsm_0_1_out_2_s bssnbl_5_out_1 n636 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01479 bsrmux_3_f1 bssnbl_4_out_1 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01478 bsoout_0_out_1_s bssnbl_5_out_1 bsrmux_3_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01477 n633 bssnbl_4_out_1 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01476 bsm_0_0_out_2_s bssnbl_5_out_1 n633 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01475 bsrmux_2_f1 bssnbl_4_out_1 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01474 bsoout_15_out_1_s bssnbl_7_out_1 bslmux_3_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01473 bslmux_3_out_2 bssnbl_6_out_1 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01472 bsm_0_15_out_2_s bssnbl_7_out_1 bslmux_3_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01471 bslmux_2_out_1 bssnbl_6_out_1 bsm_0_15_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01470 bsoout_14_out_1_s bssnbl_7_out_1 bslmux_2_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01469 bslmux_2_out_2 bssnbl_6_out_1 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01468 bsoout_14_out_2_s bssnbl_7_out_1 bslmux_2_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01467 bslmux_1_out_1 bssnbl_6_out_1 bsoout_14_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01466 bsoout_13_out_1_s bssnbl_7_out_1 bslmux_1_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01465 bslmux_1_out_2 bssnbl_6_out_1 bsoout_13_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01464 bsoout_13_out_2_s bssnbl_7_out_1 bslmux_1_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01463 bslmux_0_out_1 bssnbl_6_out_1 bsoout_13_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01462 bsoout_12_out_1_s bssnbl_7_out_1 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01461 bslmux_0_out_2 bssnbl_6_out_1 bsoout_12_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01460 bsm_0_12_out_2_s bssnbl_7_out_1 bslmux_0_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01459 bsrmux_15_f1 bssnbl_6_out_1 bsm_0_12_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01458 bsoout_11_out_1_s bssnbl_7_out_1 bsrmux_15_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01457 n681 bssnbl_6_out_1 bsoout_11_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01456 bsm_0_11_out_2_s bssnbl_7_out_1 n681 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01455 bsrmux_14_f1 bssnbl_6_out_1 bsm_0_11_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01454 bsoout_10_out_1_s bssnbl_7_out_1 bsrmux_14_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01453 n676 bssnbl_6_out_1 bsoout_10_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01452 bsm_0_10_out_2_s bssnbl_7_out_1 n676 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01451 bsrmux_13_f1 bssnbl_6_out_1 bsm_0_10_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01450 bsoout_9_out_1_s bssnbl_7_out_1 bsrmux_13_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01449 n673 bssnbl_6_out_1 bsoout_9_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01448 bsm_0_9_out_2_s bssnbl_7_out_1 n673 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01447 bsrmux_12_f1 bssnbl_6_out_1 bsm_0_9_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01446 bsoout_8_out_1_s bssnbl_7_out_1 bsrmux_12_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01445 n671 bssnbl_6_out_1 bsoout_8_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01444 bsoout_8_out_2_s bssnbl_7_out_1 n671 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01443 bsrmux_11_f1 bssnbl_6_out_1 bsoout_8_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01442 bsoout_7_out_1_s bssnbl_7_out_1 bsrmux_11_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01441 n666 bssnbl_6_out_1 bsoout_7_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01440 bsm_0_7_out_2_s bssnbl_7_out_1 n666 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01439 bsrmux_10_f1 bssnbl_6_out_1 bsm_0_7_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01438 bsoout_6_out_1_s bssnbl_7_out_1 bsrmux_10_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01437 n662 bssnbl_6_out_1 bsoout_6_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01436 bsm_0_6_out_2_s bssnbl_7_out_1 n662 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01435 bsrmux_9_f1 bssnbl_6_out_1 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01434 bsoout_5_out_1_s bssnbl_7_out_1 bsrmux_9_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01433 n656 bssnbl_6_out_1 bsoout_5_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01432 bsm_0_5_out_2_s bssnbl_7_out_1 n656 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01431 bsrmux_8_f1 bssnbl_6_out_1 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01430 bsoout_4_out_1_s bssnbl_7_out_1 bsrmux_8_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01429 n653 bssnbl_6_out_1 bsoout_4_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01428 bsm_0_4_out_2_s bssnbl_7_out_1 n653 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01427 bsrmux_7_f1 bssnbl_6_out_1 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01426 bsoout_3_out_1_s bssnbl_7_out_1 bsrmux_7_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01425 n652 bssnbl_6_out_1 bsoout_3_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01424 bsoout_3_out_2_s bssnbl_7_out_1 n652 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01423 bsrmux_6_f1 bssnbl_6_out_1 bsoout_3_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01422 bsoout_2_out_1_s bssnbl_7_out_1 bsrmux_6_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01421 n646 bssnbl_6_out_1 bsoout_2_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01420 bsm_0_2_out_2_s bssnbl_7_out_1 n646 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01419 bsrmux_5_f1 bssnbl_6_out_1 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01418 bsoout_1_out_1_s bssnbl_7_out_1 bsrmux_5_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01417 n641 bssnbl_6_out_1 bsoout_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01416 bsm_0_1_out_2_s bssnbl_7_out_1 n641 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01415 bsrmux_4_f1 bssnbl_6_out_1 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01414 bsoout_0_out_1_s bssnbl_7_out_1 bsrmux_4_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01413 n636 bssnbl_6_out_1 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01412 bsm_0_0_out_2_s bssnbl_7_out_1 n636 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01411 bsrmux_3_f1 bssnbl_6_out_1 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01410 bsoout_15_out_1_s bssnbl_9_out_1 bslmux_4_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01409 bslmux_4_out_2 bssnbl_8_out_1 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01408 bsm_0_15_out_2_s bssnbl_9_out_1 bslmux_4_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01407 bslmux_3_out_1 bssnbl_8_out_1 bsm_0_15_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01406 bsoout_14_out_1_s bssnbl_9_out_1 bslmux_3_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01405 bslmux_3_out_2 bssnbl_8_out_1 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01404 bsoout_14_out_2_s bssnbl_9_out_1 bslmux_3_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01403 bslmux_2_out_1 bssnbl_8_out_1 bsoout_14_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01402 bsoout_13_out_1_s bssnbl_9_out_1 bslmux_2_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01401 bslmux_2_out_2 bssnbl_8_out_1 bsoout_13_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01400 bsoout_13_out_2_s bssnbl_9_out_1 bslmux_2_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01399 bslmux_1_out_1 bssnbl_8_out_1 bsoout_13_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01398 bsoout_12_out_1_s bssnbl_9_out_1 bslmux_1_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01397 bslmux_1_out_2 bssnbl_8_out_1 bsoout_12_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01396 bsm_0_12_out_2_s bssnbl_9_out_1 bslmux_1_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01395 bslmux_0_out_1 bssnbl_8_out_1 bsm_0_12_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01394 bsoout_11_out_1_s bssnbl_9_out_1 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01393 bslmux_0_out_2 bssnbl_8_out_1 bsoout_11_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01392 bsm_0_11_out_2_s bssnbl_9_out_1 bslmux_0_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01391 bsrmux_15_f1 bssnbl_8_out_1 bsm_0_11_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01390 bsoout_10_out_1_s bssnbl_9_out_1 bsrmux_15_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01389 n681 bssnbl_8_out_1 bsoout_10_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01388 bsm_0_10_out_2_s bssnbl_9_out_1 n681 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01387 bsrmux_14_f1 bssnbl_8_out_1 bsm_0_10_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01386 bsoout_9_out_1_s bssnbl_9_out_1 bsrmux_14_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01385 n676 bssnbl_8_out_1 bsoout_9_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01384 bsm_0_9_out_2_s bssnbl_9_out_1 n676 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01383 bsrmux_13_f1 bssnbl_8_out_1 bsm_0_9_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01382 bsoout_8_out_1_s bssnbl_9_out_1 bsrmux_13_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01381 n673 bssnbl_8_out_1 bsoout_8_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01380 bsoout_8_out_2_s bssnbl_9_out_1 n673 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01379 bsrmux_12_f1 bssnbl_8_out_1 bsoout_8_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01378 bsoout_7_out_1_s bssnbl_9_out_1 bsrmux_12_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01377 n671 bssnbl_8_out_1 bsoout_7_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01376 bsm_0_7_out_2_s bssnbl_9_out_1 n671 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01375 bsrmux_11_f1 bssnbl_8_out_1 bsm_0_7_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01374 bsoout_6_out_1_s bssnbl_9_out_1 bsrmux_11_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01373 n666 bssnbl_8_out_1 bsoout_6_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01372 bsm_0_6_out_2_s bssnbl_9_out_1 n666 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01371 bsrmux_10_f1 bssnbl_8_out_1 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01370 bsoout_5_out_1_s bssnbl_9_out_1 bsrmux_10_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01369 n662 bssnbl_8_out_1 bsoout_5_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01368 bsm_0_5_out_2_s bssnbl_9_out_1 n662 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01367 bsrmux_9_f1 bssnbl_8_out_1 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01366 bsoout_4_out_1_s bssnbl_9_out_1 bsrmux_9_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01365 n656 bssnbl_8_out_1 bsoout_4_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01364 bsm_0_4_out_2_s bssnbl_9_out_1 n656 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01363 bsrmux_8_f1 bssnbl_8_out_1 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01362 bsoout_3_out_1_s bssnbl_9_out_1 bsrmux_8_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01361 n653 bssnbl_8_out_1 bsoout_3_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01360 bsoout_3_out_2_s bssnbl_9_out_1 n653 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01359 bsrmux_7_f1 bssnbl_8_out_1 bsoout_3_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01358 bsoout_2_out_1_s bssnbl_9_out_1 bsrmux_7_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01357 n652 bssnbl_8_out_1 bsoout_2_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01356 bsm_0_2_out_2_s bssnbl_9_out_1 n652 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01355 bsrmux_6_f1 bssnbl_8_out_1 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01354 bsoout_1_out_1_s bssnbl_9_out_1 bsrmux_6_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01353 n646 bssnbl_8_out_1 bsoout_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01352 bsm_0_1_out_2_s bssnbl_9_out_1 n646 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01351 bsrmux_5_f1 bssnbl_8_out_1 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01350 bsoout_0_out_1_s bssnbl_9_out_1 bsrmux_5_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01349 n641 bssnbl_8_out_1 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01348 bsm_0_0_out_2_s bssnbl_9_out_1 n641 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01347 bsrmux_4_f1 bssnbl_8_out_1 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01346 bsoout_15_out_1_s bssnbl_11_out_1 bslmux_5_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01345 bslmux_5_out_2 bssnbl_10_out_1 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01344 bsm_0_15_out_2_s bssnbl_11_out_1 bslmux_5_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01343 bslmux_4_out_1 bssnbl_10_out_1 bsm_0_15_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01342 bsoout_14_out_1_s bssnbl_11_out_1 bslmux_4_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01341 bslmux_4_out_2 bssnbl_10_out_1 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01340 bsoout_14_out_2_s bssnbl_11_out_1 bslmux_4_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01339 bslmux_3_out_1 bssnbl_10_out_1 bsoout_14_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01338 bsoout_13_out_1_s bssnbl_11_out_1 bslmux_3_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01337 bslmux_3_out_2 bssnbl_10_out_1 bsoout_13_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01336 bsoout_13_out_2_s bssnbl_11_out_1 bslmux_3_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01335 bslmux_2_out_1 bssnbl_10_out_1 bsoout_13_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01334 bsoout_12_out_1_s bssnbl_11_out_1 bslmux_2_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01333 bslmux_2_out_2 bssnbl_10_out_1 bsoout_12_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01332 bsm_0_12_out_2_s bssnbl_11_out_1 bslmux_2_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01331 bslmux_1_out_1 bssnbl_10_out_1 bsm_0_12_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01330 bsoout_11_out_1_s bssnbl_11_out_1 bslmux_1_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01329 bslmux_1_out_2 bssnbl_10_out_1 bsoout_11_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01328 bsm_0_11_out_2_s bssnbl_11_out_1 bslmux_1_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01327 bslmux_0_out_1 bssnbl_10_out_1 bsm_0_11_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01326 bsoout_10_out_1_s bssnbl_11_out_1 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01325 bslmux_0_out_2 bssnbl_10_out_1 bsoout_10_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01324 bsm_0_10_out_2_s bssnbl_11_out_1 bslmux_0_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01323 bsrmux_15_f1 bssnbl_10_out_1 bsm_0_10_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01322 bsoout_9_out_1_s bssnbl_11_out_1 bsrmux_15_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01321 n681 bssnbl_10_out_1 bsoout_9_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01320 bsm_0_9_out_2_s bssnbl_11_out_1 n681 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01319 bsrmux_14_f1 bssnbl_10_out_1 bsm_0_9_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01318 bsoout_8_out_1_s bssnbl_11_out_1 bsrmux_14_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01317 n676 bssnbl_10_out_1 bsoout_8_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01316 bsoout_8_out_2_s bssnbl_11_out_1 n676 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01315 bsrmux_13_f1 bssnbl_10_out_1 bsoout_8_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01314 bsoout_7_out_1_s bssnbl_11_out_1 bsrmux_13_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01313 n673 bssnbl_10_out_1 bsoout_7_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01312 bsm_0_7_out_2_s bssnbl_11_out_1 n673 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01311 bsrmux_12_f1 bssnbl_10_out_1 bsm_0_7_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01310 bsoout_6_out_1_s bssnbl_11_out_1 bsrmux_12_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01309 n671 bssnbl_10_out_1 bsoout_6_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01308 bsm_0_6_out_2_s bssnbl_11_out_1 n671 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01307 bsrmux_11_f1 bssnbl_10_out_1 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01306 bsoout_5_out_1_s bssnbl_11_out_1 bsrmux_11_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01305 n666 bssnbl_10_out_1 bsoout_5_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01304 bsm_0_5_out_2_s bssnbl_11_out_1 n666 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01303 bsrmux_10_f1 bssnbl_10_out_1 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01302 bsoout_4_out_1_s bssnbl_11_out_1 bsrmux_10_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01301 n662 bssnbl_10_out_1 bsoout_4_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01300 bsm_0_4_out_2_s bssnbl_11_out_1 n662 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01299 bsrmux_9_f1 bssnbl_10_out_1 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01298 bsoout_3_out_1_s bssnbl_11_out_1 bsrmux_9_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01297 n656 bssnbl_10_out_1 bsoout_3_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01296 bsoout_3_out_2_s bssnbl_11_out_1 n656 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01295 bsrmux_8_f1 bssnbl_10_out_1 bsoout_3_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01294 bsoout_2_out_1_s bssnbl_11_out_1 bsrmux_8_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01293 n653 bssnbl_10_out_1 bsoout_2_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01292 bsm_0_2_out_2_s bssnbl_11_out_1 n653 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01291 bsrmux_7_f1 bssnbl_10_out_1 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01290 bsoout_1_out_1_s bssnbl_11_out_1 bsrmux_7_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01289 n652 bssnbl_10_out_1 bsoout_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01288 bsm_0_1_out_2_s bssnbl_11_out_1 n652 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01287 bsrmux_6_f1 bssnbl_10_out_1 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01286 bsoout_0_out_1_s bssnbl_11_out_1 bsrmux_6_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01285 n646 bssnbl_10_out_1 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01284 bsm_0_0_out_2_s bssnbl_11_out_1 n646 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01283 bsrmux_5_f1 bssnbl_10_out_1 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01282 bsoout_15_out_1_s bssnbl_13_out_1 bslmux_6_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01281 bslmux_6_out_2 bssnbl_12_out_1 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01280 bsm_0_15_out_2_s bssnbl_13_out_1 bslmux_6_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01279 bslmux_5_out_1 bssnbl_12_out_1 bsm_0_15_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01278 bsoout_14_out_1_s bssnbl_13_out_1 bslmux_5_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01277 bslmux_5_out_2 bssnbl_12_out_1 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01276 bsoout_14_out_2_s bssnbl_13_out_1 bslmux_5_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01275 bslmux_4_out_1 bssnbl_12_out_1 bsoout_14_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01274 bsoout_13_out_1_s bssnbl_13_out_1 bslmux_4_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01273 bslmux_4_out_2 bssnbl_12_out_1 bsoout_13_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01272 bsoout_13_out_2_s bssnbl_13_out_1 bslmux_4_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01271 bslmux_3_out_1 bssnbl_12_out_1 bsoout_13_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01270 bsoout_12_out_1_s bssnbl_13_out_1 bslmux_3_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01269 bslmux_3_out_2 bssnbl_12_out_1 bsoout_12_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01268 bsm_0_12_out_2_s bssnbl_13_out_1 bslmux_3_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01267 bslmux_2_out_1 bssnbl_12_out_1 bsm_0_12_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01266 bsoout_11_out_1_s bssnbl_13_out_1 bslmux_2_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01265 bslmux_2_out_2 bssnbl_12_out_1 bsoout_11_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01264 bsm_0_11_out_2_s bssnbl_13_out_1 bslmux_2_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01263 bslmux_1_out_1 bssnbl_12_out_1 bsm_0_11_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01262 bsoout_10_out_1_s bssnbl_13_out_1 bslmux_1_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01261 bslmux_1_out_2 bssnbl_12_out_1 bsoout_10_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01260 bsm_0_10_out_2_s bssnbl_13_out_1 bslmux_1_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01259 bslmux_0_out_1 bssnbl_12_out_1 bsm_0_10_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01258 bsoout_9_out_1_s bssnbl_13_out_1 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01257 bslmux_0_out_2 bssnbl_12_out_1 bsoout_9_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01256 bsm_0_9_out_2_s bssnbl_13_out_1 bslmux_0_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01255 bsrmux_15_f1 bssnbl_12_out_1 bsm_0_9_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01254 bsoout_8_out_1_s bssnbl_13_out_1 bsrmux_15_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01253 n681 bssnbl_12_out_1 bsoout_8_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01252 bsoout_8_out_2_s bssnbl_13_out_1 n681 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01251 bsrmux_14_f1 bssnbl_12_out_1 bsoout_8_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01250 bsoout_7_out_1_s bssnbl_13_out_1 bsrmux_14_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01249 n676 bssnbl_12_out_1 bsoout_7_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01248 bsm_0_7_out_2_s bssnbl_13_out_1 n676 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01247 bsrmux_13_f1 bssnbl_12_out_1 bsm_0_7_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01246 bsoout_6_out_1_s bssnbl_13_out_1 bsrmux_13_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01245 n673 bssnbl_12_out_1 bsoout_6_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01244 bsm_0_6_out_2_s bssnbl_13_out_1 n673 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01243 bsrmux_12_f1 bssnbl_12_out_1 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01242 bsoout_5_out_1_s bssnbl_13_out_1 bsrmux_12_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01241 n671 bssnbl_12_out_1 bsoout_5_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01240 bsm_0_5_out_2_s bssnbl_13_out_1 n671 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01239 bsrmux_11_f1 bssnbl_12_out_1 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01238 bsoout_4_out_1_s bssnbl_13_out_1 bsrmux_11_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01237 n666 bssnbl_12_out_1 bsoout_4_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01236 bsm_0_4_out_2_s bssnbl_13_out_1 n666 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01235 bsrmux_10_f1 bssnbl_12_out_1 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01234 bsoout_3_out_1_s bssnbl_13_out_1 bsrmux_10_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01233 n662 bssnbl_12_out_1 bsoout_3_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01232 bsoout_3_out_2_s bssnbl_13_out_1 n662 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01231 bsrmux_9_f1 bssnbl_12_out_1 bsoout_3_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01230 bsoout_2_out_1_s bssnbl_13_out_1 bsrmux_9_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01229 n656 bssnbl_12_out_1 bsoout_2_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01228 bsm_0_2_out_2_s bssnbl_13_out_1 n656 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01227 bsrmux_8_f1 bssnbl_12_out_1 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01226 bsoout_1_out_1_s bssnbl_13_out_1 bsrmux_8_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01225 n653 bssnbl_12_out_1 bsoout_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01224 bsm_0_1_out_2_s bssnbl_13_out_1 n653 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01223 bsrmux_7_f1 bssnbl_12_out_1 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01222 bsoout_0_out_1_s bssnbl_13_out_1 bsrmux_7_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01221 n652 bssnbl_12_out_1 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01220 bsm_0_0_out_2_s bssnbl_13_out_1 n652 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01219 bsrmux_6_f1 bssnbl_12_out_1 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01218 bsoout_15_out_1_s bslmux_15_com_2 bslmux_7_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01217 bslmux_7_out_2 bssnbl_14_out_1 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01216 bsm_0_15_out_2_s bslmux_15_com_2 bslmux_7_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01215 bslmux_6_out_1 bssnbl_14_out_1 bsm_0_15_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01214 bsoout_14_out_1_s bslmux_15_com_2 bslmux_6_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01213 bslmux_6_out_2 bssnbl_14_out_1 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01212 bsoout_14_out_2_s bslmux_15_com_2 bslmux_6_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01211 bslmux_5_out_1 bssnbl_14_out_1 bsoout_14_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01210 bsoout_13_out_1_s bslmux_15_com_2 bslmux_5_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01209 bslmux_5_out_2 bssnbl_14_out_1 bsoout_13_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01208 bsoout_13_out_2_s bslmux_15_com_2 bslmux_5_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01207 bslmux_4_out_1 bssnbl_14_out_1 bsoout_13_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01206 bsoout_12_out_1_s bslmux_15_com_2 bslmux_4_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01205 bslmux_4_out_2 bssnbl_14_out_1 bsoout_12_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01204 bsm_0_12_out_2_s bslmux_15_com_2 bslmux_4_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01203 bslmux_3_out_1 bssnbl_14_out_1 bsm_0_12_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01202 bsoout_11_out_1_s bslmux_15_com_2 bslmux_3_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01201 bslmux_3_out_2 bssnbl_14_out_1 bsoout_11_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01200 bsm_0_11_out_2_s bslmux_15_com_2 bslmux_3_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01199 bslmux_2_out_1 bssnbl_14_out_1 bsm_0_11_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01198 bsoout_10_out_1_s bslmux_15_com_2 bslmux_2_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01197 bslmux_2_out_2 bssnbl_14_out_1 bsoout_10_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01196 bsm_0_10_out_2_s bslmux_15_com_2 bslmux_2_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01195 bslmux_1_out_1 bssnbl_14_out_1 bsm_0_10_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01194 bsoout_9_out_1_s bslmux_15_com_2 bslmux_1_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01193 bslmux_1_out_2 bssnbl_14_out_1 bsoout_9_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01192 bsm_0_9_out_2_s bslmux_15_com_2 bslmux_1_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01191 bslmux_0_out_1 bssnbl_14_out_1 bsm_0_9_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01190 bsoout_8_out_1_s bslmux_15_com_2 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01189 bslmux_0_out_2 bssnbl_14_out_1 bsoout_8_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01188 bsoout_8_out_2_s bslmux_15_com_2 bslmux_0_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01187 bsrmux_15_f1 bssnbl_14_out_1 bsoout_8_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01186 bsoout_7_out_1_s bslmux_15_com_2 bsrmux_15_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01185 n681 bssnbl_14_out_1 bsoout_7_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01184 bsm_0_7_out_2_s bslmux_15_com_2 n681 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01183 bsrmux_14_f1 bssnbl_14_out_1 bsm_0_7_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01182 bsoout_6_out_1_s bslmux_15_com_2 bsrmux_14_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01181 n676 bssnbl_14_out_1 bsoout_6_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01180 bsm_0_6_out_2_s bslmux_15_com_2 n676 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01179 bsrmux_13_f1 bssnbl_14_out_1 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01178 bsoout_5_out_1_s bslmux_15_com_2 bsrmux_13_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01177 n673 bssnbl_14_out_1 bsoout_5_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01176 bsm_0_5_out_2_s bslmux_15_com_2 n673 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01175 bsrmux_12_f1 bssnbl_14_out_1 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01174 bsoout_4_out_1_s bslmux_15_com_2 bsrmux_12_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01173 n671 bssnbl_14_out_1 bsoout_4_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01172 bsm_0_4_out_2_s bslmux_15_com_2 n671 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01171 bsrmux_11_f1 bssnbl_14_out_1 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01170 bsoout_3_out_1_s bslmux_15_com_2 bsrmux_11_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01169 n666 bssnbl_14_out_1 bsoout_3_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01168 bsoout_3_out_2_s bslmux_15_com_2 n666 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01167 bsrmux_10_f1 bssnbl_14_out_1 bsoout_3_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01166 bsoout_2_out_1_s bslmux_15_com_2 bsrmux_10_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01165 n662 bssnbl_14_out_1 bsoout_2_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01164 bsm_0_2_out_2_s bslmux_15_com_2 n662 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01163 bsrmux_9_f1 bssnbl_14_out_1 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01162 bsoout_1_out_1_s bslmux_15_com_2 bsrmux_9_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01161 n656 bssnbl_14_out_1 bsoout_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01160 bsm_0_1_out_2_s bslmux_15_com_2 n656 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01159 bsrmux_8_f1 bssnbl_14_out_1 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01158 bsoout_0_out_1_s bslmux_15_com_2 bsrmux_8_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01157 n653 bssnbl_14_out_1 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01156 bsm_0_0_out_2_s bslmux_15_com_2 n653 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01155 bsrmux_7_f1 bssnbl_14_out_1 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01154 bsoout_15_out_1_s bslmux_13_com_2 bslmux_8_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01153 bslmux_8_out_2 bslmux_14_com_2 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01152 bsm_0_15_out_2_s bslmux_13_com_2 bslmux_8_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01151 bslmux_7_out_1 bslmux_14_com_2 bsm_0_15_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01150 bsoout_14_out_1_s bslmux_13_com_2 bslmux_7_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01149 bslmux_7_out_2 bslmux_14_com_2 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01148 bsoout_14_out_2_s bslmux_13_com_2 bslmux_7_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01147 bslmux_6_out_1 bslmux_14_com_2 bsoout_14_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01146 bsoout_13_out_1_s bslmux_13_com_2 bslmux_6_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01145 bslmux_6_out_2 bslmux_14_com_2 bsoout_13_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01144 bsoout_13_out_2_s bslmux_13_com_2 bslmux_6_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01143 bslmux_5_out_1 bslmux_14_com_2 bsoout_13_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01142 bsoout_12_out_1_s bslmux_13_com_2 bslmux_5_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01141 bslmux_5_out_2 bslmux_14_com_2 bsoout_12_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01140 bsm_0_12_out_2_s bslmux_13_com_2 bslmux_5_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01139 bslmux_4_out_1 bslmux_14_com_2 bsm_0_12_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01138 bsoout_11_out_1_s bslmux_13_com_2 bslmux_4_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01137 bslmux_4_out_2 bslmux_14_com_2 bsoout_11_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01136 bsm_0_11_out_2_s bslmux_13_com_2 bslmux_4_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01135 bslmux_3_out_1 bslmux_14_com_2 bsm_0_11_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01134 bsoout_10_out_1_s bslmux_13_com_2 bslmux_3_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01133 bslmux_3_out_2 bslmux_14_com_2 bsoout_10_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01132 bsm_0_10_out_2_s bslmux_13_com_2 bslmux_3_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01131 bslmux_2_out_1 bslmux_14_com_2 bsm_0_10_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01130 bsoout_9_out_1_s bslmux_13_com_2 bslmux_2_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01129 bslmux_2_out_2 bslmux_14_com_2 bsoout_9_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01128 bsm_0_9_out_2_s bslmux_13_com_2 bslmux_2_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01127 bslmux_1_out_1 bslmux_14_com_2 bsm_0_9_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01126 bsoout_8_out_1_s bslmux_13_com_2 bslmux_1_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01125 bslmux_1_out_2 bslmux_14_com_2 bsoout_8_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01124 bsoout_8_out_2_s bslmux_13_com_2 bslmux_1_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01123 bslmux_0_out_1 bslmux_14_com_2 bsoout_8_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01122 bsoout_7_out_1_s bslmux_13_com_2 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01121 bslmux_0_out_2 bslmux_14_com_2 bsoout_7_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01120 bsm_0_7_out_2_s bslmux_13_com_2 bslmux_0_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01119 bsrmux_15_f1 bslmux_14_com_2 bsm_0_7_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01118 bsoout_6_out_1_s bslmux_13_com_2 bsrmux_15_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01117 n681 bslmux_14_com_2 bsoout_6_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01116 bsm_0_6_out_2_s bslmux_13_com_2 n681 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01115 bsrmux_14_f1 bslmux_14_com_2 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01114 bsoout_5_out_1_s bslmux_13_com_2 bsrmux_14_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01113 n676 bslmux_14_com_2 bsoout_5_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01112 bsm_0_5_out_2_s bslmux_13_com_2 n676 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01111 bsrmux_13_f1 bslmux_14_com_2 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01110 bsoout_4_out_1_s bslmux_13_com_2 bsrmux_13_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01109 n673 bslmux_14_com_2 bsoout_4_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01108 bsm_0_4_out_2_s bslmux_13_com_2 n673 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01107 bsrmux_12_f1 bslmux_14_com_2 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01106 bsoout_3_out_1_s bslmux_13_com_2 bsrmux_12_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01105 n671 bslmux_14_com_2 bsoout_3_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01104 bsoout_3_out_2_s bslmux_13_com_2 n671 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01103 bsrmux_11_f1 bslmux_14_com_2 bsoout_3_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01102 bsoout_2_out_1_s bslmux_13_com_2 bsrmux_11_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01101 n666 bslmux_14_com_2 bsoout_2_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01100 bsm_0_2_out_2_s bslmux_13_com_2 n666 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01099 bsrmux_10_f1 bslmux_14_com_2 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01098 bsoout_1_out_1_s bslmux_13_com_2 bsrmux_10_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01097 n662 bslmux_14_com_2 bsoout_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01096 bsm_0_1_out_2_s bslmux_13_com_2 n662 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01095 bsrmux_9_f1 bslmux_14_com_2 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01094 bsoout_0_out_1_s bslmux_13_com_2 bsrmux_9_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01093 n656 bslmux_14_com_2 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01092 bsm_0_0_out_2_s bslmux_13_com_2 n656 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01091 bsrmux_8_f1 bslmux_14_com_2 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01090 bsoout_15_out_1_s bslmux_11_com_2 bslmux_9_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01089 bsm_0_9_in_2 bslmux_12_com_2 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01088 bsm_0_15_out_2_s bslmux_11_com_2 bsm_0_9_in_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01087 bslmux_8_out_1 bslmux_12_com_2 bsm_0_15_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01086 bsoout_14_out_1_s bslmux_11_com_2 bslmux_8_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01085 bslmux_8_out_2 bslmux_12_com_2 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01084 bsoout_14_out_2_s bslmux_11_com_2 bslmux_8_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01083 bslmux_7_out_1 bslmux_12_com_2 bsoout_14_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01082 bsoout_13_out_1_s bslmux_11_com_2 bslmux_7_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01081 bslmux_7_out_2 bslmux_12_com_2 bsoout_13_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01080 bsoout_13_out_2_s bslmux_11_com_2 bslmux_7_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01079 bslmux_6_out_1 bslmux_12_com_2 bsoout_13_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01078 bsoout_12_out_1_s bslmux_11_com_2 bslmux_6_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01077 bslmux_6_out_2 bslmux_12_com_2 bsoout_12_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01076 bsm_0_12_out_2_s bslmux_11_com_2 bslmux_6_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01075 bslmux_5_out_1 bslmux_12_com_2 bsm_0_12_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01074 bsoout_11_out_1_s bslmux_11_com_2 bslmux_5_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01073 bslmux_5_out_2 bslmux_12_com_2 bsoout_11_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01072 bsm_0_11_out_2_s bslmux_11_com_2 bslmux_5_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01071 bslmux_4_out_1 bslmux_12_com_2 bsm_0_11_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01070 bsoout_10_out_1_s bslmux_11_com_2 bslmux_4_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01069 bslmux_4_out_2 bslmux_12_com_2 bsoout_10_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01068 bsm_0_10_out_2_s bslmux_11_com_2 bslmux_4_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01067 bslmux_3_out_1 bslmux_12_com_2 bsm_0_10_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01066 bsoout_9_out_1_s bslmux_11_com_2 bslmux_3_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01065 bslmux_3_out_2 bslmux_12_com_2 bsoout_9_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01064 bsm_0_9_out_2_s bslmux_11_com_2 bslmux_3_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01063 bslmux_2_out_1 bslmux_12_com_2 bsm_0_9_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01062 bsoout_8_out_1_s bslmux_11_com_2 bslmux_2_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01061 bslmux_2_out_2 bslmux_12_com_2 bsoout_8_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01060 bsoout_8_out_2_s bslmux_11_com_2 bslmux_2_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01059 bslmux_1_out_1 bslmux_12_com_2 bsoout_8_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01058 bsoout_7_out_1_s bslmux_11_com_2 bslmux_1_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01057 bslmux_1_out_2 bslmux_12_com_2 bsoout_7_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01056 bsm_0_7_out_2_s bslmux_11_com_2 bslmux_1_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01055 bslmux_0_out_1 bslmux_12_com_2 bsm_0_7_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01054 bsoout_6_out_1_s bslmux_11_com_2 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01053 bslmux_0_out_2 bslmux_12_com_2 bsoout_6_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01052 bsm_0_6_out_2_s bslmux_11_com_2 bslmux_0_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01051 bsrmux_15_f1 bslmux_12_com_2 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01050 bsoout_5_out_1_s bslmux_11_com_2 bsrmux_15_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01049 n681 bslmux_12_com_2 bsoout_5_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01048 bsm_0_5_out_2_s bslmux_11_com_2 n681 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01047 bsrmux_14_f1 bslmux_12_com_2 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01046 bsoout_4_out_1_s bslmux_11_com_2 bsrmux_14_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01045 n676 bslmux_12_com_2 bsoout_4_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01044 bsm_0_4_out_2_s bslmux_11_com_2 n676 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01043 bsrmux_13_f1 bslmux_12_com_2 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01042 bsoout_3_out_1_s bslmux_11_com_2 bsrmux_13_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01041 n673 bslmux_12_com_2 bsoout_3_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01040 bsoout_3_out_2_s bslmux_11_com_2 n673 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01039 bsrmux_12_f1 bslmux_12_com_2 bsoout_3_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01038 bsoout_2_out_1_s bslmux_11_com_2 bsrmux_12_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01037 n671 bslmux_12_com_2 bsoout_2_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01036 bsm_0_2_out_2_s bslmux_11_com_2 n671 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01035 bsrmux_11_f1 bslmux_12_com_2 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01034 bsoout_1_out_1_s bslmux_11_com_2 bsrmux_11_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01033 n666 bslmux_12_com_2 bsoout_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01032 bsm_0_1_out_2_s bslmux_11_com_2 n666 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01031 bsrmux_10_f1 bslmux_12_com_2 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01030 bsoout_0_out_1_s bslmux_11_com_2 bsrmux_10_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01029 n662 bslmux_12_com_2 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01028 bsm_0_0_out_2_s bslmux_11_com_2 n662 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01027 bsrmux_9_f1 bslmux_12_com_2 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01026 bsoout_15_out_1_s bslmux_9_com_2 bslmux_10_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01025 bsm_0_10_in_2 bslmux_10_com_2 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01024 bsm_0_15_out_2_s bslmux_9_com_2 bsm_0_10_in_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01023 bslmux_9_out_1 bslmux_10_com_2 bsm_0_15_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01022 bsoout_14_out_1_s bslmux_9_com_2 bslmux_9_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01021 bsm_0_9_in_2 bslmux_10_com_2 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01020 bsoout_14_out_2_s bslmux_9_com_2 bsm_0_9_in_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01019 bslmux_8_out_1 bslmux_10_com_2 bsoout_14_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01018 bsoout_13_out_1_s bslmux_9_com_2 bslmux_8_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01017 bslmux_8_out_2 bslmux_10_com_2 bsoout_13_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01016 bsoout_13_out_2_s bslmux_9_com_2 bslmux_8_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01015 bslmux_7_out_1 bslmux_10_com_2 bsoout_13_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01014 bsoout_12_out_1_s bslmux_9_com_2 bslmux_7_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01013 bslmux_7_out_2 bslmux_10_com_2 bsoout_12_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01012 bsm_0_12_out_2_s bslmux_9_com_2 bslmux_7_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01011 bslmux_6_out_1 bslmux_10_com_2 bsm_0_12_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01010 bsoout_11_out_1_s bslmux_9_com_2 bslmux_6_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01009 bslmux_6_out_2 bslmux_10_com_2 bsoout_11_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01008 bsm_0_11_out_2_s bslmux_9_com_2 bslmux_6_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01007 bslmux_5_out_1 bslmux_10_com_2 bsm_0_11_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01006 bsoout_10_out_1_s bslmux_9_com_2 bslmux_5_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01005 bslmux_5_out_2 bslmux_10_com_2 bsoout_10_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01004 bsm_0_10_out_2_s bslmux_9_com_2 bslmux_5_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01003 bslmux_4_out_1 bslmux_10_com_2 bsm_0_10_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01002 bsoout_9_out_1_s bslmux_9_com_2 bslmux_4_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01001 bslmux_4_out_2 bslmux_10_com_2 bsoout_9_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01000 bsm_0_9_out_2_s bslmux_9_com_2 bslmux_4_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00999 bslmux_3_out_1 bslmux_10_com_2 bsm_0_9_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00998 bsoout_8_out_1_s bslmux_9_com_2 bslmux_3_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00997 bslmux_3_out_2 bslmux_10_com_2 bsoout_8_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00996 bsoout_8_out_2_s bslmux_9_com_2 bslmux_3_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00995 bslmux_2_out_1 bslmux_10_com_2 bsoout_8_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00994 bsoout_7_out_1_s bslmux_9_com_2 bslmux_2_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00993 bslmux_2_out_2 bslmux_10_com_2 bsoout_7_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00992 bsm_0_7_out_2_s bslmux_9_com_2 bslmux_2_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00991 bslmux_1_out_1 bslmux_10_com_2 bsm_0_7_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00990 bsoout_6_out_1_s bslmux_9_com_2 bslmux_1_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00989 bslmux_1_out_2 bslmux_10_com_2 bsoout_6_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00988 bsm_0_6_out_2_s bslmux_9_com_2 bslmux_1_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00987 bslmux_0_out_1 bslmux_10_com_2 bsm_0_6_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00986 bsoout_5_out_1_s bslmux_9_com_2 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00985 bslmux_0_out_2 bslmux_10_com_2 bsoout_5_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00984 bsm_0_5_out_2_s bslmux_9_com_2 bslmux_0_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00983 bsrmux_15_f1 bslmux_10_com_2 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00982 bsoout_4_out_1_s bslmux_9_com_2 bsrmux_15_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00981 n681 bslmux_10_com_2 bsoout_4_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00980 bsm_0_4_out_2_s bslmux_9_com_2 n681 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00979 bsrmux_14_f1 bslmux_10_com_2 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00978 bsoout_3_out_1_s bslmux_9_com_2 bsrmux_14_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00977 n676 bslmux_10_com_2 bsoout_3_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00976 bsoout_3_out_2_s bslmux_9_com_2 n676 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00975 bsrmux_13_f1 bslmux_10_com_2 bsoout_3_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00974 bsoout_2_out_1_s bslmux_9_com_2 bsrmux_13_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00973 n673 bslmux_10_com_2 bsoout_2_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00972 bsm_0_2_out_2_s bslmux_9_com_2 n673 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00971 bsrmux_12_f1 bslmux_10_com_2 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00970 bsoout_1_out_1_s bslmux_9_com_2 bsrmux_12_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00969 n671 bslmux_10_com_2 bsoout_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00968 bsm_0_1_out_2_s bslmux_9_com_2 n671 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00967 bsrmux_11_f1 bslmux_10_com_2 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00966 bsoout_0_out_1_s bslmux_9_com_2 bsrmux_11_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00965 n666 bslmux_10_com_2 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00964 bsm_0_0_out_2_s bslmux_9_com_2 n666 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00963 bsrmux_10_f1 bslmux_10_com_2 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00962 bsoout_15_out_1_s bslmux_7_com_2 bslmux_11_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00961 bslmux_11_out_2 bslmux_8_com_2 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00960 bsm_0_15_out_2_s bslmux_7_com_2 bslmux_11_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00959 bslmux_10_out_1 bslmux_8_com_2 bsm_0_15_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00958 bsoout_14_out_1_s bslmux_7_com_2 bslmux_10_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00957 bsm_0_10_in_2 bslmux_8_com_2 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00956 bsoout_14_out_2_s bslmux_7_com_2 bsm_0_10_in_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00955 bslmux_9_out_1 bslmux_8_com_2 bsoout_14_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00954 bsoout_13_out_1_s bslmux_7_com_2 bslmux_9_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00953 bsm_0_9_in_2 bslmux_8_com_2 bsoout_13_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00952 bsoout_13_out_2_s bslmux_7_com_2 bsm_0_9_in_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00951 bslmux_8_out_1 bslmux_8_com_2 bsoout_13_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00950 bsoout_12_out_1_s bslmux_7_com_2 bslmux_8_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00949 bslmux_8_out_2 bslmux_8_com_2 bsoout_12_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00948 bsm_0_12_out_2_s bslmux_7_com_2 bslmux_8_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00947 bslmux_7_out_1 bslmux_8_com_2 bsm_0_12_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00946 bsoout_11_out_1_s bslmux_7_com_2 bslmux_7_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00945 bslmux_7_out_2 bslmux_8_com_2 bsoout_11_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00944 bsm_0_11_out_2_s bslmux_7_com_2 bslmux_7_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00943 bslmux_6_out_1 bslmux_8_com_2 bsm_0_11_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00942 bsoout_10_out_1_s bslmux_7_com_2 bslmux_6_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00941 bslmux_6_out_2 bslmux_8_com_2 bsoout_10_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00940 bsm_0_10_out_2_s bslmux_7_com_2 bslmux_6_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00939 bslmux_5_out_1 bslmux_8_com_2 bsm_0_10_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00938 bsoout_9_out_1_s bslmux_7_com_2 bslmux_5_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00937 bslmux_5_out_2 bslmux_8_com_2 bsoout_9_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00936 bsm_0_9_out_2_s bslmux_7_com_2 bslmux_5_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00935 bslmux_4_out_1 bslmux_8_com_2 bsm_0_9_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00934 bsoout_8_out_1_s bslmux_7_com_2 bslmux_4_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00933 bslmux_4_out_2 bslmux_8_com_2 bsoout_8_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00932 bsoout_8_out_2_s bslmux_7_com_2 bslmux_4_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00931 bslmux_3_out_1 bslmux_8_com_2 bsoout_8_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00930 bsoout_7_out_1_s bslmux_7_com_2 bslmux_3_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00929 bslmux_3_out_2 bslmux_8_com_2 bsoout_7_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00928 bsm_0_7_out_2_s bslmux_7_com_2 bslmux_3_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00927 bslmux_2_out_1 bslmux_8_com_2 bsm_0_7_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00926 bsoout_6_out_1_s bslmux_7_com_2 bslmux_2_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00925 bslmux_2_out_2 bslmux_8_com_2 bsoout_6_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00924 bsm_0_6_out_2_s bslmux_7_com_2 bslmux_2_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00923 bslmux_1_out_1 bslmux_8_com_2 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00922 bsoout_5_out_1_s bslmux_7_com_2 bslmux_1_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00921 bslmux_1_out_2 bslmux_8_com_2 bsoout_5_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00920 bsm_0_5_out_2_s bslmux_7_com_2 bslmux_1_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00919 bslmux_0_out_1 bslmux_8_com_2 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00918 bsoout_4_out_1_s bslmux_7_com_2 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00917 bslmux_0_out_2 bslmux_8_com_2 bsoout_4_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00916 bsm_0_4_out_2_s bslmux_7_com_2 bslmux_0_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00915 bsrmux_15_f1 bslmux_8_com_2 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00914 bsoout_3_out_1_s bslmux_7_com_2 bsrmux_15_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00913 n681 bslmux_8_com_2 bsoout_3_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00912 bsoout_3_out_2_s bslmux_7_com_2 n681 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00911 bsrmux_14_f1 bslmux_8_com_2 bsoout_3_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00910 bsoout_2_out_1_s bslmux_7_com_2 bsrmux_14_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00909 n676 bslmux_8_com_2 bsoout_2_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00908 bsm_0_2_out_2_s bslmux_7_com_2 n676 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00907 bsrmux_13_f1 bslmux_8_com_2 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00906 bsoout_1_out_1_s bslmux_7_com_2 bsrmux_13_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00905 n673 bslmux_8_com_2 bsoout_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00904 bsm_0_1_out_2_s bslmux_7_com_2 n673 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00903 bsrmux_12_f1 bslmux_8_com_2 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00902 bsoout_0_out_1_s bslmux_7_com_2 bsrmux_12_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00901 n671 bslmux_8_com_2 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00900 bsm_0_0_out_2_s bslmux_7_com_2 n671 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00899 bsrmux_11_f1 bslmux_8_com_2 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00898 bsoout_15_out_1_s bslmux_5_com_2 bslmux_12_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00897 bslmux_12_out_2 bslmux_6_com_2 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00896 bsm_0_15_out_2_s bslmux_5_com_2 bslmux_12_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00895 bslmux_11_out_1 bslmux_6_com_2 bsm_0_15_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00894 bsoout_14_out_1_s bslmux_5_com_2 bslmux_11_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00893 bslmux_11_out_2 bslmux_6_com_2 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00892 bsoout_14_out_2_s bslmux_5_com_2 bslmux_11_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00891 bslmux_10_out_1 bslmux_6_com_2 bsoout_14_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00890 bsoout_13_out_1_s bslmux_5_com_2 bslmux_10_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00889 bsm_0_10_in_2 bslmux_6_com_2 bsoout_13_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00888 bsoout_13_out_2_s bslmux_5_com_2 bsm_0_10_in_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00887 bslmux_9_out_1 bslmux_6_com_2 bsoout_13_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00886 bsoout_12_out_1_s bslmux_5_com_2 bslmux_9_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00885 bsm_0_9_in_2 bslmux_6_com_2 bsoout_12_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00884 bsm_0_12_out_2_s bslmux_5_com_2 bsm_0_9_in_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00883 bslmux_8_out_1 bslmux_6_com_2 bsm_0_12_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00882 bsoout_11_out_1_s bslmux_5_com_2 bslmux_8_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00881 bslmux_8_out_2 bslmux_6_com_2 bsoout_11_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00880 bsm_0_11_out_2_s bslmux_5_com_2 bslmux_8_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00879 bslmux_7_out_1 bslmux_6_com_2 bsm_0_11_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00878 bsoout_10_out_1_s bslmux_5_com_2 bslmux_7_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00877 bslmux_7_out_2 bslmux_6_com_2 bsoout_10_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00876 bsm_0_10_out_2_s bslmux_5_com_2 bslmux_7_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00875 bslmux_6_out_1 bslmux_6_com_2 bsm_0_10_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00874 bsoout_9_out_1_s bslmux_5_com_2 bslmux_6_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00873 bslmux_6_out_2 bslmux_6_com_2 bsoout_9_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00872 bsm_0_9_out_2_s bslmux_5_com_2 bslmux_6_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00871 bslmux_5_out_1 bslmux_6_com_2 bsm_0_9_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00870 bsoout_8_out_1_s bslmux_5_com_2 bslmux_5_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00869 bslmux_5_out_2 bslmux_6_com_2 bsoout_8_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00868 bsoout_8_out_2_s bslmux_5_com_2 bslmux_5_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00867 bslmux_4_out_1 bslmux_6_com_2 bsoout_8_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00866 bsoout_7_out_1_s bslmux_5_com_2 bslmux_4_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00865 bslmux_4_out_2 bslmux_6_com_2 bsoout_7_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00864 bsm_0_7_out_2_s bslmux_5_com_2 bslmux_4_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00863 bslmux_3_out_1 bslmux_6_com_2 bsm_0_7_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00862 bsoout_6_out_1_s bslmux_5_com_2 bslmux_3_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00861 bslmux_3_out_2 bslmux_6_com_2 bsoout_6_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00860 bsm_0_6_out_2_s bslmux_5_com_2 bslmux_3_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00859 bslmux_2_out_1 bslmux_6_com_2 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00858 bsoout_5_out_1_s bslmux_5_com_2 bslmux_2_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00857 bslmux_2_out_2 bslmux_6_com_2 bsoout_5_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00856 bsm_0_5_out_2_s bslmux_5_com_2 bslmux_2_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00855 bslmux_1_out_1 bslmux_6_com_2 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00854 bsoout_4_out_1_s bslmux_5_com_2 bslmux_1_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00853 bslmux_1_out_2 bslmux_6_com_2 bsoout_4_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00852 bsm_0_4_out_2_s bslmux_5_com_2 bslmux_1_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00851 bslmux_0_out_1 bslmux_6_com_2 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00850 bsoout_3_out_1_s bslmux_5_com_2 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00849 bslmux_0_out_2 bslmux_6_com_2 bsoout_3_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00848 bsoout_3_out_2_s bslmux_5_com_2 bslmux_0_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00847 bsrmux_15_f1 bslmux_6_com_2 bsoout_3_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00846 bsoout_2_out_1_s bslmux_5_com_2 bsrmux_15_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00845 n681 bslmux_6_com_2 bsoout_2_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00844 bsm_0_2_out_2_s bslmux_5_com_2 n681 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00843 bsrmux_14_f1 bslmux_6_com_2 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00842 bsoout_1_out_1_s bslmux_5_com_2 bsrmux_14_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00841 n676 bslmux_6_com_2 bsoout_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00840 bsm_0_1_out_2_s bslmux_5_com_2 n676 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00839 bsrmux_13_f1 bslmux_6_com_2 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00838 bsoout_0_out_1_s bslmux_5_com_2 bsrmux_13_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00837 n673 bslmux_6_com_2 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00836 bsm_0_0_out_2_s bslmux_5_com_2 n673 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00835 bsrmux_12_f1 bslmux_6_com_2 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00834 bsoout_15_out_1_s bslmux_3_com_2 bslmux_13_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00833 bslmux_13_out_2 bslmux_4_com_2 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00832 bsm_0_15_out_2_s bslmux_3_com_2 bslmux_13_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00831 bslmux_12_out_1 bslmux_4_com_2 bsm_0_15_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00830 bsoout_14_out_1_s bslmux_3_com_2 bslmux_12_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00829 bslmux_12_out_2 bslmux_4_com_2 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00828 bsoout_14_out_2_s bslmux_3_com_2 bslmux_12_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00827 bslmux_11_out_1 bslmux_4_com_2 bsoout_14_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00826 bsoout_13_out_1_s bslmux_3_com_2 bslmux_11_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00825 bslmux_11_out_2 bslmux_4_com_2 bsoout_13_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00824 bsoout_13_out_2_s bslmux_3_com_2 bslmux_11_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00823 bslmux_10_out_1 bslmux_4_com_2 bsoout_13_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00822 bsoout_12_out_1_s bslmux_3_com_2 bslmux_10_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00821 bsm_0_10_in_2 bslmux_4_com_2 bsoout_12_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00820 bsm_0_12_out_2_s bslmux_3_com_2 bsm_0_10_in_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00819 bslmux_9_out_1 bslmux_4_com_2 bsm_0_12_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00818 bsoout_11_out_1_s bslmux_3_com_2 bslmux_9_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00817 bsm_0_9_in_2 bslmux_4_com_2 bsoout_11_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00816 bsm_0_11_out_2_s bslmux_3_com_2 bsm_0_9_in_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00815 bslmux_8_out_1 bslmux_4_com_2 bsm_0_11_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00814 bsoout_10_out_1_s bslmux_3_com_2 bslmux_8_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00813 bslmux_8_out_2 bslmux_4_com_2 bsoout_10_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00812 bsm_0_10_out_2_s bslmux_3_com_2 bslmux_8_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00811 bslmux_7_out_1 bslmux_4_com_2 bsm_0_10_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00810 bsoout_9_out_1_s bslmux_3_com_2 bslmux_7_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00809 bslmux_7_out_2 bslmux_4_com_2 bsoout_9_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00808 bsm_0_9_out_2_s bslmux_3_com_2 bslmux_7_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00807 bslmux_6_out_1 bslmux_4_com_2 bsm_0_9_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00806 bsoout_8_out_1_s bslmux_3_com_2 bslmux_6_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00805 bslmux_6_out_2 bslmux_4_com_2 bsoout_8_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00804 bsoout_8_out_2_s bslmux_3_com_2 bslmux_6_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00803 bslmux_5_out_1 bslmux_4_com_2 bsoout_8_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00802 bsoout_7_out_1_s bslmux_3_com_2 bslmux_5_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00801 bslmux_5_out_2 bslmux_4_com_2 bsoout_7_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00800 bsm_0_7_out_2_s bslmux_3_com_2 bslmux_5_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00799 bslmux_4_out_1 bslmux_4_com_2 bsm_0_7_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00798 bsoout_6_out_1_s bslmux_3_com_2 bslmux_4_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00797 bslmux_4_out_2 bslmux_4_com_2 bsoout_6_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00796 bsm_0_6_out_2_s bslmux_3_com_2 bslmux_4_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00795 bslmux_3_out_1 bslmux_4_com_2 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00794 bsoout_5_out_1_s bslmux_3_com_2 bslmux_3_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00793 bslmux_3_out_2 bslmux_4_com_2 bsoout_5_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00792 bsm_0_5_out_2_s bslmux_3_com_2 bslmux_3_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00791 bslmux_2_out_1 bslmux_4_com_2 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00790 bsoout_4_out_1_s bslmux_3_com_2 bslmux_2_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00789 bslmux_2_out_2 bslmux_4_com_2 bsoout_4_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00788 bsm_0_4_out_2_s bslmux_3_com_2 bslmux_2_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00787 bslmux_1_out_1 bslmux_4_com_2 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00786 bsoout_3_out_1_s bslmux_3_com_2 bslmux_1_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00785 bslmux_1_out_2 bslmux_4_com_2 bsoout_3_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00784 bsoout_3_out_2_s bslmux_3_com_2 bslmux_1_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00783 bslmux_0_out_1 bslmux_4_com_2 bsoout_3_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00782 bsoout_2_out_1_s bslmux_3_com_2 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00781 bslmux_0_out_2 bslmux_4_com_2 bsoout_2_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00780 bsm_0_2_out_2_s bslmux_3_com_2 bslmux_0_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00779 bsrmux_15_f1 bslmux_4_com_2 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00778 bsoout_1_out_1_s bslmux_3_com_2 bsrmux_15_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00777 n681 bslmux_4_com_2 bsoout_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00776 bsm_0_1_out_2_s bslmux_3_com_2 n681 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00775 bsrmux_14_f1 bslmux_4_com_2 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00774 bsoout_0_out_1_s bslmux_3_com_2 bsrmux_14_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00773 n676 bslmux_4_com_2 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00772 bsm_0_0_out_2_s bslmux_3_com_2 n676 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00771 bsrmux_13_f1 bslmux_4_com_2 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00770 bsoout_15_out_1_s bslmux_1_com_2 bslmux_14_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00769 bslmux_14_out_2 bslmux_2_com_2 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00768 bsm_0_15_out_2_s bslmux_1_com_2 bslmux_14_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00767 bslmux_13_out_1 bslmux_2_com_2 bsm_0_15_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00766 bsoout_14_out_1_s bslmux_1_com_2 bslmux_13_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00765 bslmux_13_out_2 bslmux_2_com_2 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00764 bsoout_14_out_2_s bslmux_1_com_2 bslmux_13_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00763 bslmux_12_out_1 bslmux_2_com_2 bsoout_14_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00762 bsoout_13_out_1_s bslmux_1_com_2 bslmux_12_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00761 bslmux_12_out_2 bslmux_2_com_2 bsoout_13_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00760 bsoout_13_out_2_s bslmux_1_com_2 bslmux_12_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00759 bslmux_11_out_1 bslmux_2_com_2 bsoout_13_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00758 bsoout_12_out_1_s bslmux_1_com_2 bslmux_11_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00757 bslmux_11_out_2 bslmux_2_com_2 bsoout_12_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00756 bsm_0_12_out_2_s bslmux_1_com_2 bslmux_11_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00755 bslmux_10_out_1 bslmux_2_com_2 bsm_0_12_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00754 bsoout_11_out_1_s bslmux_1_com_2 bslmux_10_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00753 bsm_0_10_in_2 bslmux_2_com_2 bsoout_11_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00752 bsm_0_11_out_2_s bslmux_1_com_2 bsm_0_10_in_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00751 bslmux_9_out_1 bslmux_2_com_2 bsm_0_11_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00750 bsoout_10_out_1_s bslmux_1_com_2 bslmux_9_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00749 bsm_0_9_in_2 bslmux_2_com_2 bsoout_10_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00748 bsm_0_10_out_2_s bslmux_1_com_2 bsm_0_9_in_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00747 bslmux_8_out_1 bslmux_2_com_2 bsm_0_10_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00746 bsoout_9_out_1_s bslmux_1_com_2 bslmux_8_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00745 bslmux_8_out_2 bslmux_2_com_2 bsoout_9_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00744 bsm_0_9_out_2_s bslmux_1_com_2 bslmux_8_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00743 bslmux_7_out_1 bslmux_2_com_2 bsm_0_9_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00742 bsoout_8_out_1_s bslmux_1_com_2 bslmux_7_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00741 bslmux_7_out_2 bslmux_2_com_2 bsoout_8_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00740 bsoout_8_out_2_s bslmux_1_com_2 bslmux_7_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00739 bslmux_6_out_1 bslmux_2_com_2 bsoout_8_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00738 bsoout_7_out_1_s bslmux_1_com_2 bslmux_6_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00737 bslmux_6_out_2 bslmux_2_com_2 bsoout_7_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00736 bsm_0_7_out_2_s bslmux_1_com_2 bslmux_6_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00735 bslmux_5_out_1 bslmux_2_com_2 bsm_0_7_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00734 bsoout_6_out_1_s bslmux_1_com_2 bslmux_5_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00733 bslmux_5_out_2 bslmux_2_com_2 bsoout_6_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00732 bsm_0_6_out_2_s bslmux_1_com_2 bslmux_5_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00731 bslmux_4_out_1 bslmux_2_com_2 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00730 bsoout_5_out_1_s bslmux_1_com_2 bslmux_4_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00729 bslmux_4_out_2 bslmux_2_com_2 bsoout_5_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00728 bsm_0_5_out_2_s bslmux_1_com_2 bslmux_4_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00727 bslmux_3_out_1 bslmux_2_com_2 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00726 bsoout_4_out_1_s bslmux_1_com_2 bslmux_3_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00725 bslmux_3_out_2 bslmux_2_com_2 bsoout_4_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00724 bsm_0_4_out_2_s bslmux_1_com_2 bslmux_3_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00723 bslmux_2_out_1 bslmux_2_com_2 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00722 bsoout_3_out_1_s bslmux_1_com_2 bslmux_2_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00721 bslmux_2_out_2 bslmux_2_com_2 bsoout_3_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00720 bsoout_3_out_2_s bslmux_1_com_2 bslmux_2_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00719 bslmux_1_out_1 bslmux_2_com_2 bsoout_3_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00718 bsoout_2_out_1_s bslmux_1_com_2 bslmux_1_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00717 bslmux_1_out_2 bslmux_2_com_2 bsoout_2_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00716 bsm_0_2_out_2_s bslmux_1_com_2 bslmux_1_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00715 bslmux_0_out_1 bslmux_2_com_2 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00714 bsoout_1_out_1_s bslmux_1_com_2 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00713 bslmux_0_out_2 bslmux_2_com_2 bsoout_1_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00712 bsm_0_1_out_2_s bslmux_1_com_2 bslmux_0_out_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00711 bsrmux_15_f1 bslmux_2_com_2 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00710 bsoout_0_out_1_s bslmux_1_com_2 bsrmux_15_f1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00709 n681 bslmux_2_com_2 bsoout_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00708 bsm_0_0_out_2_s bslmux_1_com_2 n681 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00707 bsrmux_14_f1 bslmux_2_com_2 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00706 bsoout_15_out_1_s bssnbl_15_out_1 bslmux_15_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00705 bsm_0_15_in_2 bssnbl_0_out_2 bsoout_15_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00704 bsm_0_15_out_2_s bssnbl_15_out_1 bsm_0_15_in_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00703 bslmux_14_out_1 bssnbl_0_out_2 bsm_0_15_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00702 bsoout_14_out_1_s bssnbl_15_out_1 bslmux_14_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00701 bslmux_14_out_2 bssnbl_0_out_2 bsoout_14_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00700 bsoout_14_out_2_s bssnbl_15_out_1 bslmux_14_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00699 bslmux_13_out_1 bssnbl_0_out_2 bsoout_14_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00698 bsoout_13_out_1_s bssnbl_15_out_1 bslmux_13_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00697 bslmux_13_out_2 bssnbl_0_out_2 bsoout_13_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00696 bsoout_13_out_2_s bssnbl_15_out_1 bslmux_13_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00695 bslmux_12_out_1 bssnbl_0_out_2 bsoout_13_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00694 bsoout_12_out_1_s bssnbl_15_out_1 bslmux_12_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00693 bslmux_12_out_2 bssnbl_0_out_2 bsoout_12_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00692 bsm_0_12_out_2_s bssnbl_15_out_1 bslmux_12_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00691 bslmux_11_out_1 bssnbl_0_out_2 bsm_0_12_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00690 bsoout_11_out_1_s bssnbl_15_out_1 bslmux_11_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00689 bslmux_11_out_2 bssnbl_0_out_2 bsoout_11_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00688 bsm_0_11_out_2_s bssnbl_15_out_1 bslmux_11_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00687 bslmux_10_out_1 bssnbl_0_out_2 bsm_0_11_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00686 bsoout_10_out_1_s bssnbl_15_out_1 bslmux_10_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00685 bsm_0_10_in_2 bssnbl_0_out_2 bsoout_10_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00684 bsm_0_10_out_2_s bssnbl_15_out_1 bsm_0_10_in_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00683 bslmux_9_out_1 bssnbl_0_out_2 bsm_0_10_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00682 bsoout_9_out_1_s bssnbl_15_out_1 bslmux_9_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00681 bsm_0_9_in_2 bssnbl_0_out_2 bsoout_9_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00680 bsm_0_9_out_2_s bssnbl_15_out_1 bsm_0_9_in_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00679 bslmux_8_out_1 bssnbl_0_out_2 bsm_0_9_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00678 bsoout_8_out_1_s bssnbl_15_out_1 bslmux_8_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00677 bslmux_8_out_2 bssnbl_0_out_2 bsoout_8_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00676 bsoout_8_out_2_s bssnbl_15_out_1 bslmux_8_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00675 bslmux_7_out_1 bssnbl_0_out_2 bsoout_8_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00674 bsoout_7_out_1_s bssnbl_15_out_1 bslmux_7_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00673 bslmux_7_out_2 bssnbl_0_out_2 bsoout_7_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00672 bsm_0_7_out_2_s bssnbl_15_out_1 bslmux_7_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00671 bslmux_6_out_1 bssnbl_0_out_2 bsm_0_7_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00670 bsoout_6_out_1_s bssnbl_15_out_1 bslmux_6_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00669 bslmux_6_out_2 bssnbl_0_out_2 bsoout_6_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00668 bsm_0_6_out_2_s bssnbl_15_out_1 bslmux_6_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00667 bslmux_5_out_1 bssnbl_0_out_2 bsm_0_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00666 bsoout_5_out_1_s bssnbl_15_out_1 bslmux_5_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00665 bslmux_5_out_2 bssnbl_0_out_2 bsoout_5_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00664 bsm_0_5_out_2_s bssnbl_15_out_1 bslmux_5_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00663 bslmux_4_out_1 bssnbl_0_out_2 bsm_0_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00662 bsoout_4_out_1_s bssnbl_15_out_1 bslmux_4_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00661 bslmux_4_out_2 bssnbl_0_out_2 bsoout_4_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00660 bsm_0_4_out_2_s bssnbl_15_out_1 bslmux_4_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00659 bslmux_3_out_1 bssnbl_0_out_2 bsm_0_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00658 bsoout_3_out_1_s bssnbl_15_out_1 bslmux_3_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00657 bslmux_3_out_2 bssnbl_0_out_2 bsoout_3_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00656 bsoout_3_out_2_s bssnbl_15_out_1 bslmux_3_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00655 bslmux_2_out_1 bssnbl_0_out_2 bsoout_3_out_2_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00654 bsoout_2_out_1_s bssnbl_15_out_1 bslmux_2_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00653 bslmux_2_out_2 bssnbl_0_out_2 bsoout_2_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00652 bsm_0_2_out_2_s bssnbl_15_out_1 bslmux_2_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00651 bslmux_1_out_1 bssnbl_0_out_2 bsm_0_2_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00650 bsoout_1_out_1_s bssnbl_15_out_1 bslmux_1_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00649 bslmux_1_out_2 bssnbl_0_out_2 bsoout_1_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00648 bsm_0_1_out_2_s bssnbl_15_out_1 bslmux_1_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00647 bslmux_0_out_1 bssnbl_0_out_2 bsm_0_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00646 bsoout_0_out_1_s bssnbl_15_out_1 bslmux_0_out_1 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00645 bslmux_0_out_2 bssnbl_0_out_2 bsoout_0_out_1_s vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00644 bsm_0_0_out_2_s bssnbl_15_out_1 bslmux_0_out_2 vss TN L=0.18U 
+ W=1.26U AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00643 bsrmux_15_f1 bssnbl_0_out_2 bsm_0_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00642 n19 in_d_31 n31 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00641 bsm_0_15_in_2 n41 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00640 vss n41 bsm_0_15_in_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00639 bsm_0_15_in_2 n41 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00638 vss n43 n42 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00637 n42 bshlmx_0_asr n41 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00636 vss bshlmx_0_lsl n44 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00635 n44 in_d_30 n43 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00634 bslmux_15_out_1 n30 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00633 vss n30 bslmux_15_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00632 bslmux_15_out_1 n30 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00631 vss n31 n18 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00630 n18 bshlmx_0_asr n30 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00629 vss bshlmx_0_lsl n19 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00628 n58 in_d_29 n68 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00627 bslmux_14_out_2 n80 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00626 vss n80 bslmux_14_out_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00625 bslmux_14_out_2 n80 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00624 vss n84 n81 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00623 n81 bshlmx_0_asr n80 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00622 vss bshlmx_0_lsl n82 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00621 n82 in_d_28 n84 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00620 bslmux_14_out_1 n69 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00619 vss n69 bslmux_14_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00618 bslmux_14_out_1 n69 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00617 vss n68 n57 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00616 n57 bshlmx_0_asr n69 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00615 vss bshlmx_0_lsl n58 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00614 n83 in_d_27 n97 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00613 bslmux_13_out_2 n116 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00612 vss n116 bslmux_13_out_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00611 bslmux_13_out_2 n116 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00610 vss n118 n117 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00609 n117 bshlmx_0_asr n116 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00608 vss bshlmx_0_lsl n119 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00607 n119 in_d_26 n118 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00606 bslmux_13_out_1 n106 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00605 vss n106 bslmux_13_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00604 bslmux_13_out_1 n106 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00603 vss n97 n96 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00602 n96 bshlmx_0_asr n106 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00601 vss bshlmx_0_lsl n83 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00600 n124 in_d_25 n140 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00599 bslmux_12_out_2 n156 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00598 vss n156 bslmux_12_out_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00597 bslmux_12_out_2 n156 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00596 vss n158 n157 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00595 n157 bshlmx_0_asr n156 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00594 vss bshlmx_0_lsl n159 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00593 n159 in_d_24 n158 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00592 bslmux_12_out_1 n146 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00591 vss n146 bslmux_12_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00590 bslmux_12_out_1 n146 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00589 vss n140 n139 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00588 n139 bshlmx_0_asr n146 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00587 vss bshlmx_0_lsl n124 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00586 n171 in_d_23 n183 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00585 bslmux_11_out_2 n194 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00584 vss n194 bslmux_11_out_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00583 bslmux_11_out_2 n194 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00582 vss n196 n195 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00581 n195 bshlmx_0_asr n194 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00580 vss bshlmx_0_lsl n197 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00579 n197 in_d_22 n196 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00578 bslmux_11_out_1 n182 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00577 vss n182 bslmux_11_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00576 bslmux_11_out_1 n182 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00575 vss n183 n170 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00574 n170 bshlmx_0_asr n182 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00573 vss bshlmx_0_lsl n171 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00572 n210 in_d_21 n221 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00571 bsm_0_10_in_2 n232 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00570 vss n232 bsm_0_10_in_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00569 bsm_0_10_in_2 n232 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00568 vss n234 n233 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00567 n233 bshlmx_0_asr n232 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00566 vss bshlmx_0_lsl n235 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00565 n235 in_d_20 n234 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00564 bslmux_10_out_1 n220 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00563 vss n220 bslmux_10_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00562 bslmux_10_out_1 n220 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00561 vss n221 n209 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00560 n209 bshlmx_0_asr n220 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00559 vss bshlmx_0_lsl n210 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00558 n248 in_d_19 n258 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00557 bsm_0_9_in_2 n270 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00556 vss n270 bsm_0_9_in_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00555 bsm_0_9_in_2 n270 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00554 vss n273 n271 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00553 n271 bshlmx_0_asr n270 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00552 vss bshlmx_0_lsl n274 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00551 n274 in_d_18 n273 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00550 bslmux_9_out_1 n259 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00549 vss n259 bslmux_9_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00548 bslmux_9_out_1 n259 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00547 vss n258 n247 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00546 n247 bshlmx_0_asr n259 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00545 vss bshlmx_0_lsl n248 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00544 n272 in_d_17 n297 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00543 bslmux_8_out_2 n306 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00542 vss n306 bslmux_8_out_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00541 bslmux_8_out_2 n306 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00540 vss n309 n307 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00539 n307 bshlmx_0_asr n306 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00538 vss bshlmx_0_lsl n308 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00537 n308 in_d_16 n309 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00536 bslmux_8_out_1 n295 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00535 vss n295 bslmux_8_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00534 bslmux_8_out_1 n295 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00533 vss n297 n286 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00532 n286 bshlmx_0_asr n295 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00531 vss bshlmx_0_lsl n272 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00530 n314 in_d_15 n325 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00529 bslmux_7_out_2 n346 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00528 vss n346 bslmux_7_out_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00527 bslmux_7_out_2 n346 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00526 vss n348 n347 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00525 n347 bshlmx_0_asr n346 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00524 vss bshlmx_0_lsl n349 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00523 n349 in_d_14 n348 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00522 bslmux_7_out_1 n335 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00521 vss n335 bslmux_7_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00520 bslmux_7_out_1 n335 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00519 vss n325 n324 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00518 n324 bshlmx_0_asr n335 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00517 vss bshlmx_0_lsl n314 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00516 n361 in_d_13 n373 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00515 bslmux_6_out_2 n384 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00514 vss n384 bslmux_6_out_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00513 bslmux_6_out_2 n384 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00512 vss n386 n385 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00511 n385 bshlmx_0_asr n384 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00510 vss bshlmx_0_lsl n387 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00509 n387 in_d_12 n386 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00508 bslmux_6_out_1 n372 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00507 vss n372 bslmux_6_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00506 bslmux_6_out_1 n372 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00505 vss n373 n360 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00504 n360 bshlmx_0_asr n372 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00503 vss bshlmx_0_lsl n361 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00502 n400 in_d_11 n411 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00501 bslmux_5_out_2 n422 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00500 vss n422 bslmux_5_out_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00499 bslmux_5_out_2 n422 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00498 vss n424 n423 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00497 n423 bshlmx_0_asr n422 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00496 vss bshlmx_0_lsl n425 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00495 n425 in_d_10 n424 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00494 bslmux_5_out_1 n410 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00493 vss n410 bslmux_5_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00492 bslmux_5_out_1 n410 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00491 vss n411 n399 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00490 n399 bshlmx_0_asr n410 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00489 vss bshlmx_0_lsl n400 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00488 n438 in_d_9 n450 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00487 bslmux_4_out_2 n460 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00486 vss n460 bslmux_4_out_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00485 bslmux_4_out_2 n460 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00484 vss n462 n461 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00483 n461 bshlmx_0_asr n460 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00482 vss bshlmx_0_lsl n463 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00481 n463 in_d_8 n462 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00480 bslmux_4_out_1 n448 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00479 vss n448 bslmux_4_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00478 bslmux_4_out_1 n448 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00477 vss n450 n437 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00476 n437 bshlmx_0_asr n448 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00475 vss bshlmx_0_lsl n438 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00474 n478 in_d_7 n489 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00473 bslmux_3_out_2 n496 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00472 vss n496 bslmux_3_out_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00471 bslmux_3_out_2 n496 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00470 vss n502 n497 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00469 n497 bshlmx_0_asr n496 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00468 vss bshlmx_0_lsl n503 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00467 n503 in_d_6 n502 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00466 bslmux_3_out_1 n490 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00465 vss n490 bslmux_3_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00464 bslmux_3_out_1 n490 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00463 vss n489 n477 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00462 n477 bshlmx_0_asr n490 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00461 vss bshlmx_0_lsl n478 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00460 n504 in_d_5 n519 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00459 bslmux_2_out_2 n540 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00458 vss n540 bslmux_2_out_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00457 bslmux_2_out_2 n540 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00456 vss n542 n541 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00455 n541 bshlmx_0_asr n540 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00454 vss bshlmx_0_lsl n543 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00453 n543 in_d_4 n542 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00452 bslmux_2_out_1 n529 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00451 vss n529 bslmux_2_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00450 bslmux_2_out_1 n529 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00449 vss n519 n518 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00448 n518 bshlmx_0_asr n529 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00447 vss bshlmx_0_lsl n504 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00446 n556 in_d_3 n569 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00445 bslmux_1_out_2 n580 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00444 vss n580 bslmux_1_out_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00443 bslmux_1_out_2 n580 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00442 vss n582 n581 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00441 n581 bshlmx_0_asr n580 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00440 vss bshlmx_0_lsl n583 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00439 n583 in_d_2 n582 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00438 bslmux_1_out_1 n568 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00437 vss n568 bslmux_1_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00436 bslmux_1_out_1 n568 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00435 vss n569 n555 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00434 n555 bshlmx_0_asr n568 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00433 vss bshlmx_0_lsl n556 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00432 n598 in_d_1 n610 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00431 bslmux_0_out_2 n688 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00430 vss n688 bslmux_0_out_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00429 bslmux_0_out_2 n688 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00428 vss n691 n689 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00427 n689 bshlmx_0_asr n688 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00426 vss bshlmx_0_lsl n692 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00425 n692 in_d_0 n691 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00424 bslmux_0_out_1 n608 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00423 vss n608 bslmux_0_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00422 bslmux_0_out_1 n608 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00421 vss n610 n597 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00420 n597 bshlmx_0_asr n608 vss TN L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00419 vss bshlmx_0_lsl n598 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00418 vss bsdand_15_out_2 n48 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00417 vss bssnbl_15_in_2 bssnbl_15_out_1 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00416 bssnbl_15_out_1 bssnbl_15_in_2 vss vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00415 bssnbl_15_out_1 bssnbl_15_in_2 vss vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00414 bslmux_15_com_2 n48 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00413 vss n48 bslmux_15_com_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00412 bslmux_15_com_2 n48 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00411 vss bsssel_14_out_2_s n86 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00410 vss bssnbl_14_in_1 n71 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00409 vss n71 bssnbl_14_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00408 bssnbl_14_out_1 n71 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00407 bssnbl_14_out_1 n71 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00406 bslmux_14_com_2 n86 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00405 vss n86 bslmux_14_com_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00404 bslmux_14_com_2 n86 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00403 vss bssnbl_13_in_2 n126 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00402 vss bssnbl_13_in_1 n109 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00401 vss n109 bssnbl_13_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00400 bssnbl_13_out_1 n109 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00399 bssnbl_13_out_1 n109 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00398 bslmux_13_com_2 n126 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00397 vss n126 bslmux_13_com_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00396 bslmux_13_com_2 n126 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00395 vss bssnbl_12_in_2 n161 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00394 vss bssnbl_12_in_1 n148 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00393 vss n148 bssnbl_12_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00392 bssnbl_12_out_1 n148 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00391 bssnbl_12_out_1 n148 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00390 bslmux_12_com_2 n161 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00389 vss n161 bslmux_12_com_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00388 bslmux_12_com_2 n161 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00387 vss bsssel_11_out_2_s n200 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00386 vss bsssel_11_out_1_s n184 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00385 vss n184 bssnbl_11_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00384 bssnbl_11_out_1 n184 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00383 bssnbl_11_out_1 n184 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00382 bslmux_11_com_2 n200 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00381 vss n200 bslmux_11_com_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00380 bslmux_11_com_2 n200 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00379 vss bsssel_10_out_2_s n238 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00378 vss bsssel_10_out_1_s n222 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00377 vss n222 bssnbl_10_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00376 bssnbl_10_out_1 n222 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00375 bssnbl_10_out_1 n222 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00374 bslmux_10_com_2 n238 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00373 vss n238 bslmux_10_com_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00372 bslmux_10_com_2 n238 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00371 vss bsssel_9_out_2_s n276 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00370 vss bssnbl_9_in_1 n261 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00369 vss n261 bssnbl_9_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00368 bssnbl_9_out_1 n261 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00367 bssnbl_9_out_1 n261 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00366 bslmux_9_com_2 n276 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00365 vss n276 bslmux_9_com_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00364 bslmux_9_com_2 n276 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00363 vss bssnbl_8_in_2 n316 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00362 vss bssnbl_8_in_1 n299 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00361 vss n299 bssnbl_8_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00360 bssnbl_8_out_1 n299 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00359 bssnbl_8_out_1 n299 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00358 bslmux_8_com_2 n316 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00357 vss n316 bslmux_8_com_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00356 bslmux_8_com_2 n316 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00355 vss bssnbl_7_in_2 n351 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00354 vss bssnbl_7_in_1 n338 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00353 vss n338 bssnbl_7_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00352 bssnbl_7_out_1 n338 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00351 bssnbl_7_out_1 n338 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00350 bslmux_7_com_2 n351 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00349 vss n351 bslmux_7_com_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00348 bslmux_7_com_2 n351 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00347 vss bsssel_6_out_2_s n390 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00346 vss bsssel_6_out_1_s n374 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00345 vss n374 bssnbl_6_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00344 bssnbl_6_out_1 n374 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00343 bssnbl_6_out_1 n374 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00342 bslmux_6_com_2 n390 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00341 vss n390 bslmux_6_com_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00340 bslmux_6_com_2 n390 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00339 vss bsssel_5_out_2_s n428 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00338 vss bsssel_5_out_1_s n412 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00337 vss n412 bssnbl_5_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00336 bssnbl_5_out_1 n412 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00335 bssnbl_5_out_1 n412 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00334 bslmux_5_com_2 n428 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00333 vss n428 bslmux_5_com_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00332 bslmux_5_com_2 n428 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00331 vss bsssel_4_out_2_s n464 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00330 vss bssnbl_4_in_1 n452 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00329 vss n452 bssnbl_4_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00328 bssnbl_4_out_1 n452 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00327 bssnbl_4_out_1 n452 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00326 bslmux_4_com_2 n464 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00325 vss n464 bslmux_4_com_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00324 bslmux_4_com_2 n464 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00323 vss bsssel_3_out_2_s n508 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00322 vss bssnbl_3_in_1 n492 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00321 vss n492 bssnbl_3_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00320 bssnbl_3_out_1 n492 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00319 bssnbl_3_out_1 n492 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00318 bslmux_3_com_2 n508 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00317 vss n508 bslmux_3_com_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00316 bslmux_3_com_2 n508 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00315 vss bssnbl_2_in_2 n558 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00314 vss bssnbl_2_in_1 n532 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00313 vss n532 bssnbl_2_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00312 bssnbl_2_out_1 n532 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00311 bssnbl_2_out_1 n532 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00310 bslmux_2_com_2 n558 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00309 vss n558 bslmux_2_com_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00308 bslmux_2_com_2 n558 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00307 vss bsssel_1_out_2_s n586 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00306 vss bsssel_1_out_1_s n570 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00305 vss n570 bssnbl_1_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00304 bssnbl_1_out_1 n570 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00303 bssnbl_1_out_1 n570 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00302 bslmux_1_com_2 n586 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00301 vss n586 bslmux_1_com_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00300 bslmux_1_com_2 n586 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00299 vss bsssel_0_out_2_s n696 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00298 vss bsssel_0_out_1_s n611 vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00297 vss n611 bssnbl_0_out_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00296 bssnbl_0_out_1 n611 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00295 bssnbl_0_out_1 n611 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00294 bssnbl_0_out_2 n696 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00293 vss n696 bssnbl_0_out_2 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00292 bssnbl_0_out_2 n696 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00291 bssnbl_15_zero n693 n20 vss TN L=0.18U W=3.06U AS=1.1016P AD=1.1016P 
+ PS=6.84U PD=6.84U 
Mtr_00290 n20 bsdand_15_out_1 vss vss TN L=0.18U W=3.06U AS=1.1016P AD=1.1016P 
+ PS=6.84U PD=6.84U 
Mtr_00289 bssnbl_15_in_2 bsdand_15_out_1 n47 vss TN L=0.18U W=3.06U AS=1.1016P 
+ AD=1.1016P PS=6.84U PD=6.84U 
Mtr_00288 n47 n699 vss vss TN L=0.18U W=3.06U AS=1.1016P AD=1.1016P PS=6.84U 
+ PD=6.84U 
Mtr_00287 bsdand_14_out_2 n693 bssnbl_14_in_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00286 bssnbl_14_in_1 n699 bsdand_14_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00285 bsssel_14_out_2_s n693 bsdand_14_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00284 bsdand_14_out_2 n699 bsssel_14_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00283 bsdand_13_out_2 n693 bssnbl_13_in_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00282 bssnbl_13_in_1 n699 bsdand_13_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00281 bssnbl_13_in_2 n693 bsdand_13_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00280 bsdand_13_out_2 n699 bssnbl_13_in_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00279 bsdand_12_out_2 n693 bssnbl_12_in_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00278 bssnbl_12_in_1 n699 bsdand_12_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00277 bssnbl_12_in_2 n693 bsdand_12_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00276 bsdand_12_out_2 n699 bssnbl_12_in_2 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00275 bsdand_11_out_2 n693 bsssel_11_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00274 bsssel_11_out_1_s n699 bsdand_11_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00273 bsssel_11_out_2_s n693 bsdand_11_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00272 bsdand_11_out_2 n699 bsssel_11_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00271 bsdand_10_out_2 n693 bsssel_10_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00270 bsssel_10_out_1_s n699 bsdand_10_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00269 bsssel_10_out_2_s n693 bsdand_10_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00268 bsdand_10_out_2 n699 bsssel_10_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00267 bsdand_9_out_2 n693 bssnbl_9_in_1 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00266 bssnbl_9_in_1 n699 bsdand_9_out_1 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00265 bsssel_9_out_2_s n693 bsdand_9_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00264 bsdand_9_out_2 n699 bsssel_9_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00263 bsdand_8_out_2 n693 bssnbl_8_in_1 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00262 bssnbl_8_in_1 n699 bsdand_8_out_1 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00261 bssnbl_8_in_2 n693 bsdand_8_out_1 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00260 bsdand_8_out_2 n699 bssnbl_8_in_2 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00259 bsdand_7_out_2 n693 bssnbl_7_in_1 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00258 bssnbl_7_in_1 n699 bsdand_7_out_1 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00257 bssnbl_7_in_2 n693 bsdand_7_out_1 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00256 bsdand_7_out_2 n699 bssnbl_7_in_2 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00255 bsdand_6_out_2 n693 bsssel_6_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00254 bsssel_6_out_1_s n699 bsdand_6_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00253 bsssel_6_out_2_s n693 bsdand_6_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00252 bsdand_6_out_2 n699 bsssel_6_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00251 bsdand_5_out_2 n693 bsssel_5_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00250 bsssel_5_out_1_s n699 bsdand_5_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00249 bsssel_5_out_2_s n693 bsdand_5_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00248 bsdand_5_out_2 n699 bsssel_5_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00247 bsdand_4_out_2 n693 bssnbl_4_in_1 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00246 bssnbl_4_in_1 n699 bsdand_4_out_1 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00245 bsssel_4_out_2_s n693 bsdand_4_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00244 bsdand_4_out_2 n699 bsssel_4_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00243 bsdand_3_out_2 n693 bssnbl_3_in_1 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00242 bssnbl_3_in_1 n699 bsdand_3_out_1 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00241 bsssel_3_out_2_s n693 bsdand_3_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00240 bsdand_3_out_2 n699 bsssel_3_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00239 bsdand_2_out_2 n693 bssnbl_2_in_1 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00238 bssnbl_2_in_1 n699 bsdand_2_out_1 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00237 bssnbl_2_in_2 n693 bsdand_2_out_1 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00236 bsdand_2_out_2 n699 bssnbl_2_in_2 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00235 bsdand_1_out_2 n693 bsssel_1_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00234 bsssel_1_out_1_s n699 bsdand_1_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00233 bsssel_1_out_2_s n693 bsdand_1_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00232 bsdand_1_out_2 n699 bsssel_1_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00231 bsdand_0_out_2 n693 bsssel_0_out_1_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00230 bsssel_0_out_1_s n699 bsdand_0_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00229 bsssel_0_out_2_s n693 bsdand_0_out_1 vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00228 bsdand_0_out_2 n699 bsssel_0_out_2_s vss TN L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00227 bsdand_15_out_1 n33 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00226 n33 bsdand_0_v_3_2 n22 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00225 n22 bsdand_0_v_4_2 n23 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00224 n23 bsdand_0_na1 n24 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00223 n24 bsdand_1_v_0_1 n21 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00222 n21 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00221 n50 bsdand_0_v_3_2 n51 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00220 n51 bsdand_0_v_4_1 n52 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00219 n52 bsdand_0_na1 n53 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00218 n53 bsdand_1_v_0_1 n54 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00217 n54 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00216 bsdand_15_out_2 n50 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00215 bsdand_14_out_1 n72 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00214 n72 bsdand_0_v_3_2 n62 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00213 n62 bsdand_0_v_4_1 n61 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00212 n61 bsdand_0_na1 n59 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00211 n59 bsdand_0_v_0_1 n60 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00210 n60 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00209 n89 bsdand_0_v_3_1 n90 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00208 n90 bsdand_0_v_4_2 n91 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00207 n91 bsdand_0_v_1_1 n92 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00206 n92 bsdand_0_v_0_1 n93 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00205 n93 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00204 bsdand_14_out_2 n89 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00203 bsdand_13_out_1 n110 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00202 n110 bsdand_0_v_3_2 n101 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00201 n101 bsdand_0_v_4_1 n100 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00200 n100 bsdand_0_v_1_1 n98 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00199 n98 bsdand_1_v_0_1 n99 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00198 n99 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00197 n131 bsdand_0_v_3_1 n132 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00196 n132 bsdand_0_v_4_2 n133 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00195 n133 bsdand_0_v_1_1 n134 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00194 n134 bsdand_1_v_0_1 n135 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00193 n135 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00192 bsdand_13_out_2 n131 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00191 bsdand_12_out_1 n149 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00190 n149 bsdand_0_v_3_2 n127 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00189 n127 bsdand_0_v_4_1 n128 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00188 n128 bsdand_0_v_1_1 n129 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00187 n129 bsdand_0_v_0_1 n130 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00186 n130 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00185 n165 bsdand_0_v_3_1 n166 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00184 n166 bsdand_0_v_4_2 n167 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00183 n167 bsdand_0_na1 n164 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00182 n164 bsdand_0_v_0_1 n163 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00181 n163 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00180 bsdand_12_out_2 n165 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00179 bsdand_11_out_1 n186 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00178 n186 bsdand_0_v_3_2 n174 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00177 n174 bsdand_0_v_4_1 n175 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00176 n175 bsdand_0_na1 n176 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00175 n176 bsdand_1_v_0_1 n173 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00174 n173 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00173 n204 bsdand_0_v_3_1 n205 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00172 n205 bsdand_0_v_4_2 n206 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00171 n206 bsdand_0_na1 n203 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00170 n203 bsdand_1_v_0_1 n202 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00169 n202 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00168 bsdand_11_out_2 n204 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00167 bsdand_10_out_1 n224 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00166 n224 bsdand_0_v_3_2 n212 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00165 n212 bsdand_0_v_4_1 n213 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00164 n213 bsdand_0_na1 n214 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00163 n214 bsdand_0_v_0_1 n211 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00162 n211 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00161 n240 bsdand_0_v_3_1 n241 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00160 n241 bsdand_0_v_4_2 n242 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00159 n242 bsdand_0_v_1_1 n243 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00158 n243 bsdand_0_v_0_1 n244 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00157 n244 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00156 bsdand_10_out_2 n240 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00155 bsdand_9_out_1 n262 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00154 n262 bsdand_0_v_3_2 n250 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00153 n250 bsdand_0_v_4_1 n251 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00152 n251 bsdand_0_v_1_1 n252 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00151 n252 bsdand_1_v_0_1 n249 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00150 n249 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00149 n279 bsdand_0_v_3_1 n280 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00148 n280 bsdand_0_v_4_2 n281 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00147 n281 bsdand_0_v_1_1 n282 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00146 n282 bsdand_1_v_0_1 n283 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00145 n283 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00144 bsdand_9_out_2 n279 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00143 bsdand_8_out_1 n300 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00142 n300 bsdand_0_v_3_2 n290 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00141 n290 bsdand_0_v_4_1 n289 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00140 n289 bsdand_0_v_1_1 n287 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00139 n287 bsdand_0_v_0_1 n288 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00138 n288 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00137 n317 bsdand_0_v_3_1 n318 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00136 n318 bsdand_0_v_4_2 n319 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00135 n319 bsdand_0_na1 n320 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00134 n320 bsdand_0_v_0_1 n321 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00133 n321 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00132 bsdand_8_out_2 n317 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00131 bsdand_7_out_1 n339 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00130 n339 bsdand_0_v_3_1 n329 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00129 n329 bsdand_0_v_4_1 n326 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00128 n326 bsdand_0_na1 n327 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00127 n327 bsdand_1_v_0_1 n328 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00126 n328 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00125 n355 bsdand_0_v_3_1 n356 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00124 n356 bsdand_0_v_4_2 n357 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00123 n357 bsdand_0_na1 n354 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00122 n354 bsdand_1_v_0_1 n353 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00121 n353 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00120 bsdand_7_out_2 n355 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00119 bsdand_6_out_1 n376 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00118 n376 bsdand_0_v_3_1 n364 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00117 n364 bsdand_0_v_4_1 n365 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00116 n365 bsdand_0_na1 n366 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00115 n366 bsdand_0_v_0_1 n363 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00114 n363 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00113 n394 bsdand_0_v_3_2 n395 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00112 n395 bsdand_0_v_4_2 n396 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00111 n396 bsdand_0_v_1_1 n393 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00110 n393 bsdand_0_v_0_1 n392 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00109 n392 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00108 bsdand_6_out_2 n394 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00107 bsdand_5_out_1 n414 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00106 n414 bsdand_0_v_3_1 n402 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00105 n402 bsdand_0_v_4_1 n403 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00104 n403 bsdand_0_v_1_1 n404 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00103 n404 bsdand_1_v_0_1 n401 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00102 n401 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00101 n430 bsdand_0_v_3_2 n431 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00100 n431 bsdand_0_v_4_2 n432 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00099 n432 bsdand_0_v_1_1 n433 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00098 n433 bsdand_1_v_0_1 n434 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00097 n434 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00096 bsdand_5_out_2 n430 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00095 bsdand_4_out_1 n453 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00094 n453 bsdand_0_v_3_1 n440 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00093 n440 bsdand_0_v_4_1 n441 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00092 n441 bsdand_0_v_1_1 n442 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00091 n442 bsdand_0_v_0_1 n439 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00090 n439 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00089 n468 bsdand_0_v_3_2 n469 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00088 n469 bsdand_0_v_4_2 n470 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00087 n470 bsdand_0_na1 n471 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00086 n471 bsdand_0_v_0_1 n472 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00085 n472 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00084 bsdand_4_out_2 n468 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00083 bsdand_3_out_1 n493 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00082 n493 bsdand_0_v_3_1 n482 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00081 n482 bsdand_0_v_4_1 n481 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00080 n481 bsdand_0_na1 n479 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00079 n479 bsdand_1_v_0_1 n480 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00078 n480 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00077 n509 bsdand_0_v_3_2 n510 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00076 n510 bsdand_0_v_4_2 n511 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00075 n511 bsdand_0_na1 n512 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00074 n512 bsdand_1_v_0_1 n513 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00073 n513 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00072 bsdand_3_out_2 n509 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00071 bsdand_2_out_1 n533 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00070 n533 bsdand_0_v_3_1 n523 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00069 n523 bsdand_0_v_4_1 n520 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00068 n520 bsdand_0_na1 n521 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00067 n521 bsdand_0_v_0_1 n522 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00066 n522 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00065 n548 bsdand_0_v_3_2 n549 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00064 n549 bsdand_0_v_4_2 n550 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00063 n550 bsdand_0_v_1_1 n547 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00062 n547 bsdand_0_v_0_1 n546 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00061 n546 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00060 bsdand_2_out_2 n548 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00059 bsdand_1_out_1 n572 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00058 n572 bsdand_0_v_3_1 n560 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00057 n560 bsdand_0_v_4_1 n561 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00056 n561 bsdand_0_v_1_1 n562 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00055 n562 bsdand_1_v_0_1 n559 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00054 n559 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00053 n590 bsdand_0_v_3_2 n591 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00052 n591 bsdand_0_v_4_2 n592 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00051 n592 bsdand_0_v_1_1 n589 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00050 n589 bsdand_1_v_0_1 n588 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00049 n588 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00048 bsdand_1_out_2 n590 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00047 bsdand_0_out_1 n613 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00046 n613 bsdand_0_v_3_1 n600 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00045 n600 bsdand_0_v_4_1 n601 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00044 n601 bsdand_0_v_1_1 n602 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00043 n602 bsdand_0_v_0_1 n599 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00042 n599 bsdand_0_v_2_1 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00041 n705 bsdand_0_v_3_2 n706 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00040 n706 bsdand_0_v_4_2 n707 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00039 n707 bsdand_0_na1 n704 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00038 n704 bsdand_0_v_0_1 n703 vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00037 n703 bsdand_0_v_2_2 vss vss TN L=0.18U W=2.7U AS=0.972P AD=0.972P 
+ PS=6.12U PD=6.12U 
Mtr_00036 bsdand_0_out_2 n705 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00035 bsdand_0_v_4_2 bsdand_0_v_4_1 vss vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00034 vss bsdand_0_v_4_1 bsdand_0_v_4_2 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00033 bsdand_0_v_4_1 n475 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00032 vss n475 bsdand_0_v_4_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00031 bsdand_0_v_4_1 n475 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00030 bsdand_0_v_4_2 bsdand_0_v_4_1 vss vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00029 vss in_s_4 n475 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_00028 bsdand_0_v_3_2 bsdand_0_v_3_1 vss vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00027 vss bsdand_0_v_3_1 bsdand_0_v_3_2 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00026 bsdand_0_v_3_1 n516 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00025 vss n516 bsdand_0_v_3_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00024 bsdand_0_v_3_1 n516 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00023 bsdand_0_v_3_2 bsdand_0_v_3_1 vss vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00022 vss in_s_3 n516 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_00021 bsdand_0_v_2_2 bsdand_0_v_2_1 vss vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00020 vss bsdand_0_v_2_1 bsdand_0_v_2_2 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00019 bsdand_0_v_2_1 n553 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00018 vss n553 bsdand_0_v_2_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00017 bsdand_0_v_2_1 n553 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00016 bsdand_0_v_2_2 bsdand_0_v_2_1 vss vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00015 vss in_s_2 n553 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_00014 bsdand_0_na1 bsdand_0_v_1_1 vss vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00013 vss bsdand_0_v_1_1 bsdand_0_na1 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00012 bsdand_0_v_1_1 n595 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00011 vss n595 bsdand_0_v_1_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00010 bsdand_0_v_1_1 n595 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00009 bsdand_0_na1 bsdand_0_v_1_1 vss vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00008 vss in_s_1 n595 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_00007 bsdand_1_v_0_1 bsdand_0_v_0_1 vss vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00006 vss bsdand_0_v_0_1 bsdand_1_v_0_1 vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00005 bsdand_0_v_0_1 n715 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00004 vss n715 bsdand_0_v_0_1 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00003 bsdand_0_v_0_1 n715 vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00002 bsdand_1_v_0_1 bsdand_0_v_0_1 vss vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00001 vss in_s_0 n715 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
.ends ex_shift32

