
.subckt ex_m8x8 a_0 a_1 a_2 a_3 a_4 a_5 a_6 a_7 b_0 b_1 b_2 b_3 b_4 b_5 b_6 
+ b_7 p_0 p_1 p_2 p_3 p_4 p_5 p_6 p_7 p_8 p_9 p_10 p_11 p_12 p_13 p_14 p_15 
+ vdd vss 
Mtr_01824 n884 c_4_1_sum n864 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01823 n864 cla_cell0_0_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01822 cla_cell0_0_g n880 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01821 vdd c_4_1_sum n880 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01820 n880 cla_cell0_0_a vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01819 vdd n880 cla_cell0_0_g vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01818 vdd n884 p_6 vdd TP L=0.18U W=1.98U AS=0.7128P AD=0.7128P PS=4.68U 
+ PD=4.68U 
Mtr_01817 n794 c_4_2_sum n793 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01816 n793 c_4_1_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01815 cla_cell0_1_g n791 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01814 vdd c_4_2_sum n791 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01813 n791 c_4_1_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01812 vdd n791 cla_cell0_1_g vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01811 vdd n794 cla_cell0_1_p vdd TP L=0.18U W=1.98U AS=0.7128P AD=0.7128P 
+ PS=4.68U PD=4.68U 
Mtr_01810 vdd n704 cla_cell0_2_g vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01809 n704 c_4_3_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01808 vdd c_4_2_cout n704 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01807 cla_cell0_2_g n704 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01806 vdd n708 cla_cell0_2_p vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_01805 cla_cell0_2_pn cla_cell0_2_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_01804 n652 c_4_3_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01803 n708 c_4_2_cout n652 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01802 n594 c_4_4_sum n650 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01801 n650 c_4_3_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01800 cla_cell0_3_g n651 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01799 vdd c_4_4_sum n651 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01798 n651 c_4_3_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01797 vdd n651 cla_cell0_3_g vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01796 vdd n594 cla_cell1_3_p1 vdd TP L=0.18U W=1.98U AS=0.7128P AD=0.7128P 
+ PS=4.68U PD=4.68U 
Mtr_01795 n542 c_4_4_cout n432 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01794 n432 c_4_5_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01793 cla_cell0_4_g n538 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01792 vdd c_4_4_cout n538 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01791 n538 c_4_5_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01790 vdd n538 cla_cell0_4_g vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01789 vdd n542 cla_cell3_4_p1 vdd TP L=0.18U W=1.98U AS=0.7128P AD=0.7128P 
+ PS=4.68U PD=4.68U 
Mtr_01788 vdd n431 cla_cell0_5_g vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01787 n431 c_4_5_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01786 vdd c_4_6_sum n431 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01785 cla_cell0_5_g n431 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01784 vdd n433 cla_cell1_5_p1 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_01783 cla_cell5_5_p cla_cell1_5_p1 vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_01782 n430 c_4_5_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01781 n433 c_4_6_sum n430 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01780 vdd n318 cla_cell1_6_tsg vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_01779 n318 c_4_7_sum vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01778 vdd c_4_6_cout n318 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01777 cla_cell1_6_tsg n318 vdd vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_01776 vdd n321 cla_cell0_6_p vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_01775 cla_cell5_6_p cla_cell0_6_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_01774 n202 c_4_7_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01773 n321 c_4_6_cout n202 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01772 vdd n200 cla_cell0_7_g vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01771 n200 c_4_7_cout vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01770 vdd c_4_8_sum n200 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01769 cla_cell0_7_g n200 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01768 vdd n204 cla_cell0_7_p vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_01767 cla_cell0_7_pn cla_cell0_7_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_01766 n199 c_4_7_cout vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01765 n204 c_4_8_sum n199 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01764 vdd n111 cla_cell0_8_g vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01763 n111 cla_cell0_8_a vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01762 vdd c_4_8_cout n111 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01761 cla_cell0_8_g n111 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01760 vdd n114 cla_cell0_8_p vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_01759 cla_cell5_8_p cla_cell0_8_p vdd vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_01758 n22 cla_cell0_8_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01757 n114 c_4_8_cout n22 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01756 n23 cla_cell0_8_a n21 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01755 n21 cla_cell0_9_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01754 cla_cell0_9_g n18 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01753 vdd cla_cell0_8_a n18 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01752 n18 cla_cell0_9_a vdd vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01751 vdd n18 cla_cell0_9_g vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01750 vdd n23 cla_cell0_9_p vdd TP L=0.18U W=1.98U AS=0.7128P AD=0.7128P 
+ PS=4.68U PD=4.68U 
Mtr_01749 vdd cla_cell0_0_g n788 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01748 n788 cla_cell0_1_p vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01747 cla_cell1_1_co cla_cell0_1_g n788 vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01746 vdd cla_cell0_2_g cla_cell1_2_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_01745 cla_cell1_2_np cla_cell0_2_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_01744 cla_cell1_3_g cla_cell0_3_g n649 vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01743 n649 cla_cell0_3_g cla_cell1_3_g vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01742 n649 cla_cell0_2_g vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01741 n649 cla_cell0_2_g vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01740 vdd cla_cell1_3_p1 n649 vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01739 n592 cla_cell0_2_p vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01738 vdd cla_cell0_2_p n592 vdd TP L=0.18U W=0.18U AS=0.0648P AD=0.0648P 
+ PS=1.08U PD=1.08U 
Mtr_01737 n592 cla_cell1_3_p1 vdd vdd TP L=0.18U W=0.18U AS=0.0648P AD=0.0648P 
+ PS=1.08U PD=1.08U 
Mtr_01736 n592 cla_cell1_3_p1 vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01735 cla_cell2_5_tsg cla_cell0_5_g n429 vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01734 n429 cla_cell0_5_g cla_cell2_5_tsg vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01733 n429 cla_cell0_4_g vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01732 n429 cla_cell0_4_g vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01731 vdd cla_cell1_5_p1 n429 vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01730 cla_cell2_5_tsp cla_cell3_4_p1 vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01729 vdd cla_cell3_4_p1 cla_cell2_5_tsp vdd TP L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_01728 cla_cell2_5_tsp cla_cell1_5_p1 vdd vdd TP L=0.18U W=0.18U AS=0.0648P 
+ AD=0.0648P PS=1.08U PD=1.08U 
Mtr_01727 cla_cell2_5_tsp cla_cell1_5_p1 vdd vdd TP L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_01726 vdd cla_cell1_6_tsg cla_cell1_6_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_01725 cla_cell1_6_np cla_cell0_6_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_01724 cla_cell1_7_g cla_cell0_7_g n198 vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_01723 n198 cla_cell0_7_g cla_cell1_7_g vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_01722 n198 cla_cell1_6_tsg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_01721 n198 cla_cell1_6_tsg vdd vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_01720 cla_cell2_7_pl cla_cell0_6_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_01719 vdd cla_cell0_7_p n198 vdd TP L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01718 cla_cell2_7_pl cla_cell0_7_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_01717 vdd cla_cell0_8_g cla_cell1_8_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_01716 cla_cell1_8_np cla_cell0_8_p vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_01715 cla_cell1_9_g cla_cell0_9_g n17 vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_01714 n17 cla_cell0_9_g cla_cell1_9_g vdd TP L=0.18U W=0.36U AS=0.1296P 
+ AD=0.1296P PS=1.44U PD=1.44U 
Mtr_01713 n17 cla_cell0_8_g vdd vdd TP L=0.18U W=0.36U AS=0.1296P AD=0.1296P 
+ PS=1.44U PD=1.44U 
Mtr_01712 n17 cla_cell0_8_g vdd vdd TP L=0.18U W=0.36U AS=0.1296P AD=0.1296P 
+ PS=1.44U PD=1.44U 
Mtr_01711 n15 cla_cell0_8_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P AD=0.2592P 
+ PS=2.16U PD=2.16U 
Mtr_01710 vdd cla_cell0_9_p n17 vdd TP L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01709 n15 cla_cell0_9_p vdd vdd TP L=0.18U W=0.72U AS=0.2592P AD=0.2592P 
+ PS=2.16U PD=2.16U 
Mtr_01708 vdd cla_cell1_2_ng cla_cell5_2_g vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_01707 cla_cell5_2_g cla_cell1_2_np n647 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_01706 n647 cla_cell1_1_co vdd vdd TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01705 vdd n592 n589 vdd TP L=0.18U W=4.5U AS=1.62P AD=1.62P PS=9.72U 
+ PD=9.72U 
Mtr_01704 n589 cla_cell1_1_co cla_cell3_4_g2 vdd TP L=0.18U W=4.5U AS=1.62P 
+ AD=1.62P PS=9.72U PD=9.72U 
Mtr_01703 cla_cell3_4_g2 cla_cell1_3_g vdd vdd TP L=0.18U W=2.34U AS=0.8424P 
+ AD=0.8424P PS=5.4U PD=5.4U 
Mtr_01702 vdd cla_cell2_5_tsg cla_cell2_5_ng vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_01701 cla_cell2_5_np cla_cell2_5_tsp vdd vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_01700 n288 cla_cell1_6_np vdd vdd TP L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01699 cla_cell3_6_p1 cla_cell2_5_tsp n288 vdd TP L=0.18U W=1.26U 
+ AS=0.4536P AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01698 vdd cla_cell1_6_np n195 vdd TP L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01697 n195 cla_cell2_5_tsg cla_cell2_6_g vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01696 cla_cell2_6_g cla_cell1_6_ng vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_01695 n162 cla_cell2_7_pl vdd vdd TP L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01694 n192 cla_cell2_5_tsp n162 vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01693 vdd cla_cell2_7_pl n194 vdd TP L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_01692 n194 cla_cell2_5_tsg cla_cell2_7_g vdd TP L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_01691 cla_cell2_7_g cla_cell1_7_g vdd vdd TP L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_01690 vdd cla_cell3_4_g2 n497 vdd TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01689 n497 cla_cell3_4_p1 vdd vdd TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01688 cla_cell3_4_co cla_cell0_4_g n497 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_01687 vdd cla_cell3_4_g2 n424 vdd TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01686 n424 cla_cell2_5_np vdd vdd TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01685 cla_cell3_5_co cla_cell2_5_ng n424 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_01684 vdd cla_cell3_4_g2 n287 vdd TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01683 n287 cla_cell3_6_p1 vdd vdd TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01682 cla_cell3_6_co cla_cell2_6_g n287 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_01681 vdd cla_cell3_4_g2 n191 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01680 n191 n192 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_01679 cla_cell3_7_co cla_cell2_7_g n191 vdd TP L=0.18U W=3.6U AS=1.296P 
+ AD=1.296P PS=7.92U PD=7.92U 
Mtr_01678 vdd cla_cell1_8_ng cla_cell5_8_g vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_01677 cla_cell5_8_g cla_cell1_8_np n78 vdd TP L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_01676 n78 cla_cell3_7_co vdd vdd TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01675 vdd cla_cell1_9_g n14 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01674 n14 n15 n13 vdd TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P PS=6.48U 
+ PD=6.48U 
Mtr_01673 n13 cla_cell3_7_co vdd vdd TP L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_01672 n787 cla_cell0_1_p n786 vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01671 n786 cla_cell0_0_g vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01670 p_7 n787 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_01669 n646 cla_cell1_1_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01668 n697 cla_cell0_2_pn n646 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_01667 p_8 n697 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_01666 n645 cla_cell1_3_p1 n588 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_01665 n588 cla_cell5_2_g vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01664 p_9 n645 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_01663 n423 cla_cell3_4_g2 vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01662 n531 cla_cell3_4_p1 n423 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_01661 p_10 n531 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_01660 n421 cla_cell5_5_p n422 vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01659 n422 cla_cell3_4_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01658 p_11 n421 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_01657 n188 cla_cell3_5_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01656 n304 cla_cell5_6_p n188 vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01655 p_12 n304 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_01654 n190 cla_cell0_7_pn n189 vdd TP L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_01653 n189 cla_cell3_6_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01652 p_13 n190 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_01651 n77 cla_cell3_7_co vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01650 n101 cla_cell5_8_p n77 vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01649 p_14 n101 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_01648 n11 cla_cell0_9_p n12 vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01647 n12 cla_cell5_8_g vdd vdd TP L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_01646 p_15 n11 vdd vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_01645 cla_cell0_8_a n26 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01644 n34 n30 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01643 cla_cell0_9_a n35 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01642 n25 c_4_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01641 vdd p_4_9_pi2j n25 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01640 n35 c_4_8_cin n25 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01639 n35 c_4_7_a n33 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01638 n33 p_4_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01637 n26 c_4_8_cin n34 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01636 vdd n32 n30 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P PS=3.6U 
+ PD=3.6U 
Mtr_01635 n32 c_4_7_a n31 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01634 n31 p_4_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01633 n39 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01632 vdd p_4_9_t_s n29 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01631 n29 p_4_1_n2j p_4_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01630 vdd n39 n36 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01629 n36 n40 p_4_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01628 n40 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01627 vdd n126 n83 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01626 n82 p_4_1_n2j p_4_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01625 vdd p_4_8_t_s n82 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01624 vdd a_6 n84 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01623 n85 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01622 n128 p_4_2_d2j n85 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01621 n84 p_4_2_d2jbar n128 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01620 n126 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01619 n83 n128 p_4_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01618 vdd c_4_7_a n80 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01617 c_4_8_sum c_4_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01616 n81 n116 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01615 c_4_8_cout n120 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01614 n80 p_4_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01613 n120 c_4_8_cin n80 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01612 n120 p_4_8_pi2j n28 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01611 n28 c_4_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01610 c_4_8_s2_s c_4_8_cin n81 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01609 vdd c_4_8_s1_s n116 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01608 c_4_8_s1_s p_4_8_pi2j n27 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01607 n27 c_4_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01606 c_4_7_sum c_4_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01605 n219 n216 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01604 c_4_7_cout n221 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01603 n209 c_4_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01602 vdd p_4_7_pi2j n209 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01601 n221 c_4_7_cin n209 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01600 n221 c_4_7_a n218 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01599 n218 p_4_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01598 c_4_7_s2_s c_4_7_cin n219 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01597 vdd c_4_7_s1_s n216 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01596 c_4_7_s1_s c_4_7_a n217 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01595 n217 p_4_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01594 n166 p_4_2_d2j n222 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01593 n222 p_4_2_d2jbar n165 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01592 n165 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01591 vdd a_6 n166 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01590 vdd p_4_7_t_s n214 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01589 n214 p_4_1_n2j p_4_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01588 vdd n222 n223 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01587 n223 n227 p_4_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01586 n227 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01585 vdd n335 n224 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01584 n215 p_4_1_n2j p_4_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01583 vdd p_4_6_t_s n215 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01582 vdd a_4 n228 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01581 n229 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01580 n333 p_4_2_d2j n229 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01579 n228 p_4_2_d2jbar n333 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01578 n335 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01577 n224 n333 p_4_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01576 vdd c_4_6_a n289 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01575 c_4_6_sum c_4_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01574 n290 n291 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01573 c_4_6_cout n329 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01572 n289 p_4_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01571 n329 c_4_6_cin n289 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01570 n329 p_4_6_pi2j n212 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01569 n212 c_4_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01568 c_4_6_s2_s c_4_6_cin n290 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01567 vdd c_4_6_s1_s n291 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01566 c_4_6_s1_s p_4_6_pi2j n213 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01565 n213 c_4_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01564 c_4_5_sum c_4_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01563 n392 n393 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01562 c_4_5_cout n446 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01561 n437 c_4_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01560 vdd c_4_5_b n437 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01559 n446 c_4_5_cin n437 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01558 n446 c_4_5_a n445 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01557 n445 c_4_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01556 c_4_5_s2_s c_4_5_cin n392 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01555 vdd c_4_5_s1_s n393 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01554 c_4_5_s1_s c_4_5_a n444 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01553 n444 c_4_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01552 n396 p_4_2_d2j n447 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01551 n447 p_4_2_d2jbar n395 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01550 n395 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01549 vdd a_4 n396 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01548 vdd p_4_5_t_s n391 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01547 n391 p_4_1_n2j c_4_5_b vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01546 vdd n447 n394 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01545 n394 n450 p_4_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01544 n450 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01543 vdd n505 n449 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01542 n442 p_4_1_n2j p_4_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01541 vdd p_4_4_t_s n442 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01540 vdd a_2 n451 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01539 n452 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01538 n508 p_4_2_d2j n452 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01537 n451 p_4_2_d2jbar n508 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01536 n505 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01535 n449 n508 p_4_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01534 vdd c_4_4_a n436 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01533 c_4_4_sum c_4_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01532 n501 n502 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01531 c_4_4_cout n499 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01530 n436 p_4_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01529 n499 c_4_4_cin n436 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01528 n499 p_4_4_pi2j n441 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01527 n441 c_4_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01526 c_4_4_s2_s c_4_4_cin n501 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01525 vdd c_4_4_s1_s n502 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01524 c_4_4_s1_s p_4_4_pi2j n440 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01523 n440 c_4_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01522 c_4_3_sum c_4_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01521 n601 n603 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01520 c_4_3_cout n600 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01519 n655 c_4_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01518 vdd c_4_3_b n655 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01517 n600 c_4_3_cin n655 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01516 n600 c_4_3_a n661 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01515 n661 c_4_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01514 c_4_3_s2_s c_4_3_cin n601 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01513 vdd c_4_3_s1_s n603 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01512 c_4_3_s1_s c_4_3_a n662 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01511 n662 c_4_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01510 n607 p_4_2_d2j n605 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01509 n605 p_4_2_d2jbar n606 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01508 n606 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01507 vdd a_2 n607 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01506 vdd p_4_3_t_s n599 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01505 n599 p_4_1_n2j c_4_3_b vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01504 vdd n605 n604 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01503 n604 n608 p_4_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01502 n608 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01501 vdd n718 n664 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01500 n660 p_4_1_n2j c_4_2_b vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01499 vdd p_4_2_t_s n660 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01498 vdd a_0 n665 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01497 n666 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01496 n721 p_4_2_d2j n666 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01495 n665 p_4_2_d2jbar n721 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01494 n718 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01493 n664 n721 p_4_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01492 vdd c_4_2_a n654 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01491 c_4_2_sum c_4_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01490 n658 n714 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01489 c_4_2_cout n712 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01488 n654 c_4_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01487 n712 c_4_2_cin n654 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01486 n712 c_4_2_b n659 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01485 n659 c_4_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01484 c_4_2_s2_s c_4_2_cin n658 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01483 vdd c_4_2_s1_s n714 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01482 c_4_2_s1_s c_4_2_b n657 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01481 n657 c_4_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01480 c_4_1_sum c_4_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01479 n806 n804 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01478 c_4_1_cout n805 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01477 n798 c_4_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01476 vdd p_4_1_pi2j n798 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01475 n805 c_4_1_cin n798 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01474 n805 c_4_1_a n807 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01473 n807 p_4_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01472 c_4_1_s2_s c_4_1_cin n806 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01471 vdd c_4_1_s1_s n804 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01470 c_4_1_s1_s c_4_1_a n801 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01469 n801 p_4_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01468 n815 p_4_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01467 vdd a_0 n815 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01466 vdd p_4_1_t_s n802 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01465 n802 p_4_1_n2j p_4_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01464 vdd n815 n809 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01463 n809 n814 p_4_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01462 n814 p_4_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01461 n869 c_3_1_sum cl4_4_s1_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01460 vdd n908 n869 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01459 p_4 cl4_4_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01458 n897 c_3_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01457 vdd n908 n897 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01456 n896 n897 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01455 n893 c_3_1_cout n867 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01454 n867 c_3_2_sum n893 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01453 n868 c_3_2_sum n867 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01452 vdd c_3_1_cout n868 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01451 n867 c_3_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01450 vdd n908 n867 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01449 cla_cell0_0_a n893 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01448 n866 c_3_2_sum cl4_4_s2_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01447 vdd c_3_1_cout n866 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01446 n888 cl4_4_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01445 n865 n896 cl4_4_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01444 vdd n888 n865 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01443 p_5 cl4_4_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01442 n50 p_3_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01441 c_3_9_s1_s c_3_7_a n50 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01440 vdd c_3_9_s1_s n51 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01439 c_3_9_s2_s c_3_8_cin n43 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01438 n44 p_3_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01437 n42 c_3_7_a n44 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01436 n42 c_3_8_cin n46 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01435 vdd p_3_9_pi2j n46 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01434 n46 c_3_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01433 c_4_8_cin n42 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01432 n43 n51 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01431 c_4_7_a c_3_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01430 n56 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01429 vdd p_3_9_t_s n49 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01428 n49 p_3_1_n2j p_3_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01427 vdd n56 n55 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01426 n55 n53 p_3_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01425 n53 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01424 vdd n141 n89 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01423 n88 p_3_1_n2j p_3_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01422 vdd p_3_8_t_s n88 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01421 vdd a_6 n90 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01420 n91 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01419 n143 p_3_2_d2j n91 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01418 n90 p_3_2_d2jbar n143 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01417 n141 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01416 n89 n143 p_3_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01415 n47 c_3_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01414 c_3_8_s1_s p_3_8_pi2j n47 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01413 vdd c_3_8_s1_s n134 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01412 c_3_8_s2_s c_3_8_cin n87 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01411 n41 c_3_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01410 n132 p_3_8_pi2j n41 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01409 n132 c_3_8_cin n86 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01408 vdd c_3_7_a n86 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01407 n86 p_3_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01406 c_4_7_cin n132 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01405 n87 n134 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01404 c_4_6_a c_3_8_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01403 c_4_5_a c_3_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01402 n232 n243 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01401 c_4_6_cin n234 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01400 n236 c_3_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01399 vdd p_3_7_pi2j n236 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01398 n234 c_3_7_cin n236 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01397 n234 c_3_7_a n233 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01396 n233 p_3_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01395 c_3_7_s2_s c_3_7_cin n232 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01394 vdd c_3_7_s1_s n243 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01393 c_3_7_s1_s c_3_7_a n244 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01392 n244 p_3_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01391 n171 p_3_2_d2j n245 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01390 n245 p_3_2_d2jbar n170 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01389 n170 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01388 vdd a_6 n171 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01387 vdd p_3_7_t_s n241 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01386 n241 p_3_1_n2j p_3_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01385 vdd n245 n248 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01384 n248 n246 p_3_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01383 n246 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01382 vdd n348 n249 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01381 n239 p_3_1_n2j p_3_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01380 vdd p_3_6_t_s n239 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01379 vdd a_4 n250 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01378 n251 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01377 n347 p_3_2_d2j n251 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01376 n250 p_3_2_d2jbar n347 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01375 n348 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01374 n249 n347 p_3_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01373 n238 c_3_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01372 c_3_6_s1_s p_3_6_pi2j n238 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01371 vdd c_3_6_s1_s n296 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01370 c_3_6_s2_s c_2_7_cout n294 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01369 n231 c_3_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01368 n341 p_3_6_pi2j n231 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01367 n341 c_2_7_cout n295 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01366 vdd c_3_6_a n295 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01365 n295 p_3_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01364 c_4_5_cin n341 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01363 n294 n296 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01362 c_4_4_a c_3_6_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01361 c_4_3_a c_3_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01360 n398 n402 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01359 c_4_4_cin n456 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01358 n457 c_3_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01357 vdd c_3_5_b n457 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01356 n456 c_3_5_cin n457 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01355 n456 c_3_5_a n455 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01354 n455 c_3_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01353 c_3_5_s2_s c_3_5_cin n398 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01352 vdd c_3_5_s1_s n402 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01351 c_3_5_s1_s c_3_5_a n462 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01350 n462 c_3_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01349 n405 p_3_2_d2j n466 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01348 n466 p_3_2_d2jbar n404 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01347 n404 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01346 vdd a_4 n405 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01345 vdd p_3_5_t_s n401 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01344 n401 p_3_1_n2j c_3_5_b vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01343 vdd n466 n403 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01342 n403 n465 p_3_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01341 n465 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01340 vdd n515 n467 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01339 n463 p_3_1_n2j p_3_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01338 vdd p_3_4_t_s n463 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01337 vdd a_2 n468 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01336 n469 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01335 n517 p_3_2_d2j n469 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01334 n468 p_3_2_d2jbar n517 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01333 n515 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01332 n467 n517 p_3_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01331 n460 c_3_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01330 c_3_4_s1_s p_3_4_pi2j n460 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01329 vdd c_3_4_s1_s n514 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01328 c_3_4_s2_s c_2_5_cout n510 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01327 n453 c_3_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01326 n509 p_3_4_pi2j n453 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01325 n509 c_2_5_cout n454 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01324 vdd c_3_4_a n454 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01323 n454 p_3_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01322 c_4_3_cin n509 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01321 n510 n514 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01320 c_4_2_a c_3_4_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01319 c_4_1_a c_3_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01318 n609 n616 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01317 c_4_2_cin n610 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01316 n670 c_3_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01315 vdd c_3_3_b n670 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01314 n610 c_3_3_cin n670 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01313 n610 c_3_3_a n671 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01312 n671 c_3_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01311 c_3_3_s2_s c_3_3_cin n609 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01310 vdd c_3_3_s1_s n616 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01309 c_3_3_s1_s c_3_3_a n674 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01308 n674 c_3_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01307 n621 p_3_2_d2j n619 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01306 n619 p_3_2_d2jbar n620 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01305 n620 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01304 vdd a_2 n621 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01303 vdd p_3_3_t_s n614 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01302 n614 p_3_1_n2j c_3_3_b vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01301 vdd n619 n618 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01300 n618 n617 p_3_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01299 n617 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01298 vdd n731 n677 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01297 n675 p_3_1_n2j c_3_2_b vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01296 vdd p_3_2_t_s n675 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01295 vdd a_0 n678 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01294 n679 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01293 n733 p_3_2_d2j n679 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01292 n678 p_3_2_d2jbar n733 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01291 n731 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01290 n677 n733 p_3_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01289 n673 c_3_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01288 c_3_2_s1_s c_3_2_b n673 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01287 vdd c_3_2_s1_s n727 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01286 c_3_2_s2_s c_2_3_cout n669 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01285 n667 c_3_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01284 n724 c_3_2_b n667 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01283 n724 c_2_3_cout n668 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01282 vdd c_3_2_a n668 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01281 n668 c_3_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01280 c_4_1_cin n724 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01279 n669 n727 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01278 c_3_2_sum c_3_2_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01277 c_3_1_sum c_3_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01276 n818 n826 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01275 c_3_1_cout n819 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01274 n821 c_3_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01273 vdd p_3_1_pi2j n821 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01272 n819 c_3_1_cin n821 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01271 n819 c_3_1_a n817 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01270 n817 p_3_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01269 c_3_1_s2_s c_3_1_cin n818 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01268 vdd c_3_1_s1_s n826 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01267 c_3_1_s1_s c_3_1_a n827 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01266 n827 p_3_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01265 n834 p_3_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01264 vdd a_0 n834 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01263 vdd p_3_1_t_s n824 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01262 n824 p_3_1_n2j p_3_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01261 vdd n834 n831 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01260 n831 n830 p_3_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01259 n830 p_3_1_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01258 n874 c_2_1_sum cl4_3_s1_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01257 vdd n922 n874 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01256 p_2 cl4_3_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01255 n913 c_2_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01254 vdd n922 n913 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01253 n914 n913 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01252 n910 c_2_1_cout n873 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01251 n873 c_2_2_sum n910 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01250 n872 c_2_2_sum n873 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01249 vdd c_2_1_cout n872 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01248 n873 c_2_1_sum vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01247 vdd n922 n873 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01246 n908 n910 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01245 n871 c_2_2_sum cl4_3_s2_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01244 vdd c_2_1_cout n871 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01243 n906 cl4_3_s2_s vdd vdd TP L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_01242 n870 n914 cl4_3_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01241 vdd n906 n870 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01240 p_3 cl4_3_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01239 c_3_7_a c_2_9_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01238 n58 n64 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01237 c_3_8_cin n60 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01236 n57 c_2_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01235 vdd p_2_9_pi2j n57 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01234 n60 vss n57 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01233 n60 c_2_7_a n59 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01232 n59 p_2_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01231 c_2_9_s2_s vss n58 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01230 vdd c_2_9_s1_s n64 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01229 c_2_9_s1_s c_2_7_a n65 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01228 n65 p_2_9_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01227 n72 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01226 vdd p_2_9_t_s n63 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01225 n63 p_2_1_n2j p_2_9_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01224 vdd n72 n70 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01223 n70 n68 p_2_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01222 n68 n847 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01221 vdd n150 n93 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01220 n92 p_2_1_n2j p_2_8_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01219 vdd p_2_8_t_s n92 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01218 vdd a_6 n95 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01217 n94 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01216 n153 p_2_2_d2j n94 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01215 n95 p_2_2_d2jbar n153 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01214 n150 n847 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01213 n93 n153 p_2_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01212 vdd c_2_8_s1_s c_3_6_a vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01211 n146 p_2_8_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01210 vdd c_2_7_a n146 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01209 c_3_7_cin n146 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01208 c_2_8_s1_s p_2_8_pi2j n62 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01207 n62 c_2_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01206 c_3_5_a c_2_7_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01205 n254 n261 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01204 c_2_7_cout n253 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01203 n252 c_2_7_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01202 vdd p_2_7_pi2j n252 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01201 n253 vss n252 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01200 n253 c_2_7_a n255 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01199 n255 p_2_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01198 c_2_7_s2_s vss n254 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01197 vdd c_2_7_s1_s n261 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01196 c_2_7_s1_s c_2_7_a n263 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01195 n263 p_2_7_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01194 n175 p_2_2_d2j n265 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01193 n265 p_2_2_d2jbar n176 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01192 n176 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01191 vdd a_6 n175 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01190 vdd p_2_7_t_s n260 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01189 n260 p_2_1_n2j p_2_7_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01188 vdd n265 n268 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01187 n268 n266 p_2_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01186 n266 n847 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01185 vdd n360 n269 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01184 n259 p_2_1_n2j p_2_6_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01183 vdd p_2_6_t_s n259 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01182 vdd a_4 n272 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01181 n271 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01180 n359 p_2_2_d2j n271 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01179 n272 p_2_2_d2jbar n359 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01178 n360 n847 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01177 n269 n359 p_2_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01176 vdd c_2_6_s1_s c_3_4_a vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01175 n354 p_2_6_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01174 vdd c_2_6_a n354 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01173 c_3_5_cin n354 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01172 c_2_6_s1_s p_2_6_pi2j n258 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01171 n258 c_2_6_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01170 c_3_3_a c_2_5_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01169 n407 n409 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01168 c_2_5_cout n472 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01167 n470 c_2_5_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01166 vdd c_2_5_b n470 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01165 n472 p_4_1_c2j n470 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01164 n472 c_2_5_a n471 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01163 n471 c_2_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01162 c_2_5_s2_s p_4_1_c2j n407 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01161 vdd c_2_5_s1_s n409 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01160 c_2_5_s1_s c_2_5_a n478 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01159 n478 c_2_5_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01158 n413 p_2_2_d2j n479 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01157 n479 p_2_2_d2jbar n414 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01156 n414 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01155 vdd a_4 n413 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01154 vdd p_2_5_t_s n410 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01153 n410 p_2_1_n2j c_2_5_b vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01152 vdd n479 n411 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01151 n411 n480 p_2_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01150 n480 n847 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01149 vdd n520 n482 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01148 n476 p_2_1_n2j p_2_4_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01147 vdd p_2_4_t_s n476 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01146 vdd a_2 n484 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01145 n483 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01144 n523 p_2_2_d2j n483 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01143 n484 p_2_2_d2jbar n523 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01142 n520 n847 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01141 n482 n523 p_2_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01140 vdd c_2_4_s1_s c_3_2_a vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01139 n562 p_2_4_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01138 vdd c_2_4_a n562 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01137 c_3_3_cin n562 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01136 c_2_4_s1_s p_2_4_pi2j n475 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01135 n475 c_2_4_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01134 c_3_1_a c_2_3_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01133 n622 n627 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01132 c_2_3_cout n623 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01131 n680 c_2_3_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01130 vdd c_2_3_b n680 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01129 n623 p_3_1_c2j n680 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01128 n623 c_2_3_a n681 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01127 n681 c_2_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01126 c_2_3_s2_s p_3_1_c2j n622 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01125 vdd c_2_3_s1_s n627 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01124 c_2_3_s1_s c_2_3_a n684 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01123 n684 c_2_3_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01122 n632 p_2_2_d2j n634 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01121 n634 p_2_2_d2jbar n633 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01120 n633 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01119 vdd a_2 n632 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01118 vdd p_2_3_t_s n626 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01117 n626 p_2_1_n2j c_2_3_b vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01116 vdd n634 n629 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01115 n629 n630 p_2_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01114 n630 n847 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01113 vdd n739 n687 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01112 n685 p_2_1_n2j c_2_2_b vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01111 vdd p_2_2_t_s n685 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01110 vdd a_0 n689 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01109 n688 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01108 n743 p_2_2_d2j n688 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01107 n689 p_2_2_d2jbar n743 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01106 n739 n847 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01105 n687 n743 p_2_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01104 vdd c_2_2_s1_s c_2_2_sum vdd TP L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_01103 n736 c_2_2_b vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01102 vdd c_2_2_a n736 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01101 c_3_1_cin n736 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01100 c_2_2_s1_s c_2_2_b n683 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01099 n683 c_2_2_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01098 c_2_1_sum c_2_1_s2_s vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01097 n837 n844 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01096 c_2_1_cout n836 vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01095 n835 c_2_1_a vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01094 vdd p_2_1_pi2j n835 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01093 n836 n847 n835 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01092 n836 c_2_1_a n838 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01091 n838 p_2_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01090 c_2_1_s2_s n847 n837 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01089 vdd c_2_1_s1_s n844 vdd TP L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_01088 c_2_1_s1_s c_2_1_a n845 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01087 n845 p_2_1_pi2j vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01086 n849 n847 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01085 n848 n849 p_2_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01084 vdd n853 n848 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01083 n843 p_2_1_n2j p_2_1_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_01082 vdd p_2_1_t_s n843 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01081 vdd a_0 n853 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01080 n853 p_2_2_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01079 n876 n932 cl4_2_s1_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01078 vdd p_1_2_c2j n876 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01077 p_0 cl4_2_s1_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01076 n926 n932 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01075 vdd p_1_2_c2j n926 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01074 n927 n926 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01073 vdd p_1_2_pi2j n923 vdd TP L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_01072 n923 n932 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01071 vdd p_1_2_c2j n923 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01070 n922 n923 vdd vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P PS=4.32U 
+ PD=4.32U 
Mtr_01069 n875 n927 cl4_2_s3_s vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01068 vdd p_1_2_pi2j n875 vdd TP L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_01067 p_1 cl4_2_s3_s vdd vdd TP L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_01066 p_1_9_a a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01065 vdd p_1_9_t_s n71 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01064 n71 d_0_n2j c_2_7_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01063 vdd p_1_9_a n73 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01062 n73 n76 p_1_9_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01061 n76 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01060 vdd d_0_n2j n96 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01059 vdd n157 n97 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01058 n157 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01057 vdd a_6 n98 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01056 n155 d_0_d2j n99 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01055 n99 a_7 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01054 n98 d_0_d2jbar n155 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01053 n96 p_1_8_t_s c_2_6_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01052 n97 n155 p_1_8_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01051 n273 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01050 n278 n273 p_1_7_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01049 vdd p_1_7_a n278 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01048 n270 d_0_n2j c_2_5_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01047 vdd p_1_7_t_s n270 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01046 vdd a_6 n180 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01045 n179 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01044 p_1_7_a d_0_d2jbar n179 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01043 n180 d_0_d2j p_1_7_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01042 vdd d_0_n2j n275 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01041 vdd n365 n276 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01040 n365 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01039 vdd a_4 n280 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01038 n363 d_0_d2j n281 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01037 n281 a_5 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01036 n280 d_0_d2jbar n363 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01035 n275 p_1_6_t_s c_2_4_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01034 n276 n363 p_1_6_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01033 n486 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01032 n415 n486 p_1_5_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01031 vdd p_1_5_a n415 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01030 n412 d_0_n2j c_2_3_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01029 vdd p_1_5_t_s n412 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01028 vdd a_4 n418 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01027 n417 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01026 p_1_5_a d_0_d2jbar n417 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01025 n418 d_0_d2j p_1_5_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01024 vdd d_0_n2j n487 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01023 vdd n524 n488 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01022 n524 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01021 vdd a_2 n489 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01020 n527 d_0_d2j n490 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01019 n490 a_3 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01018 n489 d_0_d2jbar n527 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01017 n487 p_1_4_t_s c_2_2_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01016 n488 n527 p_1_4_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01015 n690 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01014 n635 n690 p_1_3_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01013 vdd p_1_3_a n635 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01012 n631 d_0_n2j c_2_1_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01011 vdd p_1_3_t_s n631 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01010 vdd a_2 n639 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01009 n638 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01008 p_1_3_a d_0_d2jbar n638 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01007 n639 d_0_d2j p_1_3_a vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01006 vdd d_0_n2j n691 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01005 vdd n745 n692 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01004 n745 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01003 vdd a_0 n693 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01002 n748 d_0_d2j n694 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_01001 n694 a_1 vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_01000 n693 d_0_d2jbar n748 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00999 n691 p_1_2_t_s p_1_2_pi2j vdd TP L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00998 n692 n748 p_1_2_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00997 n857 d_0_d2jbar vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00996 vdd a_0 n857 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00995 vdd p_1_1_t_s n852 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00994 n852 d_0_n2j n932 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00993 vdd n857 n855 vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00992 n855 n856 p_1_1_t_s vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00991 n856 p_1_2_c2j vdd vdd TP L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00990 n285 n369 n286 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00989 n286 b_7 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00988 vdd b_7 n283 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00987 n283 n376 n282 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00986 n282 n374 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00985 vdd b_5 n286 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00984 n286 n374 n285 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00983 n285 n376 n286 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00982 n286 b_6 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00981 vdd p_4_2_d2j p_4_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_00980 p_4_1_c2j n283 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00979 vdd n285 p_4_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00978 p_4_2_d2j n381 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00977 n369 b_7 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00976 vdd n369 n284 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00975 n284 b_7 n381 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00974 n374 b_5 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00973 n381 n374 n284 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00972 n284 b_5 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00971 n381 n376 n284 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00970 n376 b_6 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00969 n284 b_6 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00968 n494 n529 n495 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00967 n495 b_5 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00966 vdd b_5 n492 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00965 n492 n578 n491 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00964 n491 n574 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00963 vdd b_3 n495 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00962 n495 n574 n494 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00961 n494 n578 n495 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00960 n495 b_4 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00959 vdd p_3_2_d2j p_3_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_00958 p_3_1_c2j n492 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00957 vdd n494 p_3_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00956 p_3_2_d2j n584 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00955 n529 b_5 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00954 vdd n529 n493 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00953 n493 b_5 n584 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00952 n574 b_3 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00951 n584 n574 n493 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00950 n493 b_3 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00949 n584 n578 n493 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00948 n578 b_4 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00947 n493 b_4 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00946 n643 n751 n644 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00945 n644 b_3 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00944 vdd b_3 n641 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00943 n641 n758 n640 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00942 n640 n753 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00941 vdd b_1 n644 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00940 n644 n753 n643 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00939 n643 n758 n644 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00938 n644 b_2 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00937 vdd p_2_2_d2j p_2_2_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P 
+ AD=0.7776P PS=5.04U PD=5.04U 
Mtr_00936 n847 n641 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00935 vdd n643 p_2_1_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00934 p_2_2_d2j n755 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00933 n751 b_3 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00932 vdd n751 n695 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00931 n695 b_3 n755 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00930 n753 b_1 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00929 n755 n753 n695 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00928 n695 b_1 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00927 n755 n758 n695 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00926 n758 b_2 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00925 n695 b_2 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00924 n877 b_0 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00923 n946 b_0 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00922 n943 n946 n877 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00921 n877 vss vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00920 n943 n939 n877 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00919 n939 vss vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00918 n877 b_1 n943 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00917 vdd n937 n877 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00916 n937 b_1 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00915 d_0_d2j n943 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00914 vdd n863 d_0_n2j vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00913 p_1_2_c2j n860 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00912 vdd d_0_d2j d_0_d2jbar vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P 
+ PS=5.04U PD=5.04U 
Mtr_00911 n862 b_0 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00910 n863 n946 n862 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00909 n862 n939 n863 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00908 vdd vss n862 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00907 n859 n939 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00906 n860 n946 n859 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00905 vdd b_1 n860 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00904 n862 b_1 vdd vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00903 n863 n937 n862 vdd TP L=0.18U W=2.16U AS=0.7776P AD=0.7776P PS=5.04U 
+ PD=5.04U 
Mtr_00902 c_4_1_sum cla_cell0_0_a n884 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00901 n884 c_4_1_sum cla_cell0_0_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00900 vss n884 p_6 vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P PS=3.96U 
+ PD=3.96U 
Mtr_00899 vss cla_cell0_0_a n881 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00898 n881 c_4_1_sum n880 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00897 vss n880 cla_cell0_0_g vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00896 c_4_2_sum c_4_1_cout n794 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00895 n794 c_4_2_sum c_4_1_cout vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00894 vss n794 cla_cell0_1_p vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00893 vss c_4_1_cout n760 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00892 n760 c_4_2_sum n791 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00891 vss n791 cla_cell0_1_g vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00890 vss n704 cla_cell0_2_g vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00889 n705 c_4_2_cout n704 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00888 vss c_4_3_sum n705 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00887 c_4_2_cout c_4_3_sum n708 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00886 n708 c_4_2_cout c_4_3_sum vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00885 cla_cell0_2_p n708 vss vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00884 vss cla_cell0_2_p cla_cell0_2_pn vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00883 c_4_4_sum c_4_3_cout n594 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00882 n594 c_4_4_sum c_4_3_cout vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00881 vss n594 cla_cell1_3_p1 vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00880 vss c_4_3_cout n540 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00879 n540 c_4_4_sum n651 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00878 vss n651 cla_cell0_3_g vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00877 c_4_4_cout c_4_5_sum n542 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00876 n542 c_4_4_cout c_4_5_sum vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00875 vss n542 cla_cell3_4_p1 vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00874 vss c_4_5_sum n539 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00873 n539 c_4_4_cout n538 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00872 vss n538 cla_cell0_4_g vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00871 vss n431 cla_cell0_5_g vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00870 n320 c_4_6_sum n431 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00869 vss c_4_5_cout n320 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00868 c_4_6_sum c_4_5_cout n433 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00867 n433 c_4_6_sum c_4_5_cout vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00866 cla_cell1_5_p1 n433 vss vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00865 vss cla_cell1_5_p1 cla_cell5_5_p vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00864 vss n318 cla_cell1_6_tsg vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_00863 n319 c_4_6_cout n318 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00862 vss c_4_7_sum n319 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00861 c_4_6_cout c_4_7_sum n321 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00860 n321 c_4_6_cout c_4_7_sum vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00859 cla_cell0_6_p n321 vss vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00858 vss cla_cell0_6_p cla_cell5_6_p vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00857 vss n200 cla_cell0_7_g vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00856 n112 c_4_8_sum n200 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00855 vss c_4_7_cout n112 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00854 c_4_8_sum c_4_7_cout n204 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00853 n204 c_4_8_sum c_4_7_cout vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00852 cla_cell0_7_p n204 vss vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00851 vss cla_cell0_7_p cla_cell0_7_pn vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00850 vss n111 cla_cell0_8_g vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00849 n110 c_4_8_cout n111 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00848 vss cla_cell0_8_a n110 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00847 c_4_8_cout cla_cell0_8_a n114 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00846 n114 c_4_8_cout cla_cell0_8_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00845 cla_cell0_8_p n114 vss vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00844 vss cla_cell0_8_p cla_cell5_8_p vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00843 cla_cell0_8_a cla_cell0_9_a n23 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00842 n23 cla_cell0_8_a cla_cell0_9_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00841 vss n23 cla_cell0_9_p vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00840 vss cla_cell0_9_a n4 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00839 n4 cla_cell0_8_a n18 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00838 vss n18 cla_cell0_9_g vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00837 vss cla_cell0_0_g n759 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00836 n759 cla_cell0_1_p cla_cell1_1_co vss TN L=0.18U W=1.8U AS=0.648P 
+ AD=0.648P PS=4.32U PD=4.32U 
Mtr_00835 cla_cell1_1_co cla_cell0_1_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00834 cla_cell1_2_ng cla_cell0_2_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_00833 vss cla_cell0_2_p cla_cell1_2_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_00832 vss cla_cell0_2_g n536 vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00831 n536 cla_cell1_3_p1 cla_cell1_3_g vss TN L=0.18U W=1.62U AS=0.5832P 
+ AD=0.5832P PS=3.96U PD=3.96U 
Mtr_00830 cla_cell1_3_g cla_cell0_3_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00829 vss cla_cell1_3_p1 n537 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00828 n537 cla_cell0_2_p n592 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00827 n592 cla_cell0_2_p n537 vss TN L=0.18U W=0.18U AS=0.0648P AD=0.0648P 
+ PS=1.08U PD=1.08U 
Mtr_00826 vss cla_cell0_4_g n315 vss TN L=0.18U W=1.62U AS=0.5832P AD=0.5832P 
+ PS=3.96U PD=3.96U 
Mtr_00825 n315 cla_cell1_5_p1 cla_cell2_5_tsg vss TN L=0.18U W=1.62U 
+ AS=0.5832P AD=0.5832P PS=3.96U PD=3.96U 
Mtr_00824 cla_cell2_5_tsg cla_cell0_5_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00823 vss cla_cell1_5_p1 n316 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00822 n316 cla_cell3_4_p1 cla_cell2_5_tsp vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00821 cla_cell2_5_tsp cla_cell3_4_p1 n316 vss TN L=0.18U W=0.18U 
+ AS=0.0648P AD=0.0648P PS=1.08U PD=1.08U 
Mtr_00820 cla_cell1_6_ng cla_cell1_6_tsg vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_00819 vss cla_cell0_6_p cla_cell1_6_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_00818 vss cla_cell1_6_tsg n106 vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00817 n106 cla_cell0_7_p cla_cell1_7_g vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00816 cla_cell1_7_g cla_cell0_7_g vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_00815 n107 cla_cell0_6_p cla_cell2_7_pl vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00814 vss cla_cell0_7_p n107 vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00813 cla_cell1_8_ng cla_cell0_8_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_00812 vss cla_cell0_8_p cla_cell1_8_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_00811 vss cla_cell0_8_g n2 vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00810 n2 cla_cell0_9_p cla_cell1_9_g vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00809 cla_cell1_9_g cla_cell0_9_g vss vss TN L=0.18U W=0.54U AS=0.1944P 
+ AD=0.1944P PS=1.8U PD=1.8U 
Mtr_00808 n3 cla_cell0_8_p n15 vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00807 vss cla_cell0_9_p n3 vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00806 n699 cla_cell1_2_np vss vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00805 n699 cla_cell1_2_ng cla_cell5_2_g vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_00804 vss cla_cell1_1_co n699 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00803 n535 cla_cell1_3_g cla_cell3_4_g2 vss TN L=0.18U W=3.06U AS=1.1016P 
+ AD=1.1016P PS=6.84U PD=6.84U 
Mtr_00802 n535 n592 vss vss TN L=0.18U W=3.06U AS=1.1016P AD=1.1016P PS=6.84U 
+ PD=6.84U 
Mtr_00801 vss cla_cell1_1_co n535 vss TN L=0.18U W=3.06U AS=1.1016P AD=1.1016P 
+ PS=6.84U PD=6.84U 
Mtr_00800 cla_cell2_5_ng cla_cell2_5_tsg vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_00799 vss cla_cell2_5_tsp cla_cell2_5_np vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_00798 vss cla_cell2_5_tsp cla_cell3_6_p1 vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_00797 vss cla_cell1_6_np cla_cell3_6_p1 vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_00796 n310 cla_cell1_6_ng cla_cell2_6_g vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00795 vss cla_cell1_6_np n310 vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00794 n310 cla_cell2_5_tsg vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00793 vss cla_cell2_5_tsp n192 vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_00792 vss cla_cell2_7_pl n192 vss TN L=0.18U W=0.72U AS=0.2592P AD=0.2592P 
+ PS=2.16U PD=2.16U 
Mtr_00791 n163 cla_cell1_7_g cla_cell2_7_g vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00790 vss cla_cell2_7_pl n163 vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00789 n163 cla_cell2_5_tsg vss vss TN L=0.18U W=1.26U AS=0.4536P 
+ AD=0.4536P PS=3.24U PD=3.24U 
Mtr_00788 vss cla_cell3_4_g2 n533 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00787 n533 cla_cell3_4_p1 cla_cell3_4_co vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_00786 cla_cell3_4_co cla_cell0_4_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_00785 vss cla_cell3_4_g2 n308 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00784 n308 cla_cell2_5_np cla_cell3_5_co vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_00783 cla_cell3_5_co cla_cell2_5_ng vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_00782 vss cla_cell3_4_g2 n307 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00781 n307 cla_cell3_6_p1 cla_cell3_6_co vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_00780 cla_cell3_6_co cla_cell2_6_g vss vss TN L=0.18U W=0.72U AS=0.2592P 
+ AD=0.2592P PS=2.16U PD=2.16U 
Mtr_00779 vss cla_cell3_4_g2 n103 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00778 n103 n192 cla_cell3_7_co vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00777 cla_cell3_7_co cla_cell2_7_g vss vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00776 n102 cla_cell1_8_np vss vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00775 n102 cla_cell1_8_ng cla_cell5_8_g vss TN L=0.18U W=1.44U AS=0.5184P 
+ AD=0.5184P PS=3.6U PD=3.6U 
Mtr_00774 vss cla_cell3_7_co n102 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00773 n1 n15 vss vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P PS=3.6U 
+ PD=3.6U 
Mtr_00772 n1 cla_cell1_9_g n14 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00771 vss cla_cell3_7_co n1 vss TN L=0.18U W=1.44U AS=0.5184P AD=0.5184P 
+ PS=3.6U PD=3.6U 
Mtr_00770 n787 cla_cell0_0_g cla_cell0_1_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00769 n787 cla_cell0_1_p cla_cell0_0_g vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00768 p_7 n787 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_00767 n697 cla_cell0_2_pn cla_cell1_1_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00766 n697 cla_cell1_1_co cla_cell0_2_pn vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00765 p_8 n697 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_00764 n645 cla_cell5_2_g cla_cell1_3_p1 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00763 n645 cla_cell1_3_p1 cla_cell5_2_g vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00762 p_9 n645 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_00761 n531 cla_cell3_4_p1 cla_cell3_4_g2 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00760 n531 cla_cell3_4_g2 cla_cell3_4_p1 vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00759 p_10 n531 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_00758 n421 cla_cell3_4_co cla_cell5_5_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00757 n421 cla_cell5_5_p cla_cell3_4_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00756 p_11 n421 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_00755 n304 cla_cell5_6_p cla_cell3_5_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00754 n304 cla_cell3_5_co cla_cell5_6_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00753 p_12 n304 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_00752 n190 cla_cell3_6_co cla_cell0_7_pn vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00751 n190 cla_cell0_7_pn cla_cell3_6_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00750 p_13 n190 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_00749 n101 cla_cell5_8_p cla_cell3_7_co vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00748 n101 cla_cell3_7_co cla_cell5_8_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00747 p_14 n101 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_00746 n11 cla_cell5_8_g cla_cell0_9_p vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00745 n11 cla_cell0_9_p cla_cell5_8_g vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00744 p_15 n11 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P PS=7.92U 
+ PD=7.92U 
Mtr_00743 vss n35 cla_cell0_9_a vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00742 n5 p_4_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00741 vss c_4_7_a n5 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00740 n35 c_4_8_cin n5 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00739 n6 p_4_9_pi2j n35 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00738 vss c_4_7_a n6 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00737 n30 c_4_8_cin n26 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00736 n26 n30 c_4_8_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00735 c_4_7_a p_4_9_pi2j n32 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00734 n32 c_4_7_a p_4_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00733 cla_cell0_8_a n26 vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00732 vss n32 n30 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P PS=6.48U 
+ PD=6.48U 
Mtr_00731 n40 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00730 n39 a_7 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00729 vss p_4_9_t_s p_4_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00728 p_4_9_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00727 n39 n40 p_4_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00726 p_4_9_t_s n39 n40 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00725 n128 p_4_2_d2j n127 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00724 n129 p_4_2_d2jbar n128 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00723 p_4_8_t_s n128 n126 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00722 n128 n126 p_4_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00721 p_4_8_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00720 vss p_4_8_t_s p_4_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00719 n126 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00718 vss a_7 n129 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00717 n127 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00716 vss n120 c_4_8_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00715 n121 c_4_7_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00714 vss p_4_8_pi2j n121 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00713 n120 c_4_8_cin n121 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00712 n119 c_4_7_a n120 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00711 vss p_4_8_pi2j n119 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00710 n116 c_4_8_cin c_4_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00709 c_4_8_s2_s n116 c_4_8_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00708 p_4_8_pi2j c_4_7_a c_4_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00707 c_4_8_s1_s p_4_8_pi2j c_4_7_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00706 c_4_8_sum c_4_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00705 vss c_4_8_s1_s n116 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00704 vss n221 c_4_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00703 n164 p_4_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00702 vss c_4_7_a n164 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00701 n221 c_4_7_cin n164 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00700 n118 p_4_7_pi2j n221 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00699 vss c_4_7_a n118 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00698 n216 c_4_7_cin c_4_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00697 c_4_7_s2_s n216 c_4_7_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00696 c_4_7_a p_4_7_pi2j c_4_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00695 c_4_7_s1_s c_4_7_a p_4_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00694 c_4_7_sum c_4_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00693 vss c_4_7_s1_s n216 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00692 n227 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00691 vss a_5 n168 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00690 n168 p_4_2_d2j n222 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00689 n222 p_4_2_d2jbar n167 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00688 n167 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00687 vss p_4_7_t_s p_4_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00686 p_4_7_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00685 n222 n227 p_4_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00684 p_4_7_t_s n222 n227 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00683 n333 p_4_2_d2j n292 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00682 n293 p_4_2_d2jbar n333 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00681 p_4_6_t_s n333 n335 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00680 n333 n335 p_4_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00679 p_4_6_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00678 vss p_4_6_t_s p_4_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00677 n335 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00676 vss a_5 n293 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00675 n292 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00674 vss n329 c_4_6_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00673 n324 c_4_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00672 vss p_4_6_pi2j n324 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00671 n329 c_4_6_cin n324 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00670 n328 c_4_6_a n329 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00669 vss p_4_6_pi2j n328 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00668 n291 c_4_6_cin c_4_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00667 c_4_6_s2_s n291 c_4_6_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00666 p_4_6_pi2j c_4_6_a c_4_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00665 c_4_6_s1_s p_4_6_pi2j c_4_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00664 c_4_6_sum c_4_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00663 vss c_4_6_s1_s n291 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00662 vss n446 c_4_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00661 n389 c_4_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00660 vss c_4_5_a n389 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00659 n446 c_4_5_cin n389 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00658 n327 c_4_5_b n446 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00657 vss c_4_5_a n327 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00656 n393 c_4_5_cin c_4_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00655 c_4_5_s2_s n393 c_4_5_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00654 c_4_5_a c_4_5_b c_4_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00653 c_4_5_s1_s c_4_5_a c_4_5_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00652 c_4_5_sum c_4_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00651 vss c_4_5_s1_s n393 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00650 n450 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00649 vss a_3 n337 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00648 n337 p_4_2_d2j n447 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00647 n447 p_4_2_d2jbar n336 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00646 n336 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00645 vss p_4_5_t_s c_4_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00644 c_4_5_b p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00643 n447 n450 p_4_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00642 p_4_5_t_s n447 n450 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00641 n508 p_4_2_d2j n506 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00640 n507 p_4_2_d2jbar n508 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00639 p_4_4_t_s n508 n505 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00638 n508 n505 p_4_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00637 p_4_4_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00636 vss p_4_4_t_s p_4_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00635 n505 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00634 vss a_3 n507 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00633 n506 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00632 vss n499 c_4_4_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00631 n544 c_4_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00630 vss p_4_4_pi2j n544 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00629 n499 c_4_4_cin n544 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00628 n548 c_4_4_a n499 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00627 vss p_4_4_pi2j n548 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00626 n502 c_4_4_cin c_4_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00625 c_4_4_s2_s n502 c_4_4_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00624 p_4_4_pi2j c_4_4_a c_4_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00623 c_4_4_s1_s p_4_4_pi2j c_4_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00622 c_4_4_sum c_4_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00621 vss c_4_4_s1_s n502 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00620 vss n600 c_4_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00619 n547 c_4_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00618 vss c_4_3_a n547 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00617 n600 c_4_3_cin n547 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00616 n546 c_4_3_b n600 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00615 vss c_4_3_a n546 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00614 n603 c_4_3_cin c_4_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00613 c_4_3_s2_s n603 c_4_3_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00612 c_4_3_a c_4_3_b c_4_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00611 c_4_3_s1_s c_4_3_a c_4_3_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00610 c_4_3_sum c_4_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00609 vss c_4_3_s1_s n603 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00608 n608 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00607 vss a_1 n552 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00606 n552 p_4_2_d2j n605 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00605 n605 p_4_2_d2jbar n551 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00604 n551 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00603 vss p_4_3_t_s c_4_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00602 c_4_3_b p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00601 n605 n608 p_4_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00600 p_4_3_t_s n605 n608 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00599 n721 p_4_2_d2j n719 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00598 n720 p_4_2_d2jbar n721 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00597 p_4_2_t_s n721 n718 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00596 n721 n718 p_4_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00595 c_4_2_b p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00594 vss p_4_2_t_s c_4_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00593 n718 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00592 vss a_1 n720 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00591 n719 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00590 vss n712 c_4_2_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00589 n711 c_4_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00588 vss c_4_2_b n711 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00587 n712 c_4_2_cin n711 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00586 n710 c_4_2_a n712 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00585 vss c_4_2_b n710 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00584 n714 c_4_2_cin c_4_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00583 c_4_2_s2_s n714 c_4_2_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00582 c_4_2_b c_4_2_a c_4_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00581 c_4_2_s1_s c_4_2_b c_4_2_a vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00580 c_4_2_sum c_4_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00579 vss c_4_2_s1_s n714 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00578 vss n805 c_4_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00577 n763 p_4_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00576 vss c_4_1_a n763 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00575 n805 c_4_1_cin n763 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00574 n762 p_4_1_pi2j n805 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00573 vss c_4_1_a n762 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00572 n804 c_4_1_cin c_4_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00571 c_4_1_s2_s n804 c_4_1_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00570 c_4_1_a p_4_1_pi2j c_4_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00569 c_4_1_s1_s c_4_1_a p_4_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00568 c_4_1_sum c_4_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00567 vss c_4_1_s1_s n804 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00566 n814 p_4_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00565 n815 p_4_2_d2jbar n766 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00564 n766 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00563 vss p_4_1_t_s p_4_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00562 p_4_1_pi2j p_4_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00561 n815 n814 p_4_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00560 p_4_1_t_s n815 n814 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00559 cl4_4_s1_s n908 c_3_1_sum vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00558 n908 c_3_1_sum cl4_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00557 vss cl4_4_s1_s p_4 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00556 vss c_3_1_sum n898 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00555 n898 n908 n897 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00554 n896 n897 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00553 n894 c_3_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00552 vss c_3_2_sum n894 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00551 n895 c_3_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00550 n893 c_3_1_cout n895 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00549 n890 c_3_1_sum n893 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00548 n894 n908 n890 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00547 cla_cell0_0_a n893 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00546 cl4_4_s2_s c_3_1_cout c_3_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00545 c_3_1_cout c_3_2_sum cl4_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00544 vss cl4_4_s2_s n888 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00543 cl4_4_s3_s n888 n896 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00542 n888 n896 cl4_4_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00541 vss cl4_4_s3_s p_5 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00540 vss c_3_9_s1_s n51 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00539 c_4_7_a c_3_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00538 c_3_9_s1_s c_3_7_a p_3_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00537 c_3_7_a p_3_9_pi2j c_3_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00536 c_3_9_s2_s n51 c_3_8_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00535 n51 c_3_8_cin c_3_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00534 vss c_3_7_a n7 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00533 n7 p_3_9_pi2j n42 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00532 n42 c_3_8_cin n8 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00531 vss c_3_7_a n8 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00530 n8 p_3_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00529 vss n42 c_4_8_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00528 n53 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00527 n56 a_7 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00526 vss p_3_9_t_s p_3_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00525 p_3_9_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00524 n56 n53 p_3_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00523 p_3_9_t_s n56 n53 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00522 n143 p_3_2_d2j n142 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00521 n140 p_3_2_d2jbar n143 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00520 p_3_8_t_s n143 n141 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00519 n143 n141 p_3_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00518 p_3_8_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00517 vss p_3_8_t_s p_3_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00516 n141 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00515 vss a_7 n140 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00514 n142 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00513 vss c_3_8_s1_s n134 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00512 c_4_6_a c_3_8_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00511 c_3_8_s1_s p_3_8_pi2j c_3_7_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00510 c_3_8_s2_s n134 c_3_8_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00509 n134 c_3_8_cin c_3_8_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00508 vss p_3_8_pi2j n131 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00507 n131 c_3_7_a n132 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00506 n132 c_3_8_cin n133 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00505 vss p_3_8_pi2j n133 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00504 n133 c_3_7_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00503 vss n132 c_4_7_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00502 p_3_8_pi2j c_3_7_a c_3_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00501 vss n234 c_4_6_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00500 n169 p_3_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00499 vss c_3_7_a n169 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00498 n234 c_3_7_cin n169 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00497 n130 p_3_7_pi2j n234 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00496 vss c_3_7_a n130 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00495 n243 c_3_7_cin c_3_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00494 c_3_7_s2_s n243 c_3_7_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00493 c_3_7_a p_3_7_pi2j c_3_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00492 c_3_7_s1_s c_3_7_a p_3_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00491 c_4_5_a c_3_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00490 vss c_3_7_s1_s n243 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00489 n246 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00488 vss a_5 n172 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00487 n172 p_3_2_d2j n245 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00486 n245 p_3_2_d2jbar n173 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00485 n173 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00484 vss p_3_7_t_s p_3_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00483 p_3_7_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00482 n245 n246 p_3_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00481 p_3_7_t_s n245 n246 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00480 n347 p_3_2_d2j n298 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00479 n297 p_3_2_d2jbar n347 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00478 p_3_6_t_s n347 n348 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00477 n347 n348 p_3_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00476 p_3_6_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00475 vss p_3_6_t_s p_3_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00474 n348 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00473 vss a_5 n297 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00472 n298 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00471 vss c_3_6_s1_s n296 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00470 c_4_4_a c_3_6_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00469 c_3_6_s1_s p_3_6_pi2j c_3_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00468 c_3_6_s2_s n296 c_2_7_cout vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00467 n296 c_2_7_cout c_3_6_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00466 vss p_3_6_pi2j n340 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00465 n340 c_3_6_a n341 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00464 n341 c_2_7_cout n339 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00463 vss p_3_6_pi2j n339 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00462 n339 c_3_6_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00461 vss n341 c_4_5_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00460 p_3_6_pi2j c_3_6_a c_3_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00459 vss n456 c_4_4_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00458 n397 c_3_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00457 vss c_3_5_a n397 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00456 n456 c_3_5_cin n397 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00455 n338 c_3_5_b n456 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00454 vss c_3_5_a n338 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00453 n402 c_3_5_cin c_3_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00452 c_3_5_s2_s n402 c_3_5_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00451 c_3_5_a c_3_5_b c_3_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00450 c_3_5_s1_s c_3_5_a c_3_5_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00449 c_4_3_a c_3_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00448 vss c_3_5_s1_s n402 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00447 n465 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00446 vss a_3 n350 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00445 n350 p_3_2_d2j n466 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00444 n466 p_3_2_d2jbar n351 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00443 n351 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00442 vss p_3_5_t_s c_3_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00441 c_3_5_b p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00440 n466 n465 p_3_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00439 p_3_5_t_s n466 n465 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00438 n517 p_3_2_d2j n518 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00437 n516 p_3_2_d2jbar n517 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00436 p_3_4_t_s n517 n515 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00435 n517 n515 p_3_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00434 p_3_4_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00433 vss p_3_4_t_s p_3_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00432 n515 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00431 vss a_3 n516 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00430 n518 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00429 vss c_3_4_s1_s n514 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00428 c_4_2_a c_3_4_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00427 c_3_4_s1_s p_3_4_pi2j c_3_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00426 c_3_4_s2_s n514 c_2_5_cout vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00425 n514 c_2_5_cout c_3_4_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00424 vss p_3_4_pi2j n555 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00423 n555 c_3_4_a n509 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00422 n509 c_2_5_cout n556 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00421 vss p_3_4_pi2j n556 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00420 n556 c_3_4_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00419 vss n509 c_4_3_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00418 p_3_4_pi2j c_3_4_a c_3_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00417 vss n610 c_4_2_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00416 n554 c_3_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00415 vss c_3_3_a n554 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00414 n610 c_3_3_cin n554 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00413 n553 c_3_3_b n610 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00412 vss c_3_3_a n553 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00411 n616 c_3_3_cin c_3_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00410 c_3_3_s2_s n616 c_3_3_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00409 c_3_3_a c_3_3_b c_3_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00408 c_3_3_s1_s c_3_3_a c_3_3_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00407 c_4_1_a c_3_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00406 vss c_3_3_s1_s n616 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00405 n617 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00404 vss a_1 n560 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00403 n560 p_3_2_d2j n619 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00402 n619 p_3_2_d2jbar n561 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00401 n561 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00400 vss p_3_3_t_s c_3_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00399 c_3_3_b p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00398 n619 n617 p_3_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00397 p_3_3_t_s n619 n617 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00396 n733 p_3_2_d2j n734 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00395 n732 p_3_2_d2jbar n733 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00394 p_3_2_t_s n733 n731 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00393 n733 n731 p_3_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00392 c_3_2_b p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00391 vss p_3_2_t_s c_3_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00390 n731 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00389 vss a_1 n732 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00388 n734 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00387 vss c_3_2_s1_s n727 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00386 c_3_2_sum c_3_2_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00385 c_3_2_s1_s c_3_2_b c_3_2_a vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00384 c_3_2_s2_s n727 c_2_3_cout vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00383 n727 c_2_3_cout c_3_2_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00382 vss c_3_2_b n723 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00381 n723 c_3_2_a n724 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00380 n724 c_2_3_cout n722 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00379 vss c_3_2_b n722 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00378 n722 c_3_2_a vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00377 vss n724 c_4_1_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00376 c_3_2_b c_3_2_a c_3_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00375 vss n819 c_3_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00374 n768 p_3_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00373 vss c_3_1_a n768 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00372 n819 c_3_1_cin n768 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00371 n767 p_3_1_pi2j n819 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00370 vss c_3_1_a n767 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00369 n826 c_3_1_cin c_3_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00368 c_3_1_s2_s n826 c_3_1_cin vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00367 c_3_1_a p_3_1_pi2j c_3_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00366 c_3_1_s1_s c_3_1_a p_3_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00365 c_3_1_sum c_3_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00364 vss c_3_1_s1_s n826 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00363 n830 p_3_1_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00362 n834 p_3_2_d2jbar n771 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00361 n771 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00360 vss p_3_1_t_s p_3_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00359 p_3_1_pi2j p_3_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00358 n834 n830 p_3_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00357 p_3_1_t_s n834 n830 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00356 cl4_3_s1_s n922 c_2_1_sum vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00355 n922 c_2_1_sum cl4_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00354 vss cl4_3_s1_s p_2 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00353 vss c_2_1_sum n915 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00352 n915 n922 n913 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00351 n914 n913 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00350 n912 c_2_1_cout vss vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00349 vss c_2_2_sum n912 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00348 n909 c_2_2_sum vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00347 n910 c_2_1_cout n909 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00346 n907 c_2_1_sum n910 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00345 n912 n922 n907 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00344 n908 n910 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00343 cl4_3_s2_s c_2_1_cout c_2_2_sum vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00342 c_2_1_cout c_2_2_sum cl4_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00341 vss cl4_3_s2_s n906 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00340 cl4_3_s3_s n906 n914 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00339 n906 n914 cl4_3_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00338 vss cl4_3_s3_s p_3 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00337 vss n60 c_3_8_cin vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00336 n10 p_2_9_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00335 vss c_2_7_a n10 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00334 n60 vss n10 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00333 n9 p_2_9_pi2j n60 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00332 vss c_2_7_a n9 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00331 n64 vss c_2_9_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00330 c_2_9_s2_s n64 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00329 c_2_7_a p_2_9_pi2j c_2_9_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00328 c_2_9_s1_s c_2_7_a p_2_9_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00327 c_3_7_a c_2_9_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00326 vss c_2_9_s1_s n64 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00325 n68 n847 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00324 n72 a_7 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00323 vss p_2_9_t_s p_2_9_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00322 p_2_9_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00321 n72 n68 p_2_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00320 p_2_9_t_s n72 n68 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00319 n153 p_2_2_d2j n151 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00318 n152 p_2_2_d2jbar n153 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00317 p_2_8_t_s n153 n150 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00316 n153 n150 p_2_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00315 p_2_8_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00314 vss p_2_8_t_s p_2_8_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00313 n150 n847 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00312 vss a_7 n152 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00311 n151 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00310 c_3_7_cin n146 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00309 vss c_2_7_a n145 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00308 n145 p_2_8_pi2j n146 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00307 p_2_8_pi2j c_2_7_a c_2_8_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00306 c_2_8_s1_s p_2_8_pi2j c_2_7_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00305 c_3_6_a c_2_8_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00304 vss n253 c_2_7_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00303 n174 p_2_7_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00302 vss c_2_7_a n174 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00301 n253 vss n174 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00300 n144 p_2_7_pi2j n253 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00299 vss c_2_7_a n144 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00298 n261 vss c_2_7_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00297 c_2_7_s2_s n261 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00296 c_2_7_a p_2_7_pi2j c_2_7_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00295 c_2_7_s1_s c_2_7_a p_2_7_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00294 c_3_5_a c_2_7_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00293 vss c_2_7_s1_s n261 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00292 n266 n847 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00291 vss a_5 n178 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00290 n178 p_2_2_d2j n265 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00289 n265 p_2_2_d2jbar n177 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00288 n177 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00287 vss p_2_7_t_s p_2_7_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00286 p_2_7_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00285 n265 n266 p_2_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00284 p_2_7_t_s n265 n266 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00283 n359 p_2_2_d2j n300 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00282 n299 p_2_2_d2jbar n359 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00281 p_2_6_t_s n359 n360 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00280 n359 n360 p_2_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00279 p_2_6_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00278 vss p_2_6_t_s p_2_6_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00277 n360 n847 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00276 vss a_5 n299 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00275 n300 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00274 c_3_5_cin n354 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00273 vss c_2_6_a n353 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00272 n353 p_2_6_pi2j n354 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00271 p_2_6_pi2j c_2_6_a c_2_6_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00270 c_2_6_s1_s p_2_6_pi2j c_2_6_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00269 c_3_4_a c_2_6_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00268 vss n472 c_2_5_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00267 n406 c_2_5_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00266 vss c_2_5_a n406 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00265 n472 p_4_1_c2j n406 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00264 n352 c_2_5_b n472 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00263 vss c_2_5_a n352 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00262 n409 p_4_1_c2j c_2_5_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00261 c_2_5_s2_s n409 p_4_1_c2j vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00260 c_2_5_a c_2_5_b c_2_5_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00259 c_2_5_s1_s c_2_5_a c_2_5_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00258 c_3_3_a c_2_5_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00257 vss c_2_5_s1_s n409 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00256 n480 n847 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00255 vss a_3 n362 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00254 n362 p_2_2_d2j n479 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00253 n479 p_2_2_d2jbar n361 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00252 n361 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00251 vss p_2_5_t_s c_2_5_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00250 c_2_5_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00249 n479 n480 p_2_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00248 p_2_5_t_s n479 n480 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00247 n523 p_2_2_d2j n522 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00246 n521 p_2_2_d2jbar n523 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00245 p_2_4_t_s n523 n520 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00244 n523 n520 p_2_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00243 p_2_4_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00242 vss p_2_4_t_s p_2_4_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00241 n520 n847 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00240 vss a_3 n521 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00239 n522 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00238 c_3_3_cin n562 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00237 vss c_2_4_a n519 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00236 n519 p_2_4_pi2j n562 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00235 p_2_4_pi2j c_2_4_a c_2_4_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00234 c_2_4_s1_s p_2_4_pi2j c_2_4_a vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00233 c_3_2_a c_2_4_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00232 vss n623 c_2_3_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00231 n565 c_2_3_b vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00230 vss c_2_3_a n565 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00229 n623 p_3_1_c2j n565 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00228 n564 c_2_3_b n623 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00227 vss c_2_3_a n564 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00226 n627 p_3_1_c2j c_2_3_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00225 c_2_3_s2_s n627 p_3_1_c2j vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00224 c_2_3_a c_2_3_b c_2_3_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00223 c_2_3_s1_s c_2_3_a c_2_3_b vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00222 c_3_1_a c_2_3_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00221 vss c_2_3_s1_s n627 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00220 n630 n847 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00219 vss a_1 n569 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00218 n569 p_2_2_d2j n634 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00217 n634 p_2_2_d2jbar n570 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00216 n570 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00215 vss p_2_3_t_s c_2_3_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00214 c_2_3_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00213 n634 n630 p_2_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00212 p_2_3_t_s n634 n630 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00211 n743 p_2_2_d2j n742 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00210 n741 p_2_2_d2jbar n743 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00209 p_2_2_t_s n743 n739 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00208 n743 n739 p_2_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00207 c_2_2_b p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00206 vss p_2_2_t_s c_2_2_b vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00205 n739 n847 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00204 vss a_1 n741 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00203 n742 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00202 c_3_1_cin n736 vss vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00201 vss c_2_2_a n735 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00200 n735 c_2_2_b n736 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00199 c_2_2_b c_2_2_a c_2_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00198 c_2_2_s1_s c_2_2_b c_2_2_a vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00197 c_2_2_sum c_2_2_s1_s vss vss TN L=0.18U W=2.88U AS=1.0368P 
+ AD=1.0368P PS=6.48U PD=6.48U 
Mtr_00196 vss n836 c_2_1_cout vss TN L=0.18U W=1.26U AS=0.4536P AD=0.4536P 
+ PS=3.24U PD=3.24U 
Mtr_00195 n773 p_2_1_pi2j vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00194 vss c_2_1_a n773 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00193 n836 n847 n773 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00192 n772 p_2_1_pi2j n836 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00191 vss c_2_1_a n772 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00190 n844 n847 c_2_1_s2_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00189 c_2_1_s2_s n844 n847 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00188 c_2_1_a p_2_1_pi2j c_2_1_s1_s vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00187 c_2_1_s1_s c_2_1_a p_2_1_pi2j vss TN L=0.18U W=0.9U AS=0.324P 
+ AD=0.324P PS=2.52U PD=2.52U 
Mtr_00186 c_2_1_sum c_2_1_s2_s vss vss TN L=0.18U W=3.6U AS=1.296P AD=1.296P 
+ PS=7.92U PD=7.92U 
Mtr_00185 vss c_2_1_s1_s n844 vss TN L=0.18U W=2.88U AS=1.0368P AD=1.0368P 
+ PS=6.48U PD=6.48U 
Mtr_00184 p_2_1_t_s n853 n849 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00183 n853 n849 p_2_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00182 p_2_1_pi2j p_2_1_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00181 vss p_2_1_t_s p_2_1_pi2j vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00180 n776 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00179 n853 p_2_2_d2jbar n776 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00178 n849 n847 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00177 cl4_2_s1_s p_1_2_c2j n932 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00176 p_1_2_c2j n932 cl4_2_s1_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00175 vss cl4_2_s1_s p_0 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00174 vss n932 n928 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00173 n928 p_1_2_c2j n926 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00172 n927 n926 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00171 vss p_1_2_pi2j n925 vss TN L=0.18U W=1.8U AS=0.648P AD=0.648P 
+ PS=4.32U PD=4.32U 
Mtr_00170 n924 n932 n923 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00169 n925 p_1_2_c2j n924 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00168 n922 n923 vss vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P PS=2.52U 
+ PD=2.52U 
Mtr_00167 cl4_2_s3_s p_1_2_pi2j n927 vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00166 p_1_2_pi2j n927 cl4_2_s3_s vss TN L=0.18U W=0.9U AS=0.324P AD=0.324P 
+ PS=2.52U PD=2.52U 
Mtr_00165 vss cl4_2_s3_s p_1 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00164 vss p_1_9_t_s c_2_7_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00163 c_2_7_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00162 p_1_9_a n76 p_1_9_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00161 p_1_9_t_s p_1_9_a n76 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00160 n76 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00159 p_1_9_a a_7 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00158 vss d_0_n2j c_2_6_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00157 p_1_8_t_s n155 n157 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00156 vss a_7 n158 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00155 n155 d_0_d2j n156 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00154 n156 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00153 c_2_6_a p_1_8_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00152 n155 n157 p_1_8_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00151 n157 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00150 n158 d_0_d2jbar n155 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00149 p_1_7_a d_0_d2jbar n181 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00148 n182 d_0_d2j p_1_7_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00147 vss a_5 n182 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00146 n273 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00145 p_1_7_t_s p_1_7_a n273 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00144 p_1_7_a n273 p_1_7_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00143 c_2_5_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00142 vss p_1_7_t_s c_2_5_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00141 n181 a_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00140 vss d_0_n2j c_2_4_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00139 p_1_6_t_s n363 n365 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00138 vss a_5 n301 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00137 n363 d_0_d2j n302 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00136 n302 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00135 c_2_4_a p_1_6_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00134 n363 n365 p_1_6_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00133 n365 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00132 n301 d_0_d2jbar n363 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00131 p_1_5_a d_0_d2jbar n367 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00130 n368 d_0_d2j p_1_5_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00129 vss a_3 n368 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00128 n486 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00127 p_1_5_t_s p_1_5_a n486 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00126 p_1_5_a n486 p_1_5_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00125 c_2_3_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00124 vss p_1_5_t_s c_2_3_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00123 n367 a_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00122 vss d_0_n2j c_2_2_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00121 p_1_4_t_s n527 n524 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00120 vss a_3 n525 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00119 n527 d_0_d2j n526 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00118 n526 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00117 c_2_2_a p_1_4_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00116 n527 n524 p_1_4_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00115 n524 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00114 n525 d_0_d2jbar n527 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00113 p_1_3_a d_0_d2jbar n572 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00112 n573 d_0_d2j p_1_3_a vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00111 vss a_1 n573 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00110 n690 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00109 p_1_3_t_s p_1_3_a n690 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00108 p_1_3_a n690 p_1_3_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00107 c_2_1_a d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00106 vss p_1_3_t_s c_2_1_a vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00105 n572 a_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00104 vss d_0_n2j p_1_2_pi2j vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00103 p_1_2_t_s n748 n745 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00102 vss a_1 n746 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00101 n748 d_0_d2j n747 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00100 n747 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00099 p_1_2_pi2j p_1_2_t_s vss vss TN L=0.18U W=2.52U AS=0.9072P 
+ AD=0.9072P PS=5.76U PD=5.76U 
Mtr_00098 n748 n745 p_1_2_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00097 n745 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00096 n746 d_0_d2jbar n748 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00095 n777 a_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00094 vss p_1_1_t_s n932 vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00093 n932 d_0_n2j vss vss TN L=0.18U W=2.52U AS=0.9072P AD=0.9072P 
+ PS=5.76U PD=5.76U 
Mtr_00092 n857 n856 p_1_1_t_s vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00091 p_1_1_t_s n857 n856 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00090 n856 p_1_2_c2j vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00089 n857 d_0_d2jbar n777 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00088 vss n285 p_4_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00087 p_4_1_c2j n283 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00086 vss n374 n159 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00085 n159 n376 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00084 n283 b_7 n159 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00083 vss n369 n186 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00082 n186 n376 n185 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00081 n185 n374 n285 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00080 n285 b_5 n183 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00079 n183 b_6 n184 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00078 n184 b_7 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00077 p_4_2_d2j n381 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00076 vss p_4_2_d2j p_4_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00075 n372 n369 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00074 n369 b_7 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00073 vss b_7 n373 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00072 n373 n374 n382 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00071 n374 b_5 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00070 n372 b_5 n383 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00069 n376 b_6 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00068 n382 n376 n381 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00067 n381 b_6 n383 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00066 vss n494 p_3_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00065 p_3_1_c2j n492 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00064 vss n574 n371 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00063 n371 n578 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00062 n492 b_5 n371 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00061 vss n529 n379 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00060 n379 n578 n380 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00059 n380 n574 n494 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00058 n494 b_3 n378 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00057 n378 b_4 n377 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00056 n377 b_5 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00055 p_3_2_d2j n584 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00054 vss p_3_2_d2j p_3_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00053 n576 n529 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00052 n529 b_5 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00051 vss b_5 n577 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00050 n577 n574 n585 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00049 n574 b_3 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00048 n576 b_3 n586 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00047 n578 b_4 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00046 n585 n578 n584 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00045 n584 b_4 n586 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00044 vss n643 p_2_1_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00043 n847 n641 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00042 vss n753 n575 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00041 n575 n758 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00040 n641 b_3 n575 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00039 vss n751 n582 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00038 n582 n758 n583 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00037 n583 n753 n643 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00036 n643 b_1 n581 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00035 n581 b_2 n580 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00034 n580 b_3 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00033 p_2_2_d2j n755 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00032 vss p_2_2_d2j p_2_2_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P 
+ AD=0.3888P PS=2.88U PD=2.88U 
Mtr_00031 n778 n751 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00030 n751 b_3 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00029 vss b_3 n750 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00028 n750 n753 n756 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00027 n753 b_1 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00026 n778 b_1 n757 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00025 n758 b_2 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00024 n756 n758 n755 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00023 n755 b_2 n757 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00022 n943 b_0 n942 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00021 n944 n946 n943 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00020 n946 b_0 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00019 n938 vss n942 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00018 n939 vss vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00017 n940 n939 n944 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00016 vss b_1 n940 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00015 n937 b_1 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00014 n938 n937 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00013 vss d_0_d2j d_0_d2jbar vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00012 d_0_d2j n943 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00011 n782 b_1 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00010 n783 b_0 n782 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00009 n863 vss n783 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00008 n780 n939 n863 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00007 n781 n946 n780 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00006 vss n937 n781 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00005 n860 b_1 n779 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00004 n779 n946 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00003 vss n939 n779 vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P PS=2.88U 
+ PD=2.88U 
Mtr_00002 p_1_2_c2j n860 vss vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
Mtr_00001 vss n863 d_0_n2j vss TN L=0.18U W=1.08U AS=0.3888P AD=0.3888P 
+ PS=2.88U PD=2.88U 
.ends ex_m8x8

