
.subckt addaccu vss vdd sel s_3 s_2 s_1 s_0 ck b_3 b_2 
+ b_1 b_0 a_3 a_2 a_1 a_0 
M1 vdd n5912_96 s_2_24 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M2 s_2_24 n5912_99 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M3 vdd n5912_100 s_2_21 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M4 s_2_21 n5912_101 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M5 vdd n5912_81 s_2_19 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M6 s_2_19 n5912_84 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M7 vdd n5912_85 s_2_17 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M8 s_2_17 n5912_86 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M9 vdd n5912_66 s_2_15 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M10 s_2_15 n5912_69 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M11 vdd n5912_70 s_2_13 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M12 s_2_13 n5912_71 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M13 vdd n5912_51 s_2_11 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M14 s_2_11 n5912_54 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M15 vdd n5912_55 s_2_9 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M16 s_2_9 n5912_56 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M17 vdd n5912_16 s_2_7 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M18 s_2_7 n5912_19 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M19 vdd n5912_20 s_2_5 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M20 s_2_5 n5912_21 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M21 vdd n5912_1 s_2_3 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M22 s_2_3 n5912_4 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M23 vdd n5912_5 s_2_1 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M24 s_2_1 n5912_6 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M25 vdd n5373_3 n5912_50 vdd TP L=0.18U W=10.872U AS=3.91392P AD=3.91392P 
+ PS=22.464U PD=22.464U 
M26 n5912_50 n5373_4 vdd vdd TP L=0.18U W=10.872U AS=3.91392P AD=3.91392P 
+ PS=22.464U PD=22.464U 
M27 n5912_31 n5373_6 vdd vdd TP L=0.18U W=10.872U AS=3.91392P AD=3.91392P 
+ PS=22.464U PD=22.464U 
M28 vdd n5334_4 n5373_2 vdd TP L=0.18U W=10.872U AS=3.91392P AD=3.91392P 
+ PS=22.464U PD=22.464U 
M29 vdd n5373_5 n5912_31 vdd TP L=0.18U W=10.872U AS=3.91392P AD=3.91392P 
+ PS=22.464U PD=22.464U 
M30 n5334_2 ss_2_1 vdd vdd TP L=0.18U W=10.872U AS=3.91392P AD=3.91392P 
+ PS=22.464U PD=22.464U 
M31 vdd n5111_96 s_3_24 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M32 s_3_24 n5111_99 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M33 vdd n5111_100 s_3_21 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M34 s_3_21 n5111_101 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M35 vdd n5111_81 s_3_19 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M36 s_3_19 n5111_84 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M37 vdd n5111_85 s_3_17 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M38 s_3_17 n5111_86 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M39 vdd n5111_66 s_3_15 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M40 s_3_15 n5111_69 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M41 vdd n5111_70 s_3_13 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M42 s_3_13 n5111_71 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M43 vdd n5111_51 s_3_11 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M44 s_3_11 n5111_54 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M45 vdd n5111_55 s_3_9 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M46 s_3_9 n5111_56 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M47 vdd n5111_16 s_3_7 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M48 s_3_7 n5111_19 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M49 vdd n5111_20 s_3_5 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M50 s_3_5 n5111_21 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M51 vdd n5111_1 s_3_3 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M52 s_3_3 n5111_4 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M53 vdd n5111_5 s_3_1 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M54 s_3_1 n5111_6 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M55 vdd n4572_3 n5111_50 vdd TP L=0.18U W=10.872U AS=3.91392P 
+ AD=3.91392P PS=22.464U PD=22.464U 
M56 n5111_50 n4572_4 vdd vdd TP L=0.18U W=10.872U AS=3.91392P 
+ AD=3.91392P PS=22.464U PD=22.464U 
M57 n5111_31 n4572_6 vdd vdd TP L=0.18U W=10.872U AS=3.91392P 
+ AD=3.91392P PS=22.464U PD=22.464U 
M58 vdd n4533_4 n4572_2 vdd TP L=0.18U W=10.872U AS=3.91392P AD=3.91392P 
+ PS=22.464U PD=22.464U 
M59 vdd n4572_5 n5111_31 vdd TP L=0.18U W=10.872U AS=3.91392P 
+ AD=3.91392P PS=22.464U PD=22.464U 
M60 n4533_2 ss_3_3 vdd vdd TP L=0.18U W=10.872U AS=3.91392P AD=3.91392P 
+ PS=22.464U PD=22.464U 
M61 sel_1 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M62 vdd vdd sel_1 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M63 sel_3 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M64 vdd vdd sel_3 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M65 vdd sel_10 n2124_10 vdd TP L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M66 selsel_67 n2124_8 vdd vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M67 vdd n2124_7 selsel_67 vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M68 vdd vdd ck_3 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M69 ck_3 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M70 vdd vdd ck_1 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M71 ck_1 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M72 p17_logic_ck_60 n1874_19 vdd vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M73 vdd n1874_20 p17_logic_ck_84 vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M74 p17_logic_ck_84 n1874_21 vdd vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M75 p17_logic_ck_12 n1874_15 vdd vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M76 vdd n1874_16 p17_logic_ck_36 vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M77 p17_logic_ck_36 n1874_17 vdd vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M78 vdd n1874_18 p17_logic_ck_60 vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M79 vdd n1874_14 p17_logic_ck_12 vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M80 vdd ck_10 n1874_22 vdd TP L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M81 n1874_24 ck_9 vdd vdd TP L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M82 vdd ck_8 n1874_24 vdd TP L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M83 n1874_26 ck_7 vdd vdd TP L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M84 a_0_2 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M85 vdd vdd a_0_2 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M86 a_0_4 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M87 vdd vdd a_0_4 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M88 vdd a_0_6 n5983_9 vdd TP L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M89 aa_0_1 n5983_4 vdd vdd TP L=0.18U W=10.332U AS=3.71952P AD=3.71952P 
+ PS=21.384U PD=21.384U 
M90 vdd n5983_3 aa_0_1 vdd TP L=0.18U W=10.332U AS=3.71952P AD=3.71952P 
+ PS=21.384U PD=21.384U 
M91 a_1_2 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M92 vdd vdd a_1_2 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M93 a_1_4 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M94 vdd vdd a_1_4 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M95 vdd a_1_6 n5139_9 vdd TP L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M96 aa_1_1 n5139_4 vdd vdd TP L=0.18U W=10.332U AS=3.71952P AD=3.71952P 
+ PS=21.384U PD=21.384U 
M97 vdd n5139_3 aa_1_1 vdd TP L=0.18U W=10.332U AS=3.71952P AD=3.71952P 
+ PS=21.384U PD=21.384U 
M98 a_2_2 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M99 vdd vdd a_2_2 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M100 a_2_4 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M101 vdd vdd a_2_4 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M102 vdd a_2_6 n3019_9 vdd TP L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M103 aa_2_15 n3019_4 vdd vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M104 vdd n3019_3 aa_2_15 vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M105 a_3_2 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M106 vdd vdd a_3_2 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M107 a_3_4 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M108 vdd vdd a_3_4 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M109 vdd a_3_6 n1981_9 vdd TP L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M110 aa_3_20 n1981_4 vdd vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M111 vdd n1981_3 aa_3_20 vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M112 b_0_2 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M113 vdd vdd b_0_2 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M114 b_0_4 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M115 vdd vdd b_0_4 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M116 vdd b_0_6 n1644_9 vdd TP L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M117 bb_0_39 n1644_4 vdd vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M118 vdd n1644_3 bb_0_39 vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M119 n6442_1 p17_logic_ck_3 vdd vdd TP L=0.18U W=7.272U AS=2.61792P 
+ AD=2.61792P PS=15.264U PD=15.264U 
M120 clock_2 n6442_2 vdd vdd TP L=0.18U W=6.192U AS=2.22912P AD=2.22912P 
+ PS=13.104U PD=13.104U 
M121 vdd n6442_3 clock_1 vdd TP L=0.18U W=6.192U AS=2.22912P AD=2.22912P 
+ PS=13.104U PD=13.104U 
M122 clock_1 n6442_12 vdd vdd TP L=0.18U W=6.192U AS=2.22912P AD=2.22912P 
+ PS=13.104U PD=13.104U 
M123 vdd n6442_4 clock_3 vdd TP L=0.18U W=6.192U AS=2.22912P AD=2.22912P 
+ PS=13.104U PD=13.104U 
M124 clock_3 n6442_5 vdd vdd TP L=0.18U W=6.192U AS=2.22912P AD=2.22912P 
+ PS=13.104U PD=13.104U 
M125 b_1_7 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M126 vdd vdd b_1_7 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M127 b_1_8 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M128 vdd vdd b_1_8 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M129 vdd b_1_6 n1625_13 vdd TP L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M130 bb_1_57 n1625_12 vdd vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M131 vdd n1625_11 bb_1_57 vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M132 b_2_7 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M133 vdd vdd b_2_7 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M134 b_2_8 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M135 vdd vdd b_2_8 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M136 vdd b_2_6 n1496_13 vdd TP L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M137 bb_2_51 n1496_12 vdd vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M138 vdd n1496_11 bb_2_51 vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M139 b_3_7 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M140 vdd vdd b_3_7 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M141 b_3_8 vdd vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M142 vdd vdd b_3_8 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M143 vdd b_3_6 n1367_13 vdd TP L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M144 bb_3_26 n1367_12 vdd vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M145 vdd n1367_11 bb_3_26 vdd TP L=0.18U W=10.332U AS=3.71952P 
+ AD=3.71952P PS=21.384U PD=21.384U 
M146 vdd n1110_56 s_0_12 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M147 s_0_12 n1110_59 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M148 vdd n1110_60 s_0_11 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M149 s_0_11 n1110_61 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M150 vdd n1110_50 s_0_10 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M151 s_0_10 n1110_53 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M152 vdd n1110_54 s_0_9 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M153 s_0_9 n1110_55 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M154 vdd n1110_44 s_0_8 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M155 s_0_8 n1110_47 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M156 vdd n1110_48 s_0_7 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M157 s_0_7 n1110_49 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M158 vdd n1110_38 s_0_6 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M159 s_0_6 n1110_41 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M160 vdd n1110_42 s_0_5 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M161 s_0_5 n1110_43 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M162 vdd n1110_32 s_0_4 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M163 s_0_4 n1110_35 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M164 vdd n1110_36 s_0_3 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M165 s_0_3 n1110_37 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M166 vdd n1110_26 s_0_2 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M167 s_0_2 n1110_29 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M168 vdd n1110_30 s_0_1 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M169 s_0_1 n1110_31 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M170 vdd n1228_6 n1110_25 vdd TP L=0.18U W=10.872U AS=3.91392P 
+ AD=3.91392P PS=22.464U PD=22.464U 
M171 n1110_25 n1228_7 vdd vdd TP L=0.18U W=10.872U AS=3.91392P 
+ AD=3.91392P PS=22.464U PD=22.464U 
M172 n1110_24 n1228_9 vdd vdd TP L=0.18U W=10.872U AS=3.91392P 
+ AD=3.91392P PS=22.464U PD=22.464U 
M173 vdd n1191_3 n1228_13 vdd TP L=0.18U W=10.872U AS=3.91392P 
+ AD=3.91392P PS=22.464U PD=22.464U 
M174 vdd n1228_8 n1110_24 vdd TP L=0.18U W=10.872U AS=3.91392P 
+ AD=3.91392P PS=22.464U PD=22.464U 
M175 n1191_5 ss_0_24 vdd vdd TP L=0.18U W=10.872U AS=3.91392P 
+ AD=3.91392P PS=22.464U PD=22.464U 
M176 vdd n939_56 s_1_12 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M177 s_1_12 n939_59 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M178 vdd n939_60 s_1_11 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M179 s_1_11 n939_61 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M180 vdd n939_50 s_1_10 vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M181 s_1_10 n939_53 vdd vdd TP L=0.18U W=14.472U AS=5.20992P 
+ AD=5.20992P PS=29.664U PD=29.664U 
M182 vdd n939_54 s_1_9 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M183 s_1_9 n939_55 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M184 vdd n939_44 s_1_8 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M185 s_1_8 n939_47 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M186 vdd n939_48 s_1_7 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M187 s_1_7 n939_49 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M188 vdd n939_38 s_1_6 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M189 s_1_6 n939_41 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M190 vdd n939_42 s_1_5 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M191 s_1_5 n939_43 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M192 vdd n939_32 s_1_4 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M193 s_1_4 n939_35 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M194 vdd n939_36 s_1_3 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M195 s_1_3 n939_37 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M196 vdd n939_26 s_1_2 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M197 s_1_2 n939_29 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M198 vdd n939_30 s_1_1 vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M199 s_1_1 n939_31 vdd vdd TP L=0.18U W=14.472U AS=5.20992P AD=5.20992P 
+ PS=29.664U PD=29.664U 
M200 vdd n817_6 n939_25 vdd TP L=0.18U W=10.872U AS=3.91392P AD=3.91392P 
+ PS=22.464U PD=22.464U 
M201 n939_25 n817_7 vdd vdd TP L=0.18U W=10.872U AS=3.91392P AD=3.91392P 
+ PS=22.464U PD=22.464U 
M202 n939_24 n817_9 vdd vdd TP L=0.18U W=10.872U AS=3.91392P AD=3.91392P 
+ PS=22.464U PD=22.464U 
M203 vdd n780_3 n817_13 vdd TP L=0.18U W=10.872U AS=3.91392P AD=3.91392P 
+ PS=22.464U PD=22.464U 
M204 vdd n817_8 n939_24 vdd TP L=0.18U W=10.872U AS=3.91392P AD=3.91392P 
+ PS=22.464U PD=22.464U 
M205 n780_5 ss_1_11 vdd vdd TP L=0.18U W=10.872U AS=3.91392P AD=3.91392P 
+ PS=22.464U PD=22.464U 
M206 n2142 core_mux_3_14 n2333_5 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M207 vdd bb_3_1 n2142 vdd TP L=0.18U W=4.212U AS=1.51632P AD=1.51632P 
+ PS=9.144U PD=9.144U 
M208 vdd bb_3_8 n2145_1 vdd TP L=0.18U W=4.212U AS=1.51632P AD=1.51632P 
+ PS=9.144U PD=9.144U 
M209 n2145 core_mux_3_22 vdd vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M210 core_int_9_9 n2333_2 n2145 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M211 n2160 core_int_9_20 n2381_5 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M212 vdd core_carry_2_23 n2160 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M213 vdd core_carry_2_30 n2151_1 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M214 n2151 core_int_9_23 vdd vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M215 ss_3_36 n2381_2 n2151 vdd TP L=0.18U W=4.212U AS=1.51632P AD=1.51632P 
+ PS=9.144U PD=9.144U 
M216 n2157 core_int_7_3 n2163 vdd TP L=0.18U W=2.952U AS=1.06272P AD=1.06272P 
+ PS=6.624U PD=6.624U 
M217 n2400_6 core_int_8_14 n2157 vdd TP L=0.18U W=2.952U AS=1.06272P 
+ AD=1.06272P PS=6.624U PD=6.624U 
M218 vdd n2400_3 core_carry_2_2 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M219 n2163 core_int_6_18 vdd vdd TP L=0.18U W=2.952U AS=1.06272P 
+ AD=1.06272P PS=6.624U PD=6.624U 
M220 n2166 core_int_5_15 n2412_5 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M221 vdd core_carry_1_47 n2166 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M222 vdd core_carry_1_54 n2169_1 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M223 n2169 core_int_5_23 vdd vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M224 ss_2_35 n2412_2 n2169 vdd TP L=0.18U W=4.212U AS=1.51632P AD=1.51632P 
+ PS=9.144U PD=9.144U 
M225 vdd n2427_2 core_int_8_7 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M226 vdd bb_2_27 n2427_5 vdd TP L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M227 n2427_5 core_carry_1_27 vdd vdd TP L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M228 vdd n2447_2 core_int_7_18 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M229 vdd core_mux_2_54 n2447_5 vdd TP L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M230 n2447_5 core_carry_1_16 vdd vdd TP L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M231 n2178 core_int_3_3 n2175 vdd TP L=0.18U W=2.952U AS=1.06272P AD=1.06272P 
+ PS=6.624U PD=6.624U 
M232 n2489_6 core_int_4_14 n2178 vdd TP L=0.18U W=2.952U AS=1.06272P 
+ AD=1.06272P PS=6.624U PD=6.624U 
M233 vdd n2489_3 core_carry_1_7 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M234 n2175 core_int_2_14 vdd vdd TP L=0.18U W=2.952U AS=1.06272P 
+ AD=1.06272P PS=6.624U PD=6.624U 
M235 vdd n2503_2 core_int_4_7 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M236 vdd bb_1_33 n2503_5 vdd TP L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M237 n2503_5 core_carry_0_48 vdd vdd TP L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M238 vdd n2517_2 core_int_3_18 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M239 vdd core_mux_1_39 n2517_5 vdd TP L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M240 n2517_5 core_carry_0_33 vdd vdd TP L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M241 n2566_2 n2624_13 vdd vdd TP L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M242 vdd core_l2_dff_m_3 n2624_2 vdd TP L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M243 n2593_6 clock_103 vdd vdd TP L=0.18U W=3.312U AS=1.19232P 
+ AD=1.19232P PS=7.344U PD=7.344U 
M244 core_l2_dff_s_2 n2561_3 vdd vdd TP L=0.72U W=0.432U AS=0.15552P 
+ AD=0.15552P PS=1.584U PD=1.584U 
M245 vdd core_l2_dff_s_8 n2561_5 vdd TP L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M246 core_regout_2_18 core_l2_dff_s_9 vdd vdd TP L=0.18U W=4.212U 
+ AS=1.51632P AD=1.51632P PS=9.144U PD=9.144U 
M247 core_l2_dff_m_2 n2624_5 vdd vdd TP L=0.72U W=0.432U AS=0.15552P 
+ AD=0.15552P PS=1.584U PD=1.584U 
M248 n2635_2 ss_2_17 vdd vdd TP L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M249 vdd n2646_2 core_carry_0_18 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M250 vdd core_mux_0_18 n2646_5 vdd TP L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M251 n2646_5 bb_0_12 vdd vdd TP L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M252 n2187 core_mux_0_28 n2733_5 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M253 vdd bb_0_1 n2187 vdd TP L=0.18U W=4.212U AS=1.51632P AD=1.51632P 
+ PS=9.144U PD=9.144U 
M254 vdd bb_0_8 n2181_1 vdd TP L=0.18U W=4.212U AS=1.51632P AD=1.51632P 
+ PS=9.144U PD=9.144U 
M255 n2181 core_mux_0_36 vdd vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M256 ss_0_13 n2733_2 n2181 vdd TP L=0.18U W=4.212U AS=1.51632P AD=1.51632P 
+ PS=9.144U PD=9.144U 
M257 n2770_2 n2837_13 vdd vdd TP L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M258 vdd core_l0_dff_m_3 n2837_2 vdd TP L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M259 n2750_6 clock_112 vdd vdd TP L=0.18U W=3.312U AS=1.19232P 
+ AD=1.19232P PS=7.344U PD=7.344U 
M260 core_l0_dff_s_2 n2765_2 vdd vdd TP L=0.72U W=0.432U AS=0.15552P 
+ AD=0.15552P PS=1.584U PD=1.584U 
M261 vdd core_l0_dff_s_8 n2765_5 vdd TP L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M262 core_regout_0_18 core_l0_dff_s_9 vdd vdd TP L=0.18U W=4.212U 
+ AS=1.51632P AD=1.51632P PS=9.144U PD=9.144U 
M263 core_l0_dff_m_2 n2837_5 vdd vdd TP L=0.72U W=0.432U AS=0.15552P 
+ AD=0.15552P PS=1.584U PD=1.584U 
M264 n2848_2 ss_0_1 vdd vdd TP L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M265 vdd aa_3_5 n3051_2 vdd TP L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M266 n3051_1 core_nsel_49 vdd vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M267 n3197_6 selsel_48 n3051_1 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M268 n3051 core_regout_3_22 n3197_6 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M269 core_mux_3_2 n3197_2 vdd vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M270 n3245_2 n3282_13 vdd vdd TP L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M271 vdd core_l3_dff_m_3 n3282_2 vdd TP L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M272 n3223_6 clock_75 vdd vdd TP L=0.18U W=3.312U AS=1.19232P AD=1.19232P 
+ PS=7.344U PD=7.344U 
M273 core_l3_dff_s_2 n3212_3 vdd vdd TP L=0.72U W=0.432U AS=0.15552P 
+ AD=0.15552P PS=1.584U PD=1.584U 
M274 vdd core_l3_dff_s_8 n3212_5 vdd TP L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M275 core_regout_3_2 core_l3_dff_s_9 vdd vdd TP L=0.18U W=4.212U 
+ AS=1.51632P AD=1.51632P PS=9.144U PD=9.144U 
M276 core_l3_dff_m_2 n3282_5 vdd vdd TP L=0.72U W=0.432U AS=0.15552P 
+ AD=0.15552P PS=1.584U PD=1.584U 
M277 n3252_2 ss_3_18 vdd vdd TP L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M278 n3068 core_mux_2_11 n3407_5 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M279 vdd bb_2_14 n3068 vdd TP L=0.18U W=4.212U AS=1.51632P AD=1.51632P 
+ PS=9.144U PD=9.144U 
M280 vdd bb_2_21 n3062_1 vdd TP L=0.18U W=4.212U AS=1.51632P AD=1.51632P 
+ PS=9.144U PD=9.144U 
M281 n3062 core_mux_2_14 vdd vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M282 core_int_5_2 n3407_2 n3062 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M283 vdd n3422_2 core_int_6_2 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M284 vdd core_mux_2_7 n3422_5 vdd TP L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M285 n3422_5 bb_2_1 vdd vdd TP L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M286 vdd aa_2_5 n3071_2 vdd TP L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M287 n3071_1 core_nsel_23 vdd vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M288 n3558_6 selsel_23 n3071_1 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M289 n3071 core_regout_2_1 n3558_6 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M290 core_mux_2_2 n3558_2 vdd vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M291 vdd selsel_33 core_nsel_32 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M292 vdd n3595_2 core_int_2_2 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M293 vdd core_mux_1_20 n3595_5 vdd TP L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M294 n3595_5 bb_1_22 vdd vdd TP L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M295 n3088 core_mux_1_7 n3746_5 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M296 vdd bb_1_5 n3088 vdd TP L=0.18U W=4.212U AS=1.51632P AD=1.51632P 
+ PS=9.144U PD=9.144U 
M297 vdd bb_1_2 n3082_1 vdd TP L=0.18U W=4.212U AS=1.51632P AD=1.51632P 
+ PS=9.144U PD=9.144U 
M298 n3082 core_mux_1_10 vdd vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M299 core_int_1_29 n3746_2 n3082 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M300 vdd aa_1_16 n3091_2 vdd TP L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M301 n3091_1 core_nsel_13 vdd vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M302 n3810_6 selsel_13 n3091_1 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M303 n3091 core_regout_1_5 n3810_6 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M304 core_mux_1_2 n3810_2 vdd vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M305 vdd aa_0_16 n3102_2 vdd TP L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M306 n3102_1 core_nsel_8 vdd vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M307 n3914_6 selsel_3 n3102_1 vdd TP L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M308 n3102 core_regout_0_1 n3914_6 vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M309 core_mux_0_2 n3914_2 vdd vdd TP L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M310 n3119 core_int_1_1 n4048_5 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M311 vdd core_carry_0_2 n3119 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M312 vdd core_carry_0_8 n3113_1 vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M313 n3113 core_int_1_4 vdd vdd TP L=0.18U W=4.212U AS=1.51632P 
+ AD=1.51632P PS=9.144U PD=9.144U 
M314 ss_1_37 n4048_2 n3113 vdd TP L=0.18U W=4.212U AS=1.51632P AD=1.51632P 
+ PS=9.144U PD=9.144U 
M315 n4085_2 n4115_13 vdd vdd TP L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M316 vdd core_l1_dff_m_3 n4115_2 vdd TP L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M317 n4065_6 clock_66 vdd vdd TP L=0.18U W=3.312U AS=1.19232P AD=1.19232P 
+ PS=7.344U PD=7.344U 
M318 core_l1_dff_s_2 n4080_2 vdd vdd TP L=0.72U W=0.432U AS=0.15552P 
+ AD=0.15552P PS=1.584U PD=1.584U 
M319 vdd core_l1_dff_s_8 n4080_5 vdd TP L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M320 core_regout_1_14 core_l1_dff_s_9 vdd vdd TP L=0.18U W=4.212U 
+ AS=1.51632P AD=1.51632P PS=9.144U PD=9.144U 
M321 core_l1_dff_m_2 n4115_5 vdd vdd TP L=0.72U W=0.432U AS=0.15552P 
+ AD=0.15552P PS=1.584U PD=1.584U 
M322 n4126_2 ss_1_20 vdd vdd TP L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M323 vss n5912_104 s_2_25 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M324 s_2_25 n5912_108 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M325 vss n5912_109 s_2_22 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M326 s_2_22 n5912_110 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M327 vss n5912_89 s_2_20 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M328 s_2_20 n5912_93 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M329 vss n5912_94 s_2_18 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M330 s_2_18 n5912_95 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M331 vss n5912_74 s_2_16 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M332 s_2_16 n5912_78 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M333 vss n5912_79 s_2_14 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M334 s_2_14 n5912_80 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M335 vss n5912_59 s_2_12 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M336 s_2_12 n5912_63 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M337 vss n5912_64 s_2_10 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M338 s_2_10 n5912_65 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M339 vss n5912_34 s_2_8 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M340 s_2_8 n5912_38 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M341 vss n5912_39 s_2_6 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M342 s_2_6 n5912_40 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M343 vss n5912_9 s_2_4 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M344 s_2_4 n5912_13 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M345 vss n5912_14 s_2_2 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M346 s_2_2 n5912_15 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M347 vss n5373_7 n5912_41 vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M348 n5912_41 n5373_8 vss vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M349 vss n5373_9 n5912 vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M350 n5912 n5373_10 vss vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M351 vss n5334_3 n5373 vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M352 n5334 ss_2_2 vss vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M353 vss n5111_104 s_3_25 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M354 s_3_25 n5111_108 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M355 vss n5111_109 s_3_22 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M356 s_3_22 n5111_110 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M357 vss n5111_89 s_3_20 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M358 s_3_20 n5111_93 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M359 vss n5111_94 s_3_18 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M360 s_3_18 n5111_95 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M361 vss n5111_74 s_3_16 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M362 s_3_16 n5111_78 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M363 vss n5111_79 s_3_14 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M364 s_3_14 n5111_80 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M365 vss n5111_59 s_3_12 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M366 s_3_12 n5111_63 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M367 vss n5111_64 s_3_10 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M368 s_3_10 n5111_65 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M369 vss n5111_34 s_3_8 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M370 s_3_8 n5111_38 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M371 vss n5111_39 s_3_6 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M372 s_3_6 n5111_40 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M373 vss n5111_9 s_3_4 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M374 s_3_4 n5111_13 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M375 vss n5111_14 s_3_2 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M376 s_3_2 n5111_15 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M377 vss n4572_7 n5111_41 vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M378 n5111_41 n4572_8 vss vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M379 vss n4572_9 n5111 vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M380 n5111 n4572_10 vss vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M381 vss n4533_3 n4572 vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M382 n4533 ss_3_4 vss vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M383 sel_2 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M384 vss vss sel_2 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M385 sel_4 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M386 vss vss sel_4 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M387 vss sel_5 n2124_13 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M388 n2124_13 sel_7 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M389 vss sel_8 n2124_9 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M390 vss n2124_3 selsel_66 vss TN L=0.18U W=4.932U AS=1.77552P 
+ AD=1.77552P PS=10.584U PD=10.584U 
M391 selsel_66 n2124 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M392 vss vss ck_4 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M393 ck_4 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M394 vss vss ck_2 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M395 ck_2 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M396 vss n1874_6 p17_logic_ck_35 vss TN L=0.18U W=4.932U AS=1.77552P 
+ AD=1.77552P PS=10.584U PD=10.584U 
M397 p17_logic_ck_11 n1874_5 vss vss TN L=0.18U W=4.932U AS=1.77552P 
+ AD=1.77552P PS=10.584U PD=10.584U 
M398 vss n1874_4 p17_logic_ck_11 vss TN L=0.18U W=4.932U AS=1.77552P 
+ AD=1.77552P PS=10.584U PD=10.584U 
M399 vss n1874_10 p17_logic_ck_83 vss TN L=0.18U W=4.932U AS=1.77552P 
+ AD=1.77552P PS=10.584U PD=10.584U 
M400 p17_logic_ck_59 n1874_9 vss vss TN L=0.18U W=4.932U AS=1.77552P 
+ AD=1.77552P PS=10.584U PD=10.584U 
M401 p17_logic_ck_83 n1874_11 vss vss TN L=0.18U W=4.932U AS=1.77552P 
+ AD=1.77552P PS=10.584U PD=10.584U 
M402 vss n1874_8 p17_logic_ck_59 vss TN L=0.18U W=4.932U AS=1.77552P 
+ AD=1.77552P PS=10.584U PD=10.584U 
M403 p17_logic_ck_35 n1874_7 vss vss TN L=0.18U W=4.932U AS=1.77552P 
+ AD=1.77552P PS=10.584U PD=10.584U 
M404 vss ck_25 n1874_1 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M405 n1874_23 ck_24 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M406 vss ck_23 n1874_23 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M407 n1874_25 ck_22 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M408 n1874_27 ck_20 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M409 vss ck_21 n1874_25 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M410 vss ck_15 n1874_28 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M411 vss ck_18 n1874_27 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M412 n1874_28 ck_17 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M413 n1874_30 ck_11 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M414 n1874 ck_14 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M415 vss ck_12 n1874 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M416 a_0_1 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M417 vss vss a_0_1 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M418 a_0_3 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M419 vss vss a_0_3 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M420 vss a_0_7 n5983_13 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M421 n5983_13 a_0_9 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M422 vss a_0_10 n5983_10 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M423 vss n5983_7 aa_0_2 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M424 aa_0_2 n5983 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M425 a_1_1 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M426 vss vss a_1_1 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M427 a_1_3 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M428 vss vss a_1_3 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M429 vss a_1_7 n5139_13 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M430 n5139_13 a_1_9 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M431 vss a_1_10 n5139_10 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M432 vss n5139_7 aa_1_2 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M433 aa_1_2 n5139 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M434 a_2_1 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M435 vss vss a_2_1 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M436 a_2_3 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M437 vss vss a_2_3 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M438 vss a_2_7 n3019_13 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M439 n3019_13 a_2_9 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M440 vss a_2_10 n3019_10 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M441 vss n3019_7 aa_2_19 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M442 aa_2_19 n3019 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M443 a_3_1 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M444 vss vss a_3_1 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M445 a_3_3 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M446 vss vss a_3_3 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M447 vss a_3_7 n1981_13 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M448 n1981_13 a_3_9 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M449 vss a_3_10 n1981_10 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M450 vss n1981_7 aa_3_19 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M451 aa_3_19 n1981 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M452 b_0_1 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M453 vss vss b_0_1 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M454 b_0_3 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M455 vss vss b_0_3 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M456 vss b_0_7 n1644_13 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M457 n1644_13 b_0_9 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M458 vss b_0_10 n1644_10 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M459 vss n1644_7 bb_0_42 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M460 bb_0_42 n1644 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M461 vss n6442_8 clock_5 vss TN L=0.18U W=3.672U AS=1.32192P AD=1.32192P 
+ PS=8.064U PD=8.064U 
M462 clock_5 n6442_9 vss vss TN L=0.18U W=3.672U AS=1.32192P AD=1.32192P 
+ PS=8.064U PD=8.064U 
M463 n6442_13 p17_logic_ck vss vss TN L=0.18U W=3.672U AS=1.32192P 
+ AD=1.32192P PS=8.064U PD=8.064U 
M464 clock_4 n6442_6 vss vss TN L=0.18U W=3.672U AS=1.32192P AD=1.32192P 
+ PS=8.064U PD=8.064U 
M465 vss n6442_7 clock_6 vss TN L=0.18U W=3.672U AS=1.32192P AD=1.32192P 
+ PS=8.064U PD=8.064U 
M466 clock_6 n6442 vss vss TN L=0.18U W=3.672U AS=1.32192P AD=1.32192P 
+ PS=8.064U PD=8.064U 
M467 b_1_9 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M468 vss vss b_1_9 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M469 b_1_10 vss vss vss TN L=0.18U W=6.372U AS=2.29392P 
+ AD=2.29392P PS=13.464U PD=13.464U 
M470 vss vss b_1_10 vss TN L=0.18U W=6.372U AS=2.29392P 
+ AD=2.29392P PS=13.464U PD=13.464U 
M471 vss b_1_1 n1625_8 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M472 n1625_8 b_1_3 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M473 vss b_1_4 n1625_7 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M474 vss n1625_5 bb_1_56 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M475 bb_1_56 n1625 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M476 b_2_9 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M477 vss vss b_2_9 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M478 b_2_10 vss vss vss TN L=0.18U W=6.372U AS=2.29392P 
+ AD=2.29392P PS=13.464U PD=13.464U 
M479 vss vss b_2_10 vss TN L=0.18U W=6.372U AS=2.29392P 
+ AD=2.29392P PS=13.464U PD=13.464U 
M480 vss b_2_1 n1496_8 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M481 n1496_8 b_2_3 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M482 vss b_2_4 n1496_7 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M483 vss n1496_5 bb_2_50 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M484 bb_2_50 n1496 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M485 b_3_9 vss vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M486 vss vss b_3_9 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M487 b_3_10 vss vss vss TN L=0.18U W=6.372U AS=2.29392P 
+ AD=2.29392P PS=13.464U PD=13.464U 
M488 vss vss b_3_10 vss TN L=0.18U W=6.372U AS=2.29392P 
+ AD=2.29392P PS=13.464U PD=13.464U 
M489 vss b_3_1 n1367_8 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M490 n1367_8 b_3_3 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M491 vss b_3_4 n1367_7 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M492 vss n1367_5 bb_3_25 vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M493 bb_3_25 n1367 vss vss TN L=0.18U W=4.932U AS=1.77552P AD=1.77552P 
+ PS=10.584U PD=10.584U 
M494 vss n1110_109 s_0_24 vss TN L=0.18U W=6.372U AS=2.29392P 
+ AD=2.29392P PS=13.464U PD=13.464U 
M495 s_0_24 n1110_113 vss vss TN L=0.18U W=6.372U AS=2.29392P 
+ AD=2.29392P PS=13.464U PD=13.464U 
M496 vss n1110_114 s_0_23 vss TN L=0.18U W=6.372U AS=2.29392P 
+ AD=2.29392P PS=13.464U PD=13.464U 
M497 s_0_23 n1110_115 vss vss TN L=0.18U W=6.372U AS=2.29392P 
+ AD=2.29392P PS=13.464U PD=13.464U 
M498 vss n1110_100 s_0_22 vss TN L=0.18U W=6.372U AS=2.29392P 
+ AD=2.29392P PS=13.464U PD=13.464U 
M499 s_0_22 n1110_104 vss vss TN L=0.18U W=6.372U AS=2.29392P 
+ AD=2.29392P PS=13.464U PD=13.464U 
M500 vss n1110_105 s_0_21 vss TN L=0.18U W=6.372U AS=2.29392P 
+ AD=2.29392P PS=13.464U PD=13.464U 
M501 s_0_21 n1110_106 vss vss TN L=0.18U W=6.372U AS=2.29392P 
+ AD=2.29392P PS=13.464U PD=13.464U 
M502 vss n1110_91 s_0_20 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M503 s_0_20 n1110_95 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M504 vss n1110_96 s_0_19 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M505 s_0_19 n1110_97 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M506 vss n1110_82 s_0_18 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M507 s_0_18 n1110_86 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M508 vss n1110_87 s_0_17 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M509 s_0_17 n1110_88 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M510 vss n1110_73 s_0_16 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M511 s_0_16 n1110_77 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M512 vss n1110_78 s_0_15 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M513 s_0_15 n1110_79 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M514 vss n1110_64 s_0_14 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M515 s_0_14 n1110_68 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M516 vss n1110_69 s_0_13 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M517 s_0_13 n1110_70 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M518 vss n1228_2 n1110_10 vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M519 n1110_10 n1228_3 vss vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M520 vss n1228_4 n1110 vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M521 n1110 n1228_5 vss vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M522 vss n1191_2 n1228 vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M523 n1191 ss_0_25 vss vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M524 vss n939_109 s_1_24 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M525 s_1_24 n939_113 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M526 vss n939_114 s_1_23 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M527 s_1_23 n939_115 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M528 vss n939_100 s_1_22 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M529 s_1_22 n939_104 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M530 vss n939_105 s_1_21 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M531 s_1_21 n939_106 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M532 vss n939_91 s_1_20 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M533 s_1_20 n939_95 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M534 vss n939_96 s_1_19 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M535 s_1_19 n939_97 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M536 vss n939_82 s_1_18 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M537 s_1_18 n939_86 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M538 vss n939_87 s_1_17 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M539 s_1_17 n939_88 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M540 vss n939_73 s_1_16 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M541 s_1_16 n939_77 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M542 vss n939_78 s_1_15 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M543 s_1_15 n939_79 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M544 vss n939_64 s_1_14 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M545 s_1_14 n939_68 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M546 vss n939_69 s_1_13 vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M547 s_1_13 n939_70 vss vss TN L=0.18U W=6.372U AS=2.29392P AD=2.29392P 
+ PS=13.464U PD=13.464U 
M548 vss n817_2 n939_10 vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M549 n939_10 n817_3 vss vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M550 vss n817_4 n939 vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M551 n939 n817_5 vss vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M552 vss n780_2 n817 vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M553 n780 ss_1_12 vss vss TN L=0.18U W=5.472U AS=1.96992P AD=1.96992P 
+ PS=11.664U PD=11.664U 
M554 n2333_1 core_mux_3_16 vss vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M555 vss bb_3_2 n2333_1 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M556 n2277 bb_3 vss vss TN L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M557 core_int_9_3 core_mux_3_24 n2277 vss TN L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M558 vss n2333 core_int_9_3 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M559 n2381_1 core_int_9_22 vss vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M560 vss core_carry_2_24 n2381_1 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M561 n2342 core_carry_2_31 vss vss TN L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M562 ss_3_37 core_int_9 n2342 vss TN L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M563 vss n2381 ss_3_37 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M564 vss n2400_5 core_carry_2 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M565 n2400_2 core_int_8_15 vss vss TN L=0.18U W=0.792U AS=0.28512P 
+ AD=0.28512P PS=2.304U PD=2.304U 
M566 vss core_int_7_4 n2400 vss TN L=0.18U W=0.792U AS=0.28512P 
+ AD=0.28512P PS=2.304U PD=2.304U 
M567 n2400 core_int_6_19 vss vss TN L=0.18U W=0.792U AS=0.28512P 
+ AD=0.28512P PS=2.304U PD=2.304U 
M568 n2412_1 core_int_5_17 vss vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M569 vss core_carry_1_48 n2412_1 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M570 n2405 core_carry_1_55 vss vss TN L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M571 ss_2_36 core_int_5_25 n2405 vss TN L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M572 vss n2412 ss_2_36 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M573 vss n2427_4 core_int_8 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M574 n2427 bb_2_28 n2438 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M575 n2438 core_carry_1_29 vss vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M576 vss n2447_4 core_int_7 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M577 n2447 core_mux_2_55 n2435 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M578 n2435 core_carry_1_18 vss vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M579 vss n2489_5 core_carry_1 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M580 n2489_2 core_int_4_15 vss vss TN L=0.18U W=0.792U AS=0.28512P 
+ AD=0.28512P PS=2.304U PD=2.304U 
M581 vss core_int_3_4 n2489 vss TN L=0.18U W=0.792U AS=0.28512P 
+ AD=0.28512P PS=2.304U PD=2.304U 
M582 n2489 core_int_2_15 vss vss TN L=0.18U W=0.792U AS=0.28512P 
+ AD=0.28512P PS=2.304U PD=2.304U 
M583 vss n2503_4 core_int_4 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M584 n2503 bb_1_34 n2494 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M585 n2494 core_carry_0_50 vss vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M586 vss n2517_4 core_int_3 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M587 n2517 core_mux_1_40 n2525 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M588 n2525 core_carry_0_35 vss vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M589 vss n2624_8 core_l2_dff_m vss TN L=1.26U W=0.612U AS=0.22032P 
+ AD=0.22032P PS=1.944U PD=1.944U 
M590 n2566 n2624_10 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M591 core_l2_dff_s_1 n2593_2 n2566 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M592 vss n2561_2 core_l2_dff_s_1 vss TN L=1.26U W=0.612U AS=0.22032P 
+ AD=0.22032P PS=1.944U PD=1.944U 
M593 vss core_l2_dff_m_5 n2624 vss TN L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M594 core_l2_dff_m clock_100 n2635 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M595 n2593 clock_105 vss vss TN L=0.18U W=1.692U AS=0.60912P AD=0.60912P 
+ PS=4.104U PD=4.104U 
M596 vss core_l2_dff_s_10 n2561 vss TN L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M597 core_regout_2_19 core_l2_dff_s vss vss TN L=0.18U W=2.232U 
+ AS=0.80352P AD=0.80352P PS=5.184U PD=5.184U 
M598 n2635 ss_2 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M599 vss n2646_4 core_carry_0_17 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M600 n2646 core_mux_0_19 n2654 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M601 n2654 bb_0_14 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M602 n2733_1 core_mux_0_30 vss vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M603 vss bb_0_2 n2733_1 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M604 n2657 bb_0 vss vss TN L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M605 ss_0_14 core_mux_0_38 n2657 vss TN L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M606 vss n2733 ss_0_14 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M607 vss n2837_8 core_l0_dff_m vss TN L=1.26U W=0.612U AS=0.22032P 
+ AD=0.22032P PS=1.944U PD=1.944U 
M608 n2770 n2837_10 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M609 core_l0_dff_s_1 n2750_2 n2770 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M610 vss n2765_4 core_l0_dff_s_1 vss TN L=1.26U W=0.612U AS=0.22032P 
+ AD=0.22032P PS=1.944U PD=1.944U 
M611 vss core_l0_dff_m_5 n2837 vss TN L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M612 core_l0_dff_m clock_109 n2848 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M613 n2750 clock_114 vss vss TN L=0.18U W=1.692U AS=0.60912P AD=0.60912P 
+ PS=4.104U PD=4.104U 
M614 vss core_l0_dff_s_10 n2765 vss TN L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M615 core_regout_0_19 core_l0_dff_s vss vss TN L=0.18U W=2.232U 
+ AS=0.80352P AD=0.80352P PS=5.184U PD=5.184U 
M616 n2848 ss_0 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M617 n3187 aa_3 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M618 n3197_1 core_nsel_51 n3187 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M619 n3184 selsel_50 n3197_1 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M620 vss core_regout_3_24 n3184 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M621 core_mux_3 n3197 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M622 vss n3282_8 core_l3_dff_m vss TN L=1.26U W=0.612U AS=0.22032P 
+ AD=0.22032P PS=1.944U PD=1.944U 
M623 n3245 n3282_10 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M624 core_l3_dff_s_1 n3223_2 n3245 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M625 vss n3212_2 core_l3_dff_s_1 vss TN L=1.26U W=0.612U AS=0.22032P 
+ AD=0.22032P PS=1.944U PD=1.944U 
M626 vss core_l3_dff_m_5 n3282 vss TN L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M627 core_l3_dff_m clock_72 n3252 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M628 n3223 clock_77 vss vss TN L=0.18U W=1.692U AS=0.60912P AD=0.60912P 
+ PS=4.104U PD=4.104U 
M629 vss core_l3_dff_s_10 n3212 vss TN L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M630 core_regout_3 core_l3_dff_s vss vss TN L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M631 n3252 ss_3 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M632 n3407_1 core_mux_2_13 vss vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M633 vss bb_2_15 n3407_1 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M634 n3291 bb_2_22 vss vss TN L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M635 core_int_5 core_mux_2_16 n3291 vss TN L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M636 vss n3407 core_int_5 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M637 vss n3422_4 core_int_6 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M638 n3422 core_mux_2_8 n3400 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M639 n3400 bb_2 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M640 n3548 aa_2 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M641 n3558_1 core_nsel_25 n3548 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M642 n3457 selsel_25 n3558_1 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M643 vss core_regout_2 n3457 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M644 core_mux_2 n3558 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M645 vss selsel_35 core_nsel_31 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M646 vss n3595_4 core_int_2 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M647 n3595 core_mux_1_21 n3603 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M648 n3603 bb_1_24 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M649 n3746_1 core_mux_1_9 vss vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M650 vss bb_1_6 n3746_1 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M651 n3686 bb_1 vss vss TN L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M652 core_int_1_23 core_mux_1_12 n3686 vss TN L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M653 vss n3746 core_int_1_23 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M654 n3800 aa_1 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M655 n3810_1 core_nsel_15 n3800 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M656 n3816 selsel_15 n3810_1 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M657 vss core_regout_1_7 n3816 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M658 core_mux_1 n3810 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M659 n3904 aa_0 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M660 n3914_1 core_nsel n3904 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M661 n3920 selsel n3914_1 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M662 vss core_regout_0 n3920 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M663 core_mux_0 n3914 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M664 n4048_1 core_int_1_3 vss vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M665 vss core_carry_0_4 n4048_1 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M666 n3923 core_carry_0 vss vss TN L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M667 ss_1_38 core_int_1 n3923 vss TN L=0.18U W=2.232U AS=0.80352P AD=0.80352P 
+ PS=5.184U PD=5.184U 
M668 vss n4048 ss_1_38 vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M669 vss n4115_8 core_l1_dff_m vss TN L=1.26U W=0.612U AS=0.22032P 
+ AD=0.22032P PS=1.944U PD=1.944U 
M670 n4085 n4115_10 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
M671 core_l1_dff_s_1 n4065_2 n4085 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M672 vss n4080_4 core_l1_dff_s_1 vss TN L=1.26U W=0.612U AS=0.22032P 
+ AD=0.22032P PS=1.944U PD=1.944U 
M673 vss core_l1_dff_m_5 n4115 vss TN L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M674 core_l1_dff_m clock_63 n4126 vss TN L=0.18U W=1.152U AS=0.41472P 
+ AD=0.41472P PS=3.024U PD=3.024U 
M675 n4065 clock vss vss TN L=0.18U W=1.692U AS=0.60912P AD=0.60912P 
+ PS=4.104U PD=4.104U 
M676 vss core_l1_dff_s_10 n4080 vss TN L=0.18U W=0.972U AS=0.34992P 
+ AD=0.34992P PS=2.664U PD=2.664U 
M677 core_regout_1 core_l1_dff_s vss vss TN L=0.18U W=2.232U AS=0.80352P 
+ AD=0.80352P PS=5.184U PD=5.184U 
M678 n4126 ss_1 vss vss TN L=0.18U W=1.152U AS=0.41472P AD=0.41472P 
+ PS=3.024U PD=3.024U 
R39_1 s_1_53 s_1_1 0.001
R39_2 s_1_54 s_1_1 0.001
R39_3 s_1_2 s_1_379 0.001
R39_4 s_1_2 s_1_380 0.001
R39_5 s_1_111 s_1_3 0.001
R39_6 s_1_112 s_1_3 0.001
R39_7 s_1_83 s_1_4 0.001
R39_8 s_1_82 s_1_4 0.001
R39_9 s_1_140 s_1_5 0.001
R39_10 s_1_141 s_1_5 0.001
R39_11 s_1_170 s_1_6 0.001
R39_12 s_1_169 s_1_6 0.001
R39_13 s_1_228 s_1_7 0.001
R39_14 s_1_227 s_1_7 0.001
R39_15 s_1_199 s_1_8 0.001
R39_16 s_1_198 s_1_8 0.001
R39_17 s_1_285 s_1_9 0.001
R39_18 s_1_286 s_1_9 0.001
R39_19 s_1_257 s_1_10 0.001
R39_20 s_1_256 s_1_10 0.001
R39_21 s_1_343 s_1_11 0.001
R39_22 s_1_344 s_1_11 0.001
R39_23 s_1_315 s_1_12 0.001
R39_24 s_1_314 s_1_12 0.001
R39_25 s_1_52 s_1_1 0.001
R39_26 s_1_2 s_1_378 0.001
R39_27 s_1_110 s_1_3 0.001
R39_28 s_1_81 s_1_4 0.001
R39_29 s_1_139 s_1_5 0.001
R39_30 s_1_168 s_1_6 0.001
R39_31 s_1_226 s_1_7 0.001
R39_32 s_1_197 s_1_8 0.001
R39_33 s_1_284 s_1_9 0.001
R39_34 s_1_255 s_1_10 0.001
R39_35 s_1_342 s_1_11 0.001
R39_36 s_1_313 s_1_12 0.001
R39_37 s_1_51 s_1_1 0.001
R39_38 s_1_2 s_1_377 0.001
R39_39 s_1_109 s_1_3 0.001
R39_40 s_1_80 s_1_4 0.001
R39_41 s_1_138 s_1_5 0.001
R39_42 s_1_167 s_1_6 0.001
R39_43 s_1_225 s_1_7 0.001
R39_44 s_1_196 s_1_8 0.001
R39_45 s_1_283 s_1_9 0.001
R39_46 s_1_254 s_1_10 0.001
R39_47 s_1_341 s_1_11 0.001
R39_48 s_1_312 s_1_12 0.001
R39_49 s_1_49 s_1_1 0.001
R39_50 s_1_50 s_1_1 0.001
R39_51 s_1_2 s_1_375 0.001
R39_52 s_1_2 s_1_376 0.001
R39_53 s_1_107 s_1_3 0.001
R39_54 s_1_108 s_1_3 0.001
R39_55 s_1_78 s_1_4 0.001
R39_56 s_1_79 s_1_4 0.001
R39_57 s_1_137 s_1_5 0.001
R39_58 s_1_136 s_1_5 0.001
R39_59 s_1_166 s_1_6 0.001
R39_60 s_1_165 s_1_6 0.001
R39_61 s_1_223 s_1_7 0.001
R39_62 s_1_224 s_1_7 0.001
R39_63 s_1_195 s_1_8 0.001
R39_64 s_1_194 s_1_8 0.001
R39_65 s_1_281 s_1_9 0.001
R39_66 s_1_282 s_1_9 0.001
R39_67 s_1_252 s_1_10 0.001
R39_68 s_1_253 s_1_10 0.001
R39_69 s_1_339 s_1_11 0.001
R39_70 s_1_340 s_1_11 0.001
R39_71 s_1_310 s_1_12 0.001
R39_72 s_1_311 s_1_12 0.001
R39_73 s_1_48 s_1_1 0.001
R39_74 s_1_2 s_1_374 0.001
R39_75 s_1_106 s_1_3 0.001
R39_76 s_1_77 s_1_4 0.001
R39_77 s_1_135 s_1_5 0.001
R39_78 s_1_164 s_1_6 0.001
R39_79 s_1_222 s_1_7 0.001
R39_80 s_1_193 s_1_8 0.001
R39_81 s_1_280 s_1_9 0.001
R39_82 s_1_251 s_1_10 0.001
R39_83 s_1_338 s_1_11 0.001
R39_84 s_1_309 s_1_12 0.001
R39_85 s_1_46 s_1_1 0.001
R39_86 s_1_47 s_1_1 0.001
R39_87 s_1_2 s_1_372 0.001
R39_88 s_1_2 s_1_373 0.001
R39_89 s_1_104 s_1_3 0.001
R39_90 s_1_105 s_1_3 0.001
R39_91 s_1_75 s_1_4 0.001
R39_92 s_1_76 s_1_4 0.001
R39_93 s_1_133 s_1_5 0.001
R39_94 s_1_134 s_1_5 0.001
R39_95 s_1_162 s_1_6 0.001
R39_96 s_1_163 s_1_6 0.001
R39_97 s_1_220 s_1_7 0.001
R39_98 s_1_221 s_1_7 0.001
R39_99 s_1_191 s_1_8 0.001
R39_100 s_1_192 s_1_8 0.001
R39_101 s_1_278 s_1_9 0.001
R39_102 s_1_279 s_1_9 0.001
R39_103 s_1_249 s_1_10 0.001
R39_104 s_1_250 s_1_10 0.001
R39_105 s_1_336 s_1_11 0.001
R39_106 s_1_337 s_1_11 0.001
R39_107 s_1_307 s_1_12 0.001
R39_108 s_1_308 s_1_12 0.001
R39_109 s_1_45 s_1_1 0.001
R39_110 s_1_2 s_1_371 0.001
R39_111 s_1_103 s_1_3 0.001
R39_112 s_1_74 s_1_4 0.001
R39_113 s_1_132 s_1_5 0.001
R39_114 s_1_161 s_1_6 0.001
R39_115 s_1_219 s_1_7 0.001
R39_116 s_1_190 s_1_8 0.001
R39_117 s_1_277 s_1_9 0.001
R39_118 s_1_248 s_1_10 0.001
R39_119 s_1_335 s_1_11 0.001
R39_120 s_1_306 s_1_12 0.001
R39_121 s_1_44 s_1_1 0.001
R39_122 s_1_2 s_1_370 0.001
R39_123 s_1_102 s_1_3 0.001
R39_124 s_1_73 s_1_4 0.001
R39_125 s_1_131 s_1_5 0.001
R39_126 s_1_160 s_1_6 0.001
R39_127 s_1_218 s_1_7 0.001
R39_128 s_1_189 s_1_8 0.001
R39_129 s_1_276 s_1_9 0.001
R39_130 s_1_247 s_1_10 0.001
R39_131 s_1_334 s_1_11 0.001
R39_132 s_1_305 s_1_12 0.001
R39_133 s_1_43 s_1_1 0.001
R39_134 s_1_42 s_1_1 0.001
R39_135 s_1_2 s_1_369 0.001
R39_136 s_1_2 s_1_368 0.001
R39_137 s_1_101 s_1_3 0.001
R39_138 s_1_100 s_1_3 0.001
R39_139 s_1_72 s_1_4 0.001
R39_140 s_1_71 s_1_4 0.001
R39_141 s_1_130 s_1_5 0.001
R39_142 s_1_129 s_1_5 0.001
R39_143 s_1_159 s_1_6 0.001
R39_144 s_1_158 s_1_6 0.001
R39_145 s_1_217 s_1_7 0.001
R39_146 s_1_216 s_1_7 0.001
R39_147 s_1_188 s_1_8 0.001
R39_148 s_1_187 s_1_8 0.001
R39_149 s_1_275 s_1_9 0.001
R39_150 s_1_274 s_1_9 0.001
R39_151 s_1_246 s_1_10 0.001
R39_152 s_1_245 s_1_10 0.001
R39_153 s_1_333 s_1_11 0.001
R39_154 s_1_332 s_1_11 0.001
R39_155 s_1_304 s_1_12 0.001
R39_156 s_1_303 s_1_12 0.001
R39_157 s_1_41 s_1_1 0.001
R39_158 s_1_2 s_1_367 0.001
R39_159 s_1_99 s_1_3 0.001
R39_160 s_1_70 s_1_4 0.001
R39_161 s_1_128 s_1_5 0.001
R39_162 s_1_157 s_1_6 0.001
R39_163 s_1_215 s_1_7 0.001
R39_164 s_1_186 s_1_8 0.001
R39_165 s_1_273 s_1_9 0.001
R39_166 s_1_244 s_1_10 0.001
R39_167 s_1_331 s_1_11 0.001
R39_168 s_1_302 s_1_12 0.001
R39_169 s_1_39 s_1_1 0.001
R39_170 s_1_40 s_1_1 0.001
R39_171 s_1_2 s_1_365 0.001
R39_172 s_1_2 s_1_366 0.001
R39_173 s_1_97 s_1_3 0.001
R39_174 s_1_98 s_1_3 0.001
R39_175 s_1_68 s_1_4 0.001
R39_176 s_1_69 s_1_4 0.001
R39_177 s_1_127 s_1_5 0.001
R39_178 s_1_126 s_1_5 0.001
R39_179 s_1_155 s_1_6 0.001
R39_180 s_1_156 s_1_6 0.001
R39_181 s_1_214 s_1_7 0.001
R39_182 s_1_213 s_1_7 0.001
R39_183 s_1_185 s_1_8 0.001
R39_184 s_1_184 s_1_8 0.001
R39_185 s_1_272 s_1_9 0.001
R39_186 s_1_271 s_1_9 0.001
R39_187 s_1_243 s_1_10 0.001
R39_188 s_1_242 s_1_10 0.001
R39_189 s_1_329 s_1_11 0.001
R39_190 s_1_330 s_1_11 0.001
R39_191 s_1_301 s_1_12 0.001
R39_192 s_1_300 s_1_12 0.001
R39_193 s_1_38 s_1_1 0.001
R39_194 s_1_2 s_1_364 0.001
R39_195 s_1_96 s_1_3 0.001
R39_196 s_1_67 s_1_4 0.001
R39_197 s_1_125 s_1_5 0.001
R39_198 s_1_154 s_1_6 0.001
R39_199 s_1_212 s_1_7 0.001
R39_200 s_1_183 s_1_8 0.001
R39_201 s_1_270 s_1_9 0.001
R39_202 s_1_241 s_1_10 0.001
R39_203 s_1_328 s_1_11 0.001
R39_204 s_1_299 s_1_12 0.001
R39_205 s_1_37 s_1_1 0.001
R39_206 s_1_2 s_1_363 0.001
R39_207 s_1_95 s_1_3 0.001
R39_208 s_1_66 s_1_4 0.001
R39_209 s_1_124 s_1_5 0.001
R39_210 s_1_153 s_1_6 0.001
R39_211 s_1_211 s_1_7 0.001
R39_212 s_1_182 s_1_8 0.001
R39_213 s_1_269 s_1_9 0.001
R39_214 s_1_240 s_1_10 0.001
R39_215 s_1_327 s_1_11 0.001
R39_216 s_1_298 s_1_12 0.001
R39_217 s_1_35 s_1_1 0.001
R39_218 s_1_36 s_1_1 0.001
R39_219 s_1_2 s_1_361 0.001
R39_220 s_1_2 s_1_362 0.001
R39_221 s_1_93 s_1_3 0.001
R39_222 s_1_94 s_1_3 0.001
R39_223 s_1_64 s_1_4 0.001
R39_224 s_1_65 s_1_4 0.001
R39_225 s_1_122 s_1_5 0.001
R39_226 s_1_123 s_1_5 0.001
R39_227 s_1_152 s_1_6 0.001
R39_228 s_1_151 s_1_6 0.001
R39_229 s_1_209 s_1_7 0.001
R39_230 s_1_210 s_1_7 0.001
R39_231 s_1_181 s_1_8 0.001
R39_232 s_1_180 s_1_8 0.001
R39_233 s_1_267 s_1_9 0.001
R39_234 s_1_268 s_1_9 0.001
R39_235 s_1_238 s_1_10 0.001
R39_236 s_1_239 s_1_10 0.001
R39_237 s_1_325 s_1_11 0.001
R39_238 s_1_326 s_1_11 0.001
R39_239 s_1_296 s_1_12 0.001
R39_240 s_1_297 s_1_12 0.001
R39_241 s_1_34 s_1_13 0.001
R39_242 s_1_33 s_1_13 0.001
R39_243 s_1_359 s_1_14 0.001
R39_244 s_1_360 s_1_14 0.001
R39_245 s_1_92 s_1_15 0.001
R39_246 s_1_91 s_1_15 0.001
R39_247 s_1_62 s_1_16 0.001
R39_248 s_1_63 s_1_16 0.001
R39_249 s_1_121 s_1_17 0.001
R39_250 s_1_120 s_1_17 0.001
R39_251 s_1_150 s_1_18 0.001
R39_252 s_1_149 s_1_18 0.001
R39_253 s_1_208 s_1_19 0.001
R39_254 s_1_207 s_1_19 0.001
R39_255 s_1_178 s_1_20 0.001
R39_256 s_1_179 s_1_20 0.001
R39_257 s_1_265 s_1_21 0.001
R39_258 s_1_266 s_1_21 0.001
R39_259 s_1_236 s_1_22 0.001
R39_260 s_1_237 s_1_22 0.001
R39_261 s_1_324 s_1_23 0.001
R39_262 s_1_323 s_1_23 0.001
R39_263 s_1_294 s_1_24 0.001
R39_264 s_1_295 s_1_24 0.001
R39_265 s_1_32 s_1_13 0.001
R39_266 s_1_358 s_1_14 0.001
R39_267 s_1_90 s_1_15 0.001
R39_268 s_1_61 s_1_16 0.001
R39_269 s_1_119 s_1_17 0.001
R39_270 s_1_148 s_1_18 0.001
R39_271 s_1_206 s_1_19 0.001
R39_272 s_1_177 s_1_20 0.001
R39_273 s_1_264 s_1_21 0.001
R39_274 s_1_235 s_1_22 0.001
R39_275 s_1_322 s_1_23 0.001
R39_276 s_1_293 s_1_24 0.001
R39_277 s_1_31 s_1_13 0.001
R39_278 s_1_357 s_1_14 0.001
R39_279 s_1_89 s_1_15 0.001
R39_280 s_1_60 s_1_16 0.001
R39_281 s_1_118 s_1_17 0.001
R39_282 s_1_147 s_1_18 0.001
R39_283 s_1_205 s_1_19 0.001
R39_284 s_1_176 s_1_20 0.001
R39_285 s_1_263 s_1_21 0.001
R39_286 s_1_234 s_1_22 0.001
R39_287 s_1_321 s_1_23 0.001
R39_288 s_1_292 s_1_24 0.001
R39_289 s_1_30 s_1_13 0.001
R39_290 s_1_29 s_1_13 0.001
R39_291 s_1_356 s_1_14 0.001
R39_292 s_1_355 s_1_14 0.001
R39_293 s_1_87 s_1_15 0.001
R39_294 s_1_88 s_1_15 0.001
R39_295 s_1_59 s_1_16 0.001
R39_296 s_1_58 s_1_16 0.001
R39_297 s_1_117 s_1_17 0.001
R39_298 s_1_116 s_1_17 0.001
R39_299 s_1_146 s_1_18 0.001
R39_300 s_1_145 s_1_18 0.001
R39_301 s_1_204 s_1_19 0.001
R39_302 s_1_203 s_1_19 0.001
R39_303 s_1_175 s_1_20 0.001
R39_304 s_1_174 s_1_20 0.001
R39_305 s_1_262 s_1_21 0.001
R39_306 s_1_261 s_1_21 0.001
R39_307 s_1_233 s_1_22 0.001
R39_308 s_1_232 s_1_22 0.001
R39_309 s_1_320 s_1_23 0.001
R39_310 s_1_319 s_1_23 0.001
R39_311 s_1_291 s_1_24 0.001
R39_312 s_1_290 s_1_24 0.001
R39_313 s_1_28 s_1_13 0.001
R39_314 s_1_354 s_1_14 0.001
R39_315 s_1_86 s_1_15 0.001
R39_316 s_1_57 s_1_16 0.001
R39_317 s_1_115 s_1_17 0.001
R39_318 s_1_144 s_1_18 0.001
R39_319 s_1_202 s_1_19 0.001
R39_320 s_1_173 s_1_20 0.001
R39_321 s_1_260 s_1_21 0.001
R39_322 s_1_231 s_1_22 0.001
R39_323 s_1_318 s_1_23 0.001
R39_324 s_1_289 s_1_24 0.001
R39_325 s_1_27 s_1_13 0.001
R39_326 s_1_353 s_1_14 0.001
R39_327 s_1_85 s_1_15 0.001
R39_328 s_1_56 s_1_16 0.001
R39_329 s_1_114 s_1_17 0.001
R39_330 s_1_143 s_1_18 0.001
R39_331 s_1_201 s_1_19 0.001
R39_332 s_1_172 s_1_20 0.001
R39_333 s_1_259 s_1_21 0.001
R39_334 s_1_230 s_1_22 0.001
R39_335 s_1_317 s_1_23 0.001
R39_336 s_1_288 s_1_24 0.001
R39_337 s_1 s_1_25 0.001
R39_338 s_1_349 s_1 0.108
R39_339 s_1_27 s_1_351 0.54
R39_340 s_1_28 s_1_27 0.108
R39_341 s_1_29 s_1_28 0.108
R39_342 s_1_30 s_1_29 0.108
R39_343 s_1_31 s_1_30 0.108
R39_344 s_1_32 s_1_31 0.108
R39_345 s_1_33 s_1_32 0.108
R39_346 s_1_34 s_1_33 0.108
R39_347 s_1_35 s_1_34 0.864
R39_348 s_1_36 s_1_35 0.108
R39_349 s_1_37 s_1_36 0.108
R39_350 s_1_38 s_1_37 0.108
R39_351 s_1_39 s_1_38 0.108
R39_352 s_1_40 s_1_39 0.108
R39_353 s_1_41 s_1_40 0.108
R39_354 s_1_42 s_1_41 0.108
R39_355 s_1_43 s_1_42 0.108
R39_356 s_1_44 s_1_43 0.108
R39_357 s_1_45 s_1_44 0.108
R39_358 s_1_46 s_1_45 0.108
R39_359 s_1_47 s_1_46 0.108
R39_360 s_1_48 s_1_47 0.108
R39_361 s_1_49 s_1_48 0.108
R39_362 s_1_50 s_1_49 0.108
R39_363 s_1_51 s_1_50 0.108
R39_364 s_1_52 s_1_51 0.108
R39_365 s_1_53 s_1_52 0.108
R39_366 s_1_54 s_1_53 0.108
R39_367 s_1_55 s_1_54 0.001
R39_368 s_1_56 s_1_349 1.296
R39_369 s_1_57 s_1_56 0.108
R39_370 s_1_58 s_1_57 0.108
R39_371 s_1_59 s_1_58 0.108
R39_372 s_1_60 s_1_59 0.108
R39_373 s_1_61 s_1_60 0.108
R39_374 s_1_62 s_1_61 0.108
R39_375 s_1_63 s_1_62 0.108
R39_376 s_1_64 s_1_63 0.864
R39_377 s_1_65 s_1_64 0.108
R39_378 s_1_66 s_1_65 0.108
R39_379 s_1_67 s_1_66 0.108
R39_380 s_1_68 s_1_67 0.108
R39_381 s_1_69 s_1_68 0.108
R39_382 s_1_70 s_1_69 0.108
R39_383 s_1_71 s_1_70 0.108
R39_384 s_1_72 s_1_71 0.108
R39_385 s_1_73 s_1_72 0.108
R39_386 s_1_74 s_1_73 0.108
R39_387 s_1_75 s_1_74 0.108
R39_388 s_1_76 s_1_75 0.108
R39_389 s_1_77 s_1_76 0.108
R39_390 s_1_78 s_1_77 0.108
R39_391 s_1_79 s_1_78 0.108
R39_392 s_1_80 s_1_79 0.108
R39_393 s_1_81 s_1_80 0.108
R39_394 s_1_82 s_1_81 0.108
R39_395 s_1_83 s_1_82 0.108
R39_396 s_1_84 s_1_83 0.001
R39_397 s_1_85 s_1_349 1.296
R39_398 s_1_86 s_1_85 0.108
R39_399 s_1_87 s_1_86 0.108
R39_400 s_1_88 s_1_87 0.108
R39_401 s_1_89 s_1_88 0.108
R39_402 s_1_90 s_1_89 0.108
R39_403 s_1_91 s_1_90 0.108
R39_404 s_1_92 s_1_91 0.108
R39_405 s_1_93 s_1_92 0.864
R39_406 s_1_94 s_1_93 0.108
R39_407 s_1_95 s_1_94 0.108
R39_408 s_1_96 s_1_95 0.108
R39_409 s_1_97 s_1_96 0.108
R39_410 s_1_98 s_1_97 0.108
R39_411 s_1_99 s_1_98 0.108
R39_412 s_1_100 s_1_99 0.108
R39_413 s_1_101 s_1_100 0.108
R39_414 s_1_102 s_1_101 0.108
R39_415 s_1_103 s_1_102 0.108
R39_416 s_1_104 s_1_103 0.108
R39_417 s_1_105 s_1_104 0.108
R39_418 s_1_106 s_1_105 0.108
R39_419 s_1_107 s_1_106 0.108
R39_420 s_1_108 s_1_107 0.108
R39_421 s_1_109 s_1_108 0.108
R39_422 s_1_110 s_1_109 0.108
R39_423 s_1_111 s_1_110 0.108
R39_424 s_1_112 s_1_111 0.108
R39_425 s_1_113 s_1_112 0.001
R39_426 s_1_114 s_1_349 1.296
R39_427 s_1_115 s_1_114 0.108
R39_428 s_1_116 s_1_115 0.108
R39_429 s_1_117 s_1_116 0.108
R39_430 s_1_118 s_1_117 0.108
R39_431 s_1_119 s_1_118 0.108
R39_432 s_1_120 s_1_119 0.108
R39_433 s_1_121 s_1_120 0.108
R39_434 s_1_122 s_1_121 0.864
R39_435 s_1_123 s_1_122 0.108
R39_436 s_1_124 s_1_123 0.108
R39_437 s_1_125 s_1_124 0.108
R39_438 s_1_126 s_1_125 0.108
R39_439 s_1_127 s_1_126 0.108
R39_440 s_1_128 s_1_127 0.108
R39_441 s_1_129 s_1_128 0.108
R39_442 s_1_130 s_1_129 0.108
R39_443 s_1_131 s_1_130 0.108
R39_444 s_1_132 s_1_131 0.108
R39_445 s_1_133 s_1_132 0.108
R39_446 s_1_134 s_1_133 0.108
R39_447 s_1_135 s_1_134 0.108
R39_448 s_1_136 s_1_135 0.108
R39_449 s_1_137 s_1_136 0.108
R39_450 s_1_138 s_1_137 0.108
R39_451 s_1_139 s_1_138 0.108
R39_452 s_1_140 s_1_139 0.108
R39_453 s_1_141 s_1_140 0.108
R39_454 s_1_142 s_1_141 0.001
R39_455 s_1_143 s_1_349 1.296
R39_456 s_1_144 s_1_143 0.108
R39_457 s_1_145 s_1_144 0.108
R39_458 s_1_146 s_1_145 0.108
R39_459 s_1_147 s_1_146 0.108
R39_460 s_1_148 s_1_147 0.108
R39_461 s_1_149 s_1_148 0.108
R39_462 s_1_150 s_1_149 0.108
R39_463 s_1_151 s_1_150 0.864
R39_464 s_1_152 s_1_151 0.108
R39_465 s_1_153 s_1_152 0.108
R39_466 s_1_154 s_1_153 0.108
R39_467 s_1_155 s_1_154 0.108
R39_468 s_1_156 s_1_155 0.108
R39_469 s_1_157 s_1_156 0.108
R39_470 s_1_158 s_1_157 0.108
R39_471 s_1_159 s_1_158 0.108
R39_472 s_1_160 s_1_159 0.108
R39_473 s_1_161 s_1_160 0.108
R39_474 s_1_162 s_1_161 0.108
R39_475 s_1_163 s_1_162 0.108
R39_476 s_1_164 s_1_163 0.108
R39_477 s_1_165 s_1_164 0.108
R39_478 s_1_166 s_1_165 0.108
R39_479 s_1_167 s_1_166 0.108
R39_480 s_1_168 s_1_167 0.108
R39_481 s_1_169 s_1_168 0.108
R39_482 s_1_170 s_1_169 0.108
R39_483 s_1_171 s_1_170 0.001
R39_484 s_1_172 s_1_349 1.296
R39_485 s_1_173 s_1_172 0.108
R39_486 s_1_174 s_1_173 0.108
R39_487 s_1_175 s_1_174 0.108
R39_488 s_1_176 s_1_175 0.108
R39_489 s_1_177 s_1_176 0.108
R39_490 s_1_178 s_1_177 0.108
R39_491 s_1_179 s_1_178 0.108
R39_492 s_1_180 s_1_179 0.864
R39_493 s_1_181 s_1_180 0.108
R39_494 s_1_182 s_1_181 0.108
R39_495 s_1_183 s_1_182 0.108
R39_496 s_1_184 s_1_183 0.108
R39_497 s_1_185 s_1_184 0.108
R39_498 s_1_186 s_1_185 0.108
R39_499 s_1_187 s_1_186 0.108
R39_500 s_1_188 s_1_187 0.108
R39_501 s_1_189 s_1_188 0.108
R39_502 s_1_190 s_1_189 0.108
R39_503 s_1_191 s_1_190 0.108
R39_504 s_1_192 s_1_191 0.108
R39_505 s_1_193 s_1_192 0.108
R39_506 s_1_194 s_1_193 0.108
R39_507 s_1_195 s_1_194 0.108
R39_508 s_1_196 s_1_195 0.108
R39_509 s_1_197 s_1_196 0.108
R39_510 s_1_198 s_1_197 0.108
R39_511 s_1_199 s_1_198 0.108
R39_512 s_1_200 s_1_199 0.001
R39_513 s_1_201 s_1_349 1.296
R39_514 s_1_202 s_1_201 0.108
R39_515 s_1_203 s_1_202 0.108
R39_516 s_1_204 s_1_203 0.108
R39_517 s_1_205 s_1_204 0.108
R39_518 s_1_206 s_1_205 0.108
R39_519 s_1_207 s_1_206 0.108
R39_520 s_1_208 s_1_207 0.108
R39_521 s_1_209 s_1_208 0.864
R39_522 s_1_210 s_1_209 0.108
R39_523 s_1_211 s_1_210 0.108
R39_524 s_1_212 s_1_211 0.108
R39_525 s_1_213 s_1_212 0.108
R39_526 s_1_214 s_1_213 0.108
R39_527 s_1_215 s_1_214 0.108
R39_528 s_1_216 s_1_215 0.108
R39_529 s_1_217 s_1_216 0.108
R39_530 s_1_218 s_1_217 0.108
R39_531 s_1_219 s_1_218 0.108
R39_532 s_1_220 s_1_219 0.108
R39_533 s_1_221 s_1_220 0.108
R39_534 s_1_222 s_1_221 0.108
R39_535 s_1_223 s_1_222 0.108
R39_536 s_1_224 s_1_223 0.108
R39_537 s_1_225 s_1_224 0.108
R39_538 s_1_226 s_1_225 0.108
R39_539 s_1_227 s_1_226 0.108
R39_540 s_1_228 s_1_227 0.108
R39_541 s_1_229 s_1_228 0.001
R39_542 s_1_230 s_1_349 1.296
R39_543 s_1_231 s_1_230 0.108
R39_544 s_1_232 s_1_231 0.108
R39_545 s_1_233 s_1_232 0.108
R39_546 s_1_234 s_1_233 0.108
R39_547 s_1_235 s_1_234 0.108
R39_548 s_1_236 s_1_235 0.108
R39_549 s_1_237 s_1_236 0.108
R39_550 s_1_238 s_1_237 0.864
R39_551 s_1_239 s_1_238 0.108
R39_552 s_1_240 s_1_239 0.108
R39_553 s_1_241 s_1_240 0.108
R39_554 s_1_242 s_1_241 0.108
R39_555 s_1_243 s_1_242 0.108
R39_556 s_1_244 s_1_243 0.108
R39_557 s_1_245 s_1_244 0.108
R39_558 s_1_246 s_1_245 0.108
R39_559 s_1_247 s_1_246 0.108
R39_560 s_1_248 s_1_247 0.108
R39_561 s_1_249 s_1_248 0.108
R39_562 s_1_250 s_1_249 0.108
R39_563 s_1_251 s_1_250 0.108
R39_564 s_1_252 s_1_251 0.108
R39_565 s_1_253 s_1_252 0.108
R39_566 s_1_254 s_1_253 0.108
R39_567 s_1_255 s_1_254 0.108
R39_568 s_1_256 s_1_255 0.108
R39_569 s_1_257 s_1_256 0.108
R39_570 s_1_258 s_1_257 0.001
R39_571 s_1_259 s_1_349 1.296
R39_572 s_1_260 s_1_259 0.108
R39_573 s_1_261 s_1_260 0.108
R39_574 s_1_262 s_1_261 0.108
R39_575 s_1_263 s_1_262 0.108
R39_576 s_1_264 s_1_263 0.108
R39_577 s_1_265 s_1_264 0.108
R39_578 s_1_266 s_1_265 0.108
R39_579 s_1_267 s_1_266 0.864
R39_580 s_1_268 s_1_267 0.108
R39_581 s_1_269 s_1_268 0.108
R39_582 s_1_270 s_1_269 0.108
R39_583 s_1_271 s_1_270 0.108
R39_584 s_1_272 s_1_271 0.108
R39_585 s_1_273 s_1_272 0.108
R39_586 s_1_274 s_1_273 0.108
R39_587 s_1_275 s_1_274 0.108
R39_588 s_1_276 s_1_275 0.108
R39_589 s_1_277 s_1_276 0.108
R39_590 s_1_278 s_1_277 0.108
R39_591 s_1_279 s_1_278 0.108
R39_592 s_1_280 s_1_279 0.108
R39_593 s_1_281 s_1_280 0.108
R39_594 s_1_282 s_1_281 0.108
R39_595 s_1_283 s_1_282 0.108
R39_596 s_1_284 s_1_283 0.108
R39_597 s_1_285 s_1_284 0.108
R39_598 s_1_286 s_1_285 0.108
R39_599 s_1_287 s_1_286 0.001
R39_600 s_1_288 s_1_346 0.54
R39_601 s_1_289 s_1_288 0.108
R39_602 s_1_290 s_1_289 0.108
R39_603 s_1_291 s_1_290 0.108
R39_604 s_1_292 s_1_291 0.108
R39_605 s_1_293 s_1_292 0.108
R39_606 s_1_294 s_1_293 0.108
R39_607 s_1_295 s_1_294 0.108
R39_608 s_1_296 s_1_295 0.864
R39_609 s_1_297 s_1_296 0.108
R39_610 s_1_298 s_1_297 0.108
R39_611 s_1_299 s_1_298 0.108
R39_612 s_1_300 s_1_299 0.108
R39_613 s_1_301 s_1_300 0.108
R39_614 s_1_302 s_1_301 0.108
R39_615 s_1_303 s_1_302 0.108
R39_616 s_1_304 s_1_303 0.108
R39_617 s_1_305 s_1_304 0.108
R39_618 s_1_306 s_1_305 0.108
R39_619 s_1_307 s_1_306 0.108
R39_620 s_1_308 s_1_307 0.108
R39_621 s_1_309 s_1_308 0.108
R39_622 s_1_310 s_1_309 0.108
R39_623 s_1_311 s_1_310 0.108
R39_624 s_1_312 s_1_311 0.108
R39_625 s_1_313 s_1_312 0.108
R39_626 s_1_314 s_1_313 0.108
R39_627 s_1_315 s_1_314 0.108
R39_628 s_1_316 s_1_315 0.001
R39_629 s_1_317 s_1_348 0.54
R39_630 s_1_318 s_1_317 0.108
R39_631 s_1_319 s_1_318 0.108
R39_632 s_1_320 s_1_319 0.108
R39_633 s_1_321 s_1_320 0.108
R39_634 s_1_322 s_1_321 0.108
R39_635 s_1_323 s_1_322 0.108
R39_636 s_1_324 s_1_323 0.108
R39_637 s_1_325 s_1_324 0.864
R39_638 s_1_326 s_1_325 0.108
R39_639 s_1_327 s_1_326 0.108
R39_640 s_1_328 s_1_327 0.108
R39_641 s_1_329 s_1_328 0.108
R39_642 s_1_330 s_1_329 0.108
R39_643 s_1_331 s_1_330 0.108
R39_644 s_1_332 s_1_331 0.108
R39_645 s_1_333 s_1_332 0.108
R39_646 s_1_334 s_1_333 0.108
R39_647 s_1_335 s_1_334 0.108
R39_648 s_1_336 s_1_335 0.108
R39_649 s_1_337 s_1_336 0.108
R39_650 s_1_338 s_1_337 0.108
R39_651 s_1_339 s_1_338 0.108
R39_652 s_1_340 s_1_339 0.108
R39_653 s_1_341 s_1_340 0.108
R39_654 s_1_342 s_1_341 0.108
R39_655 s_1_343 s_1_342 0.108
R39_656 s_1_344 s_1_343 0.108
R39_657 s_1_345 s_1_344 0.001
R39_658 s_1_347 s_1_346 0.001
R39_659 s_1_348 s_1_347 0.001
R39_660 s_1_349 s_1_348 0.001
R39_661 s_1_352 s_1_349 0.001
R39_662 s_1_350 s_1_352 0.001
R39_663 s_1_351 s_1_350 0.001
R39_664 s_1_353 s_1_352 0.54
R39_665 s_1_354 s_1_353 0.108
R39_666 s_1_355 s_1_354 0.108
R39_667 s_1_356 s_1_355 0.108
R39_668 s_1_357 s_1_356 0.108
R39_669 s_1_358 s_1_357 0.108
R39_670 s_1_359 s_1_358 0.108
R39_671 s_1_360 s_1_359 0.108
R39_672 s_1_361 s_1_360 0.864
R39_673 s_1_362 s_1_361 0.108
R39_674 s_1_363 s_1_362 0.108
R39_675 s_1_364 s_1_363 0.108
R39_676 s_1_365 s_1_364 0.108
R39_677 s_1_366 s_1_365 0.108
R39_678 s_1_367 s_1_366 0.108
R39_679 s_1_368 s_1_367 0.108
R39_680 s_1_369 s_1_368 0.108
R39_681 s_1_370 s_1_369 0.108
R39_682 s_1_371 s_1_370 0.108
R39_683 s_1_372 s_1_371 0.108
R39_684 s_1_373 s_1_372 0.108
R39_685 s_1_374 s_1_373 0.108
R39_686 s_1_375 s_1_374 0.108
R39_687 s_1_376 s_1_375 0.108
R39_688 s_1_377 s_1_376 0.108
R39_689 s_1_378 s_1_377 0.108
R39_690 s_1_379 s_1_378 0.108
R39_691 s_1_380 s_1_379 0.108
R39_692 s_1_381 s_1_380 0.001

C0 s_1_349 vss 6.29069e-15
C1 s_1 vss 6.29069e-15
C2 s_1_27 vss 1.40901e-16
C3 s_1_351 vss 1.40901e-16
C4 s_1_28 vss 3.13114e-17
C5 s_1_27 vss 3.13114e-17
C6 s_1_29 vss 3.13114e-17
C7 s_1_28 vss 3.13114e-17
C8 s_1_30 vss 3.13114e-17
C9 s_1_29 vss 3.13114e-17
C10 s_1_31 vss 3.13114e-17
C11 s_1_30 vss 3.13114e-17
C12 s_1_32 vss 3.13114e-17
C13 s_1_31 vss 3.13114e-17
C14 s_1_33 vss 3.13114e-17
C15 s_1_32 vss 3.13114e-17
C16 s_1_34 vss 3.13114e-17
C17 s_1_33 vss 3.13114e-17
C18 s_1_35 vss 2.42663e-16
C19 s_1_34 vss 2.42663e-16
C20 s_1_36 vss 3.13114e-17
C21 s_1_35 vss 3.13114e-17
C22 s_1_37 vss 3.13114e-17
C23 s_1_36 vss 3.13114e-17
C24 s_1_38 vss 3.13114e-17
C25 s_1_37 vss 3.13114e-17
C26 s_1_39 vss 3.13114e-17
C27 s_1_38 vss 3.13114e-17
C28 s_1_40 vss 3.13114e-17
C29 s_1_39 vss 3.13114e-17
C30 s_1_41 vss 3.13114e-17
C31 s_1_40 vss 3.13114e-17
C32 s_1_42 vss 3.13114e-17
C33 s_1_41 vss 3.13114e-17
C34 s_1_43 vss 3.13114e-17
C35 s_1_42 vss 3.13114e-17
C36 s_1_44 vss 3.13114e-17
C37 s_1_43 vss 3.13114e-17
C38 s_1_45 vss 3.13114e-17
C39 s_1_44 vss 3.13114e-17
C40 s_1_46 vss 3.13114e-17
C41 s_1_45 vss 3.13114e-17
C42 s_1_47 vss 3.13114e-17
C43 s_1_46 vss 3.13114e-17
C44 s_1_48 vss 3.13114e-17
C45 s_1_47 vss 3.13114e-17
C46 s_1_49 vss 3.13114e-17
C47 s_1_48 vss 3.13114e-17
C48 s_1_50 vss 3.13114e-17
C49 s_1_49 vss 3.13114e-17
C50 s_1_51 vss 3.13114e-17
C51 s_1_50 vss 3.13114e-17
C52 s_1_52 vss 3.13114e-17
C53 s_1_51 vss 3.13114e-17
C54 s_1_53 vss 3.13114e-17
C55 s_1_52 vss 3.13114e-17
C56 s_1_54 vss 3.13114e-17
C57 s_1_53 vss 3.13114e-17
C58 s_1_55 vss 1.40901e-17
C59 s_1_54 vss 1.40901e-17
C60 s_1_56 vss 3.60081e-16
C61 s_1_349 vss 3.60081e-16
C62 s_1_57 vss 3.13114e-17
C63 s_1_56 vss 3.13114e-17
C64 s_1_58 vss 3.13114e-17
C65 s_1_57 vss 3.13114e-17
C66 s_1_59 vss 3.13114e-17
C67 s_1_58 vss 3.13114e-17
C68 s_1_60 vss 3.13114e-17
C69 s_1_59 vss 3.13114e-17
C70 s_1_61 vss 3.13114e-17
C71 s_1_60 vss 3.13114e-17
C72 s_1_62 vss 3.13114e-17
C73 s_1_61 vss 3.13114e-17
C74 s_1_63 vss 3.13114e-17
C75 s_1_62 vss 3.13114e-17
C76 s_1_64 vss 2.42663e-16
C77 s_1_63 vss 2.42663e-16
C78 s_1_65 vss 3.13114e-17
C79 s_1_64 vss 3.13114e-17
C80 s_1_66 vss 3.13114e-17
C81 s_1_65 vss 3.13114e-17
C82 s_1_67 vss 3.13114e-17
C83 s_1_66 vss 3.13114e-17
C84 s_1_68 vss 3.13114e-17
C85 s_1_67 vss 3.13114e-17
C86 s_1_69 vss 3.13114e-17
C87 s_1_68 vss 3.13114e-17
C88 s_1_70 vss 3.13114e-17
C89 s_1_69 vss 3.13114e-17
C90 s_1_71 vss 3.13114e-17
C91 s_1_70 vss 3.13114e-17
C92 s_1_72 vss 3.13114e-17
C93 s_1_71 vss 3.13114e-17
C94 s_1_73 vss 3.13114e-17
C95 s_1_72 vss 3.13114e-17
C96 s_1_74 vss 3.13114e-17
C97 s_1_73 vss 3.13114e-17
C98 s_1_75 vss 3.13114e-17
C99 s_1_74 vss 3.13114e-17
C100 s_1_76 vss 3.13114e-17
C101 s_1_75 vss 3.13114e-17
C102 s_1_77 vss 3.13114e-17
C103 s_1_76 vss 3.13114e-17
C104 s_1_78 vss 3.13114e-17
C105 s_1_77 vss 3.13114e-17
C106 s_1_79 vss 3.13114e-17
C107 s_1_78 vss 3.13114e-17
C108 s_1_80 vss 3.13114e-17
C109 s_1_79 vss 3.13114e-17
C110 s_1_81 vss 3.13114e-17
C111 s_1_80 vss 3.13114e-17
C112 s_1_82 vss 3.13114e-17
C113 s_1_81 vss 3.13114e-17
C114 s_1_83 vss 3.13114e-17
C115 s_1_82 vss 3.13114e-17
C116 s_1_84 vss 1.40901e-17
C117 s_1_83 vss 1.40901e-17
C118 s_1_85 vss 3.60081e-16
C119 s_1_349 vss 3.60081e-16
C120 s_1_86 vss 3.13114e-17
C121 s_1_85 vss 3.13114e-17
C122 s_1_87 vss 3.13114e-17
C123 s_1_86 vss 3.13114e-17
C124 s_1_88 vss 3.13114e-17
C125 s_1_87 vss 3.13114e-17
C126 s_1_89 vss 3.13114e-17
C127 s_1_88 vss 3.13114e-17
C128 s_1_90 vss 3.13114e-17
C129 s_1_89 vss 3.13114e-17
C130 s_1_91 vss 3.13114e-17
C131 s_1_90 vss 3.13114e-17
C132 s_1_92 vss 3.13114e-17
C133 s_1_91 vss 3.13114e-17
C134 s_1_93 vss 2.42663e-16
C135 s_1_92 vss 2.42663e-16
C136 s_1_94 vss 3.13114e-17
C137 s_1_93 vss 3.13114e-17
C138 s_1_95 vss 3.13114e-17
C139 s_1_94 vss 3.13114e-17
C140 s_1_96 vss 3.13114e-17
C141 s_1_95 vss 3.13114e-17
C142 s_1_97 vss 3.13114e-17
C143 s_1_96 vss 3.13114e-17
C144 s_1_98 vss 3.13114e-17
C145 s_1_97 vss 3.13114e-17
C146 s_1_99 vss 3.13114e-17
C147 s_1_98 vss 3.13114e-17
C148 s_1_100 vss 3.13114e-17
C149 s_1_99 vss 3.13114e-17
C150 s_1_101 vss 3.13114e-17
C151 s_1_100 vss 3.13114e-17
C152 s_1_102 vss 3.13114e-17
C153 s_1_101 vss 3.13114e-17
C154 s_1_103 vss 3.13114e-17
C155 s_1_102 vss 3.13114e-17
C156 s_1_104 vss 3.13114e-17
C157 s_1_103 vss 3.13114e-17
C158 s_1_105 vss 3.13114e-17
C159 s_1_104 vss 3.13114e-17
C160 s_1_106 vss 3.13114e-17
C161 s_1_105 vss 3.13114e-17
C162 s_1_107 vss 3.13114e-17
C163 s_1_106 vss 3.13114e-17
C164 s_1_108 vss 3.13114e-17
C165 s_1_107 vss 3.13114e-17
C166 s_1_109 vss 3.13114e-17
C167 s_1_108 vss 3.13114e-17
C168 s_1_110 vss 3.13114e-17
C169 s_1_109 vss 3.13114e-17
C170 s_1_111 vss 3.13114e-17
C171 s_1_110 vss 3.13114e-17
C172 s_1_112 vss 3.13114e-17
C173 s_1_111 vss 3.13114e-17
C174 s_1_113 vss 1.40901e-17
C175 s_1_112 vss 1.40901e-17
C176 s_1_114 vss 3.60081e-16
C177 s_1_349 vss 3.60081e-16
C178 s_1_115 vss 3.13114e-17
C179 s_1_114 vss 3.13114e-17
C180 s_1_116 vss 3.13114e-17
C181 s_1_115 vss 3.13114e-17
C182 s_1_117 vss 3.13114e-17
C183 s_1_116 vss 3.13114e-17
C184 s_1_118 vss 3.13114e-17
C185 s_1_117 vss 3.13114e-17
C186 s_1_119 vss 3.13114e-17
C187 s_1_118 vss 3.13114e-17
C188 s_1_120 vss 3.13114e-17
C189 s_1_119 vss 3.13114e-17
C190 s_1_121 vss 3.13114e-17
C191 s_1_120 vss 3.13114e-17
C192 s_1_122 vss 2.42663e-16
C193 s_1_121 vss 2.42663e-16
C194 s_1_123 vss 3.13114e-17
C195 s_1_122 vss 3.13114e-17
C196 s_1_124 vss 3.13114e-17
C197 s_1_123 vss 3.13114e-17
C198 s_1_125 vss 3.13114e-17
C199 s_1_124 vss 3.13114e-17
C200 s_1_126 vss 3.13114e-17
C201 s_1_125 vss 3.13114e-17
C202 s_1_127 vss 3.13114e-17
C203 s_1_126 vss 3.13114e-17
C204 s_1_128 vss 3.13114e-17
C205 s_1_127 vss 3.13114e-17
C206 s_1_129 vss 3.13114e-17
C207 s_1_128 vss 3.13114e-17
C208 s_1_130 vss 3.13114e-17
C209 s_1_129 vss 3.13114e-17
C210 s_1_131 vss 3.13114e-17
C211 s_1_130 vss 3.13114e-17
C212 s_1_132 vss 3.13114e-17
C213 s_1_131 vss 3.13114e-17
C214 s_1_133 vss 3.13114e-17
C215 s_1_132 vss 3.13114e-17
C216 s_1_134 vss 3.13114e-17
C217 s_1_133 vss 3.13114e-17
C218 s_1_135 vss 3.13114e-17
C219 s_1_134 vss 3.13114e-17
C220 s_1_136 vss 3.13114e-17
C221 s_1_135 vss 3.13114e-17
C222 s_1_137 vss 3.13114e-17
C223 s_1_136 vss 3.13114e-17
C224 s_1_138 vss 3.13114e-17
C225 s_1_137 vss 3.13114e-17
C226 s_1_139 vss 3.13114e-17
C227 s_1_138 vss 3.13114e-17
C228 s_1_140 vss 3.13114e-17
C229 s_1_139 vss 3.13114e-17
C230 s_1_141 vss 3.13114e-17
C231 s_1_140 vss 3.13114e-17
C232 s_1_142 vss 1.40901e-17
C233 s_1_141 vss 1.40901e-17
C234 s_1_143 vss 3.60081e-16
C235 s_1_349 vss 3.60081e-16
C236 s_1_144 vss 3.13114e-17
C237 s_1_143 vss 3.13114e-17
C238 s_1_145 vss 3.13114e-17
C239 s_1_144 vss 3.13114e-17
C240 s_1_146 vss 3.13114e-17
C241 s_1_145 vss 3.13114e-17
C242 s_1_147 vss 3.13114e-17
C243 s_1_146 vss 3.13114e-17
C244 s_1_148 vss 3.13114e-17
C245 s_1_147 vss 3.13114e-17
C246 s_1_149 vss 3.13114e-17
C247 s_1_148 vss 3.13114e-17
C248 s_1_150 vss 3.13114e-17
C249 s_1_149 vss 3.13114e-17
C250 s_1_151 vss 2.42663e-16
C251 s_1_150 vss 2.42663e-16
C252 s_1_152 vss 3.13114e-17
C253 s_1_151 vss 3.13114e-17
C254 s_1_153 vss 3.13114e-17
C255 s_1_152 vss 3.13114e-17
C256 s_1_154 vss 3.13114e-17
C257 s_1_153 vss 3.13114e-17
C258 s_1_155 vss 3.13114e-17
C259 s_1_154 vss 3.13114e-17
C260 s_1_156 vss 3.13114e-17
C261 s_1_155 vss 3.13114e-17
C262 s_1_157 vss 3.13114e-17
C263 s_1_156 vss 3.13114e-17
C264 s_1_158 vss 3.13114e-17
C265 s_1_157 vss 3.13114e-17
C266 s_1_159 vss 3.13114e-17
C267 s_1_158 vss 3.13114e-17
C268 s_1_160 vss 3.13114e-17
C269 s_1_159 vss 3.13114e-17
C270 s_1_161 vss 3.13114e-17
C271 s_1_160 vss 3.13114e-17
C272 s_1_162 vss 3.13114e-17
C273 s_1_161 vss 3.13114e-17
C274 s_1_163 vss 3.13114e-17
C275 s_1_162 vss 3.13114e-17
C276 s_1_164 vss 3.13114e-17
C277 s_1_163 vss 3.13114e-17
C278 s_1_165 vss 3.13114e-17
C279 s_1_164 vss 3.13114e-17
C280 s_1_166 vss 3.13114e-17
C281 s_1_165 vss 3.13114e-17
C282 s_1_167 vss 3.13114e-17
C283 s_1_166 vss 3.13114e-17
C284 s_1_168 vss 3.13114e-17
C285 s_1_167 vss 3.13114e-17
C286 s_1_169 vss 3.13114e-17
C287 s_1_168 vss 3.13114e-17
C288 s_1_170 vss 3.13114e-17
C289 s_1_169 vss 3.13114e-17
C290 s_1_171 vss 1.40901e-17
C291 s_1_170 vss 1.40901e-17
C292 s_1_172 vss 3.60081e-16
C293 s_1_349 vss 3.60081e-16
C294 s_1_173 vss 3.13114e-17
C295 s_1_172 vss 3.13114e-17
C296 s_1_174 vss 3.13114e-17
C297 s_1_173 vss 3.13114e-17
C298 s_1_175 vss 3.13114e-17
C299 s_1_174 vss 3.13114e-17
C300 s_1_176 vss 3.13114e-17
C301 s_1_175 vss 3.13114e-17
C302 s_1_177 vss 3.13114e-17
C303 s_1_176 vss 3.13114e-17
C304 s_1_178 vss 3.13114e-17
C305 s_1_177 vss 3.13114e-17
C306 s_1_179 vss 3.13114e-17
C307 s_1_178 vss 3.13114e-17
C308 s_1_180 vss 2.42663e-16
C309 s_1_179 vss 2.42663e-16
C310 s_1_181 vss 3.13114e-17
C311 s_1_180 vss 3.13114e-17
C312 s_1_182 vss 3.13114e-17
C313 s_1_181 vss 3.13114e-17
C314 s_1_183 vss 3.13114e-17
C315 s_1_182 vss 3.13114e-17
C316 s_1_184 vss 3.13114e-17
C317 s_1_183 vss 3.13114e-17
C318 s_1_185 vss 3.13114e-17
C319 s_1_184 vss 3.13114e-17
C320 s_1_186 vss 3.13114e-17
C321 s_1_185 vss 3.13114e-17
C322 s_1_187 vss 3.13114e-17
C323 s_1_186 vss 3.13114e-17
C324 s_1_188 vss 3.13114e-17
C325 s_1_187 vss 3.13114e-17
C326 s_1_189 vss 3.13114e-17
C327 s_1_188 vss 3.13114e-17
C328 s_1_190 vss 3.13114e-17
C329 s_1_189 vss 3.13114e-17
C330 s_1_191 vss 3.13114e-17
C331 s_1_190 vss 3.13114e-17
C332 s_1_192 vss 3.13114e-17
C333 s_1_191 vss 3.13114e-17
C334 s_1_193 vss 3.13114e-17
C335 s_1_192 vss 3.13114e-17
C336 s_1_194 vss 3.13114e-17
C337 s_1_193 vss 3.13114e-17
C338 s_1_195 vss 3.13114e-17
C339 s_1_194 vss 3.13114e-17
C340 s_1_196 vss 3.13114e-17
C341 s_1_195 vss 3.13114e-17
C342 s_1_197 vss 3.13114e-17
C343 s_1_196 vss 3.13114e-17
C344 s_1_198 vss 3.13114e-17
C345 s_1_197 vss 3.13114e-17
C346 s_1_199 vss 3.13114e-17
C347 s_1_198 vss 3.13114e-17
C348 s_1_200 vss 1.40901e-17
C349 s_1_199 vss 1.40901e-17
C350 s_1_201 vss 3.60081e-16
C351 s_1_349 vss 3.60081e-16
C352 s_1_202 vss 3.13114e-17
C353 s_1_201 vss 3.13114e-17
C354 s_1_203 vss 3.13114e-17
C355 s_1_202 vss 3.13114e-17
C356 s_1_204 vss 3.13114e-17
C357 s_1_203 vss 3.13114e-17
C358 s_1_205 vss 3.13114e-17
C359 s_1_204 vss 3.13114e-17
C360 s_1_206 vss 3.13114e-17
C361 s_1_205 vss 3.13114e-17
C362 s_1_207 vss 3.13114e-17
C363 s_1_206 vss 3.13114e-17
C364 s_1_208 vss 3.13114e-17
C365 s_1_207 vss 3.13114e-17
C366 s_1_209 vss 2.42663e-16
C367 s_1_208 vss 2.42663e-16
C368 s_1_210 vss 3.13114e-17
C369 s_1_209 vss 3.13114e-17
C370 s_1_211 vss 3.13114e-17
C371 s_1_210 vss 3.13114e-17
C372 s_1_212 vss 3.13114e-17
C373 s_1_211 vss 3.13114e-17
C374 s_1_213 vss 3.13114e-17
C375 s_1_212 vss 3.13114e-17
C376 s_1_214 vss 3.13114e-17
C377 s_1_213 vss 3.13114e-17
C378 s_1_215 vss 3.13114e-17
C379 s_1_214 vss 3.13114e-17
C380 s_1_216 vss 3.13114e-17
C381 s_1_215 vss 3.13114e-17
C382 s_1_217 vss 3.13114e-17
C383 s_1_216 vss 3.13114e-17
C384 s_1_218 vss 3.13114e-17
C385 s_1_217 vss 3.13114e-17
C386 s_1_219 vss 3.13114e-17
C387 s_1_218 vss 3.13114e-17
C388 s_1_220 vss 3.13114e-17
C389 s_1_219 vss 3.13114e-17
C390 s_1_221 vss 3.13114e-17
C391 s_1_220 vss 3.13114e-17
C392 s_1_222 vss 3.13114e-17
C393 s_1_221 vss 3.13114e-17
C394 s_1_223 vss 3.13114e-17
C395 s_1_222 vss 3.13114e-17
C396 s_1_224 vss 3.13114e-17
C397 s_1_223 vss 3.13114e-17
C398 s_1_225 vss 3.13114e-17
C399 s_1_224 vss 3.13114e-17
C400 s_1_226 vss 3.13114e-17
C401 s_1_225 vss 3.13114e-17
C402 s_1_227 vss 3.13114e-17
C403 s_1_226 vss 3.13114e-17
C404 s_1_228 vss 3.13114e-17
C405 s_1_227 vss 3.13114e-17
C406 s_1_229 vss 1.40901e-17
C407 s_1_228 vss 1.40901e-17
C408 s_1_230 vss 3.60081e-16
C409 s_1_349 vss 3.60081e-16
C410 s_1_231 vss 3.13114e-17
C411 s_1_230 vss 3.13114e-17
C412 s_1_232 vss 3.13114e-17
C413 s_1_231 vss 3.13114e-17
C414 s_1_233 vss 3.13114e-17
C415 s_1_232 vss 3.13114e-17
C416 s_1_234 vss 3.13114e-17
C417 s_1_233 vss 3.13114e-17
C418 s_1_235 vss 3.13114e-17
C419 s_1_234 vss 3.13114e-17
C420 s_1_236 vss 3.13114e-17
C421 s_1_235 vss 3.13114e-17
C422 s_1_237 vss 3.13114e-17
C423 s_1_236 vss 3.13114e-17
C424 s_1_238 vss 2.42663e-16
C425 s_1_237 vss 2.42663e-16
C426 s_1_239 vss 3.13114e-17
C427 s_1_238 vss 3.13114e-17
C428 s_1_240 vss 3.13114e-17
C429 s_1_239 vss 3.13114e-17
C430 s_1_241 vss 3.13114e-17
C431 s_1_240 vss 3.13114e-17
C432 s_1_242 vss 3.13114e-17
C433 s_1_241 vss 3.13114e-17
C434 s_1_243 vss 3.13114e-17
C435 s_1_242 vss 3.13114e-17
C436 s_1_244 vss 3.13114e-17
C437 s_1_243 vss 3.13114e-17
C438 s_1_245 vss 3.13114e-17
C439 s_1_244 vss 3.13114e-17
C440 s_1_246 vss 3.13114e-17
C441 s_1_245 vss 3.13114e-17
C442 s_1_247 vss 3.13114e-17
C443 s_1_246 vss 3.13114e-17
C444 s_1_248 vss 3.13114e-17
C445 s_1_247 vss 3.13114e-17
C446 s_1_249 vss 3.13114e-17
C447 s_1_248 vss 3.13114e-17
C448 s_1_250 vss 3.13114e-17
C449 s_1_249 vss 3.13114e-17
C450 s_1_251 vss 3.13114e-17
C451 s_1_250 vss 3.13114e-17
C452 s_1_252 vss 3.13114e-17
C453 s_1_251 vss 3.13114e-17
C454 s_1_253 vss 3.13114e-17
C455 s_1_252 vss 3.13114e-17
C456 s_1_254 vss 3.13114e-17
C457 s_1_253 vss 3.13114e-17
C458 s_1_255 vss 3.13114e-17
C459 s_1_254 vss 3.13114e-17
C460 s_1_256 vss 3.13114e-17
C461 s_1_255 vss 3.13114e-17
C462 s_1_257 vss 3.13114e-17
C463 s_1_256 vss 3.13114e-17
C464 s_1_258 vss 1.40901e-17
C465 s_1_257 vss 1.40901e-17
C466 s_1_259 vss 3.60081e-16
C467 s_1_349 vss 3.60081e-16
C468 s_1_260 vss 3.13114e-17
C469 s_1_259 vss 3.13114e-17
C470 s_1_261 vss 3.13114e-17
C471 s_1_260 vss 3.13114e-17
C472 s_1_262 vss 3.13114e-17
C473 s_1_261 vss 3.13114e-17
C474 s_1_263 vss 3.13114e-17
C475 s_1_262 vss 3.13114e-17
C476 s_1_264 vss 3.13114e-17
C477 s_1_263 vss 3.13114e-17
C478 s_1_265 vss 3.13114e-17
C479 s_1_264 vss 3.13114e-17
C480 s_1_266 vss 3.13114e-17
C481 s_1_265 vss 3.13114e-17
C482 s_1_267 vss 2.42663e-16
C483 s_1_266 vss 2.42663e-16
C484 s_1_268 vss 3.13114e-17
C485 s_1_267 vss 3.13114e-17
C486 s_1_269 vss 3.13114e-17
C487 s_1_268 vss 3.13114e-17
C488 s_1_270 vss 3.13114e-17
C489 s_1_269 vss 3.13114e-17
C490 s_1_271 vss 3.13114e-17
C491 s_1_270 vss 3.13114e-17
C492 s_1_272 vss 3.13114e-17
C493 s_1_271 vss 3.13114e-17
C494 s_1_273 vss 3.13114e-17
C495 s_1_272 vss 3.13114e-17
C496 s_1_274 vss 3.13114e-17
C497 s_1_273 vss 3.13114e-17
C498 s_1_275 vss 3.13114e-17
C499 s_1_274 vss 3.13114e-17
C500 s_1_276 vss 3.13114e-17
C501 s_1_275 vss 3.13114e-17
C502 s_1_277 vss 3.13114e-17
C503 s_1_276 vss 3.13114e-17
C504 s_1_278 vss 3.13114e-17
C505 s_1_277 vss 3.13114e-17
C506 s_1_279 vss 3.13114e-17
C507 s_1_278 vss 3.13114e-17
C508 s_1_280 vss 3.13114e-17
C509 s_1_279 vss 3.13114e-17
C510 s_1_281 vss 3.13114e-17
C511 s_1_280 vss 3.13114e-17
C512 s_1_282 vss 3.13114e-17
C513 s_1_281 vss 3.13114e-17
C514 s_1_283 vss 3.13114e-17
C515 s_1_282 vss 3.13114e-17
C516 s_1_284 vss 3.13114e-17
C517 s_1_283 vss 3.13114e-17
C518 s_1_285 vss 3.13114e-17
C519 s_1_284 vss 3.13114e-17
C520 s_1_286 vss 3.13114e-17
C521 s_1_285 vss 3.13114e-17
C522 s_1_287 vss 1.40901e-17
C523 s_1_286 vss 1.40901e-17
C524 s_1_288 vss 1.40901e-16
C525 s_1_346 vss 1.40901e-16
C526 s_1_289 vss 3.13114e-17
C527 s_1_288 vss 3.13114e-17
C528 s_1_290 vss 3.13114e-17
C529 s_1_289 vss 3.13114e-17
C530 s_1_291 vss 3.13114e-17
C531 s_1_290 vss 3.13114e-17
C532 s_1_292 vss 3.13114e-17
C533 s_1_291 vss 3.13114e-17
C534 s_1_293 vss 3.13114e-17
C535 s_1_292 vss 3.13114e-17
C536 s_1_294 vss 3.13114e-17
C537 s_1_293 vss 3.13114e-17
C538 s_1_295 vss 3.13114e-17
C539 s_1_294 vss 3.13114e-17
C540 s_1_296 vss 2.42663e-16
C541 s_1_295 vss 2.42663e-16
C542 s_1_297 vss 3.13114e-17
C543 s_1_296 vss 3.13114e-17
C544 s_1_298 vss 3.13114e-17
C545 s_1_297 vss 3.13114e-17
C546 s_1_299 vss 3.13114e-17
C547 s_1_298 vss 3.13114e-17
C548 s_1_300 vss 3.13114e-17
C549 s_1_299 vss 3.13114e-17
C550 s_1_301 vss 3.13114e-17
C551 s_1_300 vss 3.13114e-17
C552 s_1_302 vss 3.13114e-17
C553 s_1_301 vss 3.13114e-17
C554 s_1_303 vss 3.13114e-17
C555 s_1_302 vss 3.13114e-17
C556 s_1_304 vss 3.13114e-17
C557 s_1_303 vss 3.13114e-17
C558 s_1_305 vss 3.13114e-17
C559 s_1_304 vss 3.13114e-17
C560 s_1_306 vss 3.13114e-17
C561 s_1_305 vss 3.13114e-17
C562 s_1_307 vss 3.13114e-17
C563 s_1_306 vss 3.13114e-17
C564 s_1_308 vss 3.13114e-17
C565 s_1_307 vss 3.13114e-17
C566 s_1_309 vss 3.13114e-17
C567 s_1_308 vss 3.13114e-17
C568 s_1_310 vss 3.13114e-17
C569 s_1_309 vss 3.13114e-17
C570 s_1_311 vss 3.13114e-17
C571 s_1_310 vss 3.13114e-17
C572 s_1_312 vss 3.13114e-17
C573 s_1_311 vss 3.13114e-17
C574 s_1_313 vss 3.13114e-17
C575 s_1_312 vss 3.13114e-17
C576 s_1_314 vss 3.13114e-17
C577 s_1_313 vss 3.13114e-17
C578 s_1_315 vss 3.13114e-17
C579 s_1_314 vss 3.13114e-17
C580 s_1_316 vss 1.40901e-17
C581 s_1_315 vss 1.40901e-17
C582 s_1_317 vss 1.40901e-16
C583 s_1_348 vss 1.40901e-16
C584 s_1_318 vss 3.13114e-17
C585 s_1_317 vss 3.13114e-17
C586 s_1_319 vss 3.13114e-17
C587 s_1_318 vss 3.13114e-17
C588 s_1_320 vss 3.13114e-17
C589 s_1_319 vss 3.13114e-17
C590 s_1_321 vss 3.13114e-17
C591 s_1_320 vss 3.13114e-17
C592 s_1_322 vss 3.13114e-17
C593 s_1_321 vss 3.13114e-17
C594 s_1_323 vss 3.13114e-17
C595 s_1_322 vss 3.13114e-17
C596 s_1_324 vss 3.13114e-17
C597 s_1_323 vss 3.13114e-17
C598 s_1_325 vss 2.42663e-16
C599 s_1_324 vss 2.42663e-16
C600 s_1_326 vss 3.13114e-17
C601 s_1_325 vss 3.13114e-17
C602 s_1_327 vss 3.13114e-17
C603 s_1_326 vss 3.13114e-17
C604 s_1_328 vss 3.13114e-17
C605 s_1_327 vss 3.13114e-17
C606 s_1_329 vss 3.13114e-17
C607 s_1_328 vss 3.13114e-17
C608 s_1_330 vss 3.13114e-17
C609 s_1_329 vss 3.13114e-17
C610 s_1_331 vss 3.13114e-17
C611 s_1_330 vss 3.13114e-17
C612 s_1_332 vss 3.13114e-17
C613 s_1_331 vss 3.13114e-17
C614 s_1_333 vss 3.13114e-17
C615 s_1_332 vss 3.13114e-17
C616 s_1_334 vss 3.13114e-17
C617 s_1_333 vss 3.13114e-17
C618 s_1_335 vss 3.13114e-17
C619 s_1_334 vss 3.13114e-17
C620 s_1_336 vss 3.13114e-17
C621 s_1_335 vss 3.13114e-17
C622 s_1_337 vss 3.13114e-17
C623 s_1_336 vss 3.13114e-17
C624 s_1_338 vss 3.13114e-17
C625 s_1_337 vss 3.13114e-17
C626 s_1_339 vss 3.13114e-17
C627 s_1_338 vss 3.13114e-17
C628 s_1_340 vss 3.13114e-17
C629 s_1_339 vss 3.13114e-17
C630 s_1_341 vss 3.13114e-17
C631 s_1_340 vss 3.13114e-17
C632 s_1_342 vss 3.13114e-17
C633 s_1_341 vss 3.13114e-17
C634 s_1_343 vss 3.13114e-17
C635 s_1_342 vss 3.13114e-17
C636 s_1_344 vss 3.13114e-17
C637 s_1_343 vss 3.13114e-17
C638 s_1_345 vss 1.40901e-17
C639 s_1_344 vss 1.40901e-17
C640 s_1_347 vss 2.95333e-17
C641 s_1_346 vss 2.95333e-17
C642 s_1_348 vss 3.71708e-16
C643 s_1_347 vss 3.71708e-16
C644 s_1_349 vss 2.15831e-15
C645 s_1_348 vss 2.15831e-15
C646 s_1_352 vss 2.15831e-15
C647 s_1_349 vss 2.15831e-15
C648 s_1_350 vss 3.71708e-16
C649 s_1_352 vss 3.71708e-16
C650 s_1_351 vss 2.95333e-17
C651 s_1_350 vss 2.95333e-17
C652 s_1_353 vss 1.40901e-16
C653 s_1_352 vss 1.40901e-16
C654 s_1_354 vss 3.13114e-17
C655 s_1_353 vss 3.13114e-17
C656 s_1_355 vss 3.13114e-17
C657 s_1_354 vss 3.13114e-17
C658 s_1_356 vss 3.13114e-17
C659 s_1_355 vss 3.13114e-17
C660 s_1_357 vss 3.13114e-17
C661 s_1_356 vss 3.13114e-17
C662 s_1_358 vss 3.13114e-17
C663 s_1_357 vss 3.13114e-17
C664 s_1_359 vss 3.13114e-17
C665 s_1_358 vss 3.13114e-17
C666 s_1_360 vss 3.13114e-17
C667 s_1_359 vss 3.13114e-17
C668 s_1_361 vss 2.42663e-16
C669 s_1_360 vss 2.42663e-16
C670 s_1_362 vss 3.13114e-17
C671 s_1_361 vss 3.13114e-17
C672 s_1_363 vss 3.13114e-17
C673 s_1_362 vss 3.13114e-17
C674 s_1_364 vss 3.13114e-17
C675 s_1_363 vss 3.13114e-17
C676 s_1_365 vss 3.13114e-17
C677 s_1_364 vss 3.13114e-17
C678 s_1_366 vss 3.13114e-17
C679 s_1_365 vss 3.13114e-17
C680 s_1_367 vss 3.13114e-17
C681 s_1_366 vss 3.13114e-17
C682 s_1_368 vss 3.13114e-17
C683 s_1_367 vss 3.13114e-17
C684 s_1_369 vss 3.13114e-17
C685 s_1_368 vss 3.13114e-17
C686 s_1_370 vss 3.13114e-17
C687 s_1_369 vss 3.13114e-17
C688 s_1_371 vss 3.13114e-17
C689 s_1_370 vss 3.13114e-17
C690 s_1_372 vss 3.13114e-17
C691 s_1_371 vss 3.13114e-17
C692 s_1_373 vss 3.13114e-17
C693 s_1_372 vss 3.13114e-17
C694 s_1_374 vss 3.13114e-17
C695 s_1_373 vss 3.13114e-17
C696 s_1_375 vss 3.13114e-17
C697 s_1_374 vss 3.13114e-17
C698 s_1_376 vss 3.13114e-17
C699 s_1_375 vss 3.13114e-17
C700 s_1_377 vss 3.13114e-17
C701 s_1_376 vss 3.13114e-17
C702 s_1_378 vss 3.13114e-17
C703 s_1_377 vss 3.13114e-17
C704 s_1_379 vss 3.13114e-17
C705 s_1_378 vss 3.13114e-17
C706 s_1_380 vss 3.13114e-17
C707 s_1_379 vss 3.13114e-17
C708 s_1_381 vss 1.40901e-17
C709 s_1_380 vss 1.40901e-17

R40_1 s_0_1 s_0_379 0.001
R40_2 s_0_1 s_0_380 0.001
R40_3 s_0_54 s_0_2 0.001
R40_4 s_0_53 s_0_2 0.001
R40_5 s_0_82 s_0_3 0.001
R40_6 s_0_83 s_0_3 0.001
R40_7 s_0_141 s_0_4 0.001
R40_8 s_0_140 s_0_4 0.001
R40_9 s_0_111 s_0_5 0.001
R40_10 s_0_112 s_0_5 0.001
R40_11 s_0_169 s_0_6 0.001
R40_12 s_0_170 s_0_6 0.001
R40_13 s_0_228 s_0_7 0.001
R40_14 s_0_227 s_0_7 0.001
R40_15 s_0_199 s_0_8 0.001
R40_16 s_0_198 s_0_8 0.001
R40_17 s_0_256 s_0_9 0.001
R40_18 s_0_257 s_0_9 0.001
R40_19 s_0_286 s_0_10 0.001
R40_20 s_0_285 s_0_10 0.001
R40_21 s_0_315 s_0_11 0.001
R40_22 s_0_314 s_0_11 0.001
R40_23 s_0_344 s_0_12 0.001
R40_24 s_0_343 s_0_12 0.001
R40_25 s_0_1 s_0_378 0.001
R40_26 s_0_52 s_0_2 0.001
R40_27 s_0_81 s_0_3 0.001
R40_28 s_0_139 s_0_4 0.001
R40_29 s_0_110 s_0_5 0.001
R40_30 s_0_168 s_0_6 0.001
R40_31 s_0_226 s_0_7 0.001
R40_32 s_0_197 s_0_8 0.001
R40_33 s_0_255 s_0_9 0.001
R40_34 s_0_284 s_0_10 0.001
R40_35 s_0_313 s_0_11 0.001
R40_36 s_0_342 s_0_12 0.001
R40_37 s_0_1 s_0_377 0.001
R40_38 s_0_51 s_0_2 0.001
R40_39 s_0_80 s_0_3 0.001
R40_40 s_0_138 s_0_4 0.001
R40_41 s_0_109 s_0_5 0.001
R40_42 s_0_167 s_0_6 0.001
R40_43 s_0_225 s_0_7 0.001
R40_44 s_0_196 s_0_8 0.001
R40_45 s_0_254 s_0_9 0.001
R40_46 s_0_283 s_0_10 0.001
R40_47 s_0_312 s_0_11 0.001
R40_48 s_0_341 s_0_12 0.001
R40_49 s_0_1 s_0_375 0.001
R40_50 s_0_1 s_0_376 0.001
R40_51 s_0_49 s_0_2 0.001
R40_52 s_0_50 s_0_2 0.001
R40_53 s_0_78 s_0_3 0.001
R40_54 s_0_79 s_0_3 0.001
R40_55 s_0_136 s_0_4 0.001
R40_56 s_0_137 s_0_4 0.001
R40_57 s_0_107 s_0_5 0.001
R40_58 s_0_108 s_0_5 0.001
R40_59 s_0_165 s_0_6 0.001
R40_60 s_0_166 s_0_6 0.001
R40_61 s_0_223 s_0_7 0.001
R40_62 s_0_224 s_0_7 0.001
R40_63 s_0_194 s_0_8 0.001
R40_64 s_0_195 s_0_8 0.001
R40_65 s_0_252 s_0_9 0.001
R40_66 s_0_253 s_0_9 0.001
R40_67 s_0_281 s_0_10 0.001
R40_68 s_0_282 s_0_10 0.001
R40_69 s_0_310 s_0_11 0.001
R40_70 s_0_311 s_0_11 0.001
R40_71 s_0_340 s_0_12 0.001
R40_72 s_0_339 s_0_12 0.001
R40_73 s_0_1 s_0_374 0.001
R40_74 s_0_48 s_0_2 0.001
R40_75 s_0_77 s_0_3 0.001
R40_76 s_0_135 s_0_4 0.001
R40_77 s_0_106 s_0_5 0.001
R40_78 s_0_164 s_0_6 0.001
R40_79 s_0_222 s_0_7 0.001
R40_80 s_0_193 s_0_8 0.001
R40_81 s_0_251 s_0_9 0.001
R40_82 s_0_280 s_0_10 0.001
R40_83 s_0_309 s_0_11 0.001
R40_84 s_0_338 s_0_12 0.001
R40_85 s_0_1 s_0_372 0.001
R40_86 s_0_1 s_0_373 0.001
R40_87 s_0_46 s_0_2 0.001
R40_88 s_0_47 s_0_2 0.001
R40_89 s_0_75 s_0_3 0.001
R40_90 s_0_76 s_0_3 0.001
R40_91 s_0_133 s_0_4 0.001
R40_92 s_0_134 s_0_4 0.001
R40_93 s_0_104 s_0_5 0.001
R40_94 s_0_105 s_0_5 0.001
R40_95 s_0_162 s_0_6 0.001
R40_96 s_0_163 s_0_6 0.001
R40_97 s_0_220 s_0_7 0.001
R40_98 s_0_221 s_0_7 0.001
R40_99 s_0_191 s_0_8 0.001
R40_100 s_0_192 s_0_8 0.001
R40_101 s_0_250 s_0_9 0.001
R40_102 s_0_249 s_0_9 0.001
R40_103 s_0_278 s_0_10 0.001
R40_104 s_0_279 s_0_10 0.001
R40_105 s_0_307 s_0_11 0.001
R40_106 s_0_308 s_0_11 0.001
R40_107 s_0_336 s_0_12 0.001
R40_108 s_0_337 s_0_12 0.001
R40_109 s_0_1 s_0_371 0.001
R40_110 s_0_45 s_0_2 0.001
R40_111 s_0_74 s_0_3 0.001
R40_112 s_0_132 s_0_4 0.001
R40_113 s_0_103 s_0_5 0.001
R40_114 s_0_161 s_0_6 0.001
R40_115 s_0_219 s_0_7 0.001
R40_116 s_0_190 s_0_8 0.001
R40_117 s_0_248 s_0_9 0.001
R40_118 s_0_277 s_0_10 0.001
R40_119 s_0_306 s_0_11 0.001
R40_120 s_0_335 s_0_12 0.001
R40_121 s_0_1 s_0_370 0.001
R40_122 s_0_44 s_0_2 0.001
R40_123 s_0_73 s_0_3 0.001
R40_124 s_0_131 s_0_4 0.001
R40_125 s_0_102 s_0_5 0.001
R40_126 s_0_160 s_0_6 0.001
R40_127 s_0_218 s_0_7 0.001
R40_128 s_0_189 s_0_8 0.001
R40_129 s_0_247 s_0_9 0.001
R40_130 s_0_276 s_0_10 0.001
R40_131 s_0_305 s_0_11 0.001
R40_132 s_0_334 s_0_12 0.001
R40_133 s_0_1 s_0_369 0.001
R40_134 s_0_1 s_0_368 0.001
R40_135 s_0_43 s_0_2 0.001
R40_136 s_0_42 s_0_2 0.001
R40_137 s_0_72 s_0_3 0.001
R40_138 s_0_71 s_0_3 0.001
R40_139 s_0_130 s_0_4 0.001
R40_140 s_0_129 s_0_4 0.001
R40_141 s_0_101 s_0_5 0.001
R40_142 s_0_100 s_0_5 0.001
R40_143 s_0_159 s_0_6 0.001
R40_144 s_0_158 s_0_6 0.001
R40_145 s_0_217 s_0_7 0.001
R40_146 s_0_216 s_0_7 0.001
R40_147 s_0_188 s_0_8 0.001
R40_148 s_0_187 s_0_8 0.001
R40_149 s_0_246 s_0_9 0.001
R40_150 s_0_245 s_0_9 0.001
R40_151 s_0_275 s_0_10 0.001
R40_152 s_0_274 s_0_10 0.001
R40_153 s_0_304 s_0_11 0.001
R40_154 s_0_303 s_0_11 0.001
R40_155 s_0_333 s_0_12 0.001
R40_156 s_0_332 s_0_12 0.001
R40_157 s_0_1 s_0_367 0.001
R40_158 s_0_41 s_0_2 0.001
R40_159 s_0_70 s_0_3 0.001
R40_160 s_0_128 s_0_4 0.001
R40_161 s_0_99 s_0_5 0.001
R40_162 s_0_157 s_0_6 0.001
R40_163 s_0_215 s_0_7 0.001
R40_164 s_0_186 s_0_8 0.001
R40_165 s_0_244 s_0_9 0.001
R40_166 s_0_273 s_0_10 0.001
R40_167 s_0_302 s_0_11 0.001
R40_168 s_0_331 s_0_12 0.001
R40_169 s_0_1 s_0_366 0.001
R40_170 s_0_1 s_0_365 0.001
R40_171 s_0_40 s_0_2 0.001
R40_172 s_0_39 s_0_2 0.001
R40_173 s_0_69 s_0_3 0.001
R40_174 s_0_68 s_0_3 0.001
R40_175 s_0_126 s_0_4 0.001
R40_176 s_0_127 s_0_4 0.001
R40_177 s_0_98 s_0_5 0.001
R40_178 s_0_97 s_0_5 0.001
R40_179 s_0_156 s_0_6 0.001
R40_180 s_0_155 s_0_6 0.001
R40_181 s_0_213 s_0_7 0.001
R40_182 s_0_214 s_0_7 0.001
R40_183 s_0_184 s_0_8 0.001
R40_184 s_0_185 s_0_8 0.001
R40_185 s_0_243 s_0_9 0.001
R40_186 s_0_242 s_0_9 0.001
R40_187 s_0_272 s_0_10 0.001
R40_188 s_0_271 s_0_10 0.001
R40_189 s_0_301 s_0_11 0.001
R40_190 s_0_300 s_0_11 0.001
R40_191 s_0_330 s_0_12 0.001
R40_192 s_0_329 s_0_12 0.001
R40_193 s_0_1 s_0_364 0.001
R40_194 s_0_38 s_0_2 0.001
R40_195 s_0_67 s_0_3 0.001
R40_196 s_0_125 s_0_4 0.001
R40_197 s_0_96 s_0_5 0.001
R40_198 s_0_154 s_0_6 0.001
R40_199 s_0_212 s_0_7 0.001
R40_200 s_0_183 s_0_8 0.001
R40_201 s_0_241 s_0_9 0.001
R40_202 s_0_270 s_0_10 0.001
R40_203 s_0_299 s_0_11 0.001
R40_204 s_0_328 s_0_12 0.001
R40_205 s_0_1 s_0_363 0.001
R40_206 s_0_37 s_0_2 0.001
R40_207 s_0_66 s_0_3 0.001
R40_208 s_0_124 s_0_4 0.001
R40_209 s_0_95 s_0_5 0.001
R40_210 s_0_153 s_0_6 0.001
R40_211 s_0_211 s_0_7 0.001
R40_212 s_0_182 s_0_8 0.001
R40_213 s_0_240 s_0_9 0.001
R40_214 s_0_269 s_0_10 0.001
R40_215 s_0_298 s_0_11 0.001
R40_216 s_0_327 s_0_12 0.001
R40_217 s_0_1 s_0_362 0.001
R40_218 s_0_1 s_0_361 0.001
R40_219 s_0_35 s_0_2 0.001
R40_220 s_0_36 s_0_2 0.001
R40_221 s_0_64 s_0_3 0.001
R40_222 s_0_65 s_0_3 0.001
R40_223 s_0_122 s_0_4 0.001
R40_224 s_0_123 s_0_4 0.001
R40_225 s_0_93 s_0_5 0.001
R40_226 s_0_94 s_0_5 0.001
R40_227 s_0_151 s_0_6 0.001
R40_228 s_0_152 s_0_6 0.001
R40_229 s_0_209 s_0_7 0.001
R40_230 s_0_210 s_0_7 0.001
R40_231 s_0_180 s_0_8 0.001
R40_232 s_0_181 s_0_8 0.001
R40_233 s_0_239 s_0_9 0.001
R40_234 s_0_238 s_0_9 0.001
R40_235 s_0_267 s_0_10 0.001
R40_236 s_0_268 s_0_10 0.001
R40_237 s_0_296 s_0_11 0.001
R40_238 s_0_297 s_0_11 0.001
R40_239 s_0_325 s_0_12 0.001
R40_240 s_0_326 s_0_12 0.001
R40_241 s_0_360 s_0_13 0.001
R40_242 s_0_359 s_0_13 0.001
R40_243 s_0_33 s_0_14 0.001
R40_244 s_0_34 s_0_14 0.001
R40_245 s_0_62 s_0_15 0.001
R40_246 s_0_63 s_0_15 0.001
R40_247 s_0_121 s_0_16 0.001
R40_248 s_0_120 s_0_16 0.001
R40_249 s_0_91 s_0_17 0.001
R40_250 s_0_92 s_0_17 0.001
R40_251 s_0_149 s_0_18 0.001
R40_252 s_0_150 s_0_18 0.001
R40_253 s_0_208 s_0_19 0.001
R40_254 s_0_207 s_0_19 0.001
R40_255 s_0_178 s_0_20 0.001
R40_256 s_0_179 s_0_20 0.001
R40_257 s_0_237 s_0_21 0.001
R40_258 s_0_236 s_0_21 0.001
R40_259 s_0_265 s_0_22 0.001
R40_260 s_0_266 s_0_22 0.001
R40_261 s_0_294 s_0_23 0.001
R40_262 s_0_295 s_0_23 0.001
R40_263 s_0_323 s_0_24 0.001
R40_264 s_0_324 s_0_24 0.001
R40_265 s_0_358 s_0_13 0.001
R40_266 s_0_32 s_0_14 0.001
R40_267 s_0_61 s_0_15 0.001
R40_268 s_0_119 s_0_16 0.001
R40_269 s_0_90 s_0_17 0.001
R40_270 s_0_148 s_0_18 0.001
R40_271 s_0_206 s_0_19 0.001
R40_272 s_0_177 s_0_20 0.001
R40_273 s_0_235 s_0_21 0.001
R40_274 s_0_264 s_0_22 0.001
R40_275 s_0_293 s_0_23 0.001
R40_276 s_0_322 s_0_24 0.001
R40_277 s_0_357 s_0_13 0.001
R40_278 s_0_31 s_0_14 0.001
R40_279 s_0_60 s_0_15 0.001
R40_280 s_0_118 s_0_16 0.001
R40_281 s_0_89 s_0_17 0.001
R40_282 s_0_147 s_0_18 0.001
R40_283 s_0_205 s_0_19 0.001
R40_284 s_0_176 s_0_20 0.001
R40_285 s_0_234 s_0_21 0.001
R40_286 s_0_263 s_0_22 0.001
R40_287 s_0_292 s_0_23 0.001
R40_288 s_0_321 s_0_24 0.001
R40_289 s_0_356 s_0_13 0.001
R40_290 s_0_355 s_0_13 0.001
R40_291 s_0_30 s_0_14 0.001
R40_292 s_0_29 s_0_14 0.001
R40_293 s_0_59 s_0_15 0.001
R40_294 s_0_58 s_0_15 0.001
R40_295 s_0_117 s_0_16 0.001
R40_296 s_0_116 s_0_16 0.001
R40_297 s_0_88 s_0_17 0.001
R40_298 s_0_87 s_0_17 0.001
R40_299 s_0_146 s_0_18 0.001
R40_300 s_0_145 s_0_18 0.001
R40_301 s_0_203 s_0_19 0.001
R40_302 s_0_204 s_0_19 0.001
R40_303 s_0_175 s_0_20 0.001
R40_304 s_0_174 s_0_20 0.001
R40_305 s_0_233 s_0_21 0.001
R40_306 s_0_232 s_0_21 0.001
R40_307 s_0_262 s_0_22 0.001
R40_308 s_0_261 s_0_22 0.001
R40_309 s_0_291 s_0_23 0.001
R40_310 s_0_290 s_0_23 0.001
R40_311 s_0_320 s_0_24 0.001
R40_312 s_0_319 s_0_24 0.001
R40_313 s_0_354 s_0_13 0.001
R40_314 s_0_28 s_0_14 0.001
R40_315 s_0_57 s_0_15 0.001
R40_316 s_0_115 s_0_16 0.001
R40_317 s_0_86 s_0_17 0.001
R40_318 s_0_144 s_0_18 0.001
R40_319 s_0_202 s_0_19 0.001
R40_320 s_0_173 s_0_20 0.001
R40_321 s_0_231 s_0_21 0.001
R40_322 s_0_260 s_0_22 0.001
R40_323 s_0_289 s_0_23 0.001
R40_324 s_0_318 s_0_24 0.001
R40_325 s_0_353 s_0_13 0.001
R40_326 s_0_27 s_0_14 0.001
R40_327 s_0_56 s_0_15 0.001
R40_328 s_0_114 s_0_16 0.001
R40_329 s_0_85 s_0_17 0.001
R40_330 s_0_143 s_0_18 0.001
R40_331 s_0_201 s_0_19 0.001
R40_332 s_0_172 s_0_20 0.001
R40_333 s_0_230 s_0_21 0.001
R40_334 s_0_259 s_0_22 0.001
R40_335 s_0_288 s_0_23 0.001
R40_336 s_0_317 s_0_24 0.001
R40_337 s_0 s_0_25 0.001
R40_338 s_0_349 s_0 0.108
R40_339 s_0_27 s_0_350 0.54
R40_340 s_0_28 s_0_27 0.108
R40_341 s_0_29 s_0_28 0.108
R40_342 s_0_30 s_0_29 0.108
R40_343 s_0_31 s_0_30 0.108
R40_344 s_0_32 s_0_31 0.108
R40_345 s_0_33 s_0_32 0.108
R40_346 s_0_34 s_0_33 0.108
R40_347 s_0_35 s_0_34 0.864
R40_348 s_0_36 s_0_35 0.108
R40_349 s_0_37 s_0_36 0.108
R40_350 s_0_38 s_0_37 0.108
R40_351 s_0_39 s_0_38 0.108
R40_352 s_0_40 s_0_39 0.108
R40_353 s_0_41 s_0_40 0.108
R40_354 s_0_42 s_0_41 0.108
R40_355 s_0_43 s_0_42 0.108
R40_356 s_0_44 s_0_43 0.108
R40_357 s_0_45 s_0_44 0.108
R40_358 s_0_46 s_0_45 0.108
R40_359 s_0_47 s_0_46 0.108
R40_360 s_0_48 s_0_47 0.108
R40_361 s_0_49 s_0_48 0.108
R40_362 s_0_50 s_0_49 0.108
R40_363 s_0_51 s_0_50 0.108
R40_364 s_0_52 s_0_51 0.108
R40_365 s_0_53 s_0_52 0.108
R40_366 s_0_54 s_0_53 0.108
R40_367 s_0_55 s_0_54 0.001
R40_368 s_0_56 s_0_349 1.296
R40_369 s_0_57 s_0_56 0.108
R40_370 s_0_58 s_0_57 0.108
R40_371 s_0_59 s_0_58 0.108
R40_372 s_0_60 s_0_59 0.108
R40_373 s_0_61 s_0_60 0.108
R40_374 s_0_62 s_0_61 0.108
R40_375 s_0_63 s_0_62 0.108
R40_376 s_0_64 s_0_63 0.864
R40_377 s_0_65 s_0_64 0.108
R40_378 s_0_66 s_0_65 0.108
R40_379 s_0_67 s_0_66 0.108
R40_380 s_0_68 s_0_67 0.108
R40_381 s_0_69 s_0_68 0.108
R40_382 s_0_70 s_0_69 0.108
R40_383 s_0_71 s_0_70 0.108
R40_384 s_0_72 s_0_71 0.108
R40_385 s_0_73 s_0_72 0.108
R40_386 s_0_74 s_0_73 0.108
R40_387 s_0_75 s_0_74 0.108
R40_388 s_0_76 s_0_75 0.108
R40_389 s_0_77 s_0_76 0.108
R40_390 s_0_78 s_0_77 0.108
R40_391 s_0_79 s_0_78 0.108
R40_392 s_0_80 s_0_79 0.108
R40_393 s_0_81 s_0_80 0.108
R40_394 s_0_82 s_0_81 0.108
R40_395 s_0_83 s_0_82 0.108
R40_396 s_0_84 s_0_83 0.001
R40_397 s_0_85 s_0_349 1.296
R40_398 s_0_86 s_0_85 0.108
R40_399 s_0_87 s_0_86 0.108
R40_400 s_0_88 s_0_87 0.108
R40_401 s_0_89 s_0_88 0.108
R40_402 s_0_90 s_0_89 0.108
R40_403 s_0_91 s_0_90 0.108
R40_404 s_0_92 s_0_91 0.108
R40_405 s_0_93 s_0_92 0.864
R40_406 s_0_94 s_0_93 0.108
R40_407 s_0_95 s_0_94 0.108
R40_408 s_0_96 s_0_95 0.108
R40_409 s_0_97 s_0_96 0.108
R40_410 s_0_98 s_0_97 0.108
R40_411 s_0_99 s_0_98 0.108
R40_412 s_0_100 s_0_99 0.108
R40_413 s_0_101 s_0_100 0.108
R40_414 s_0_102 s_0_101 0.108
R40_415 s_0_103 s_0_102 0.108
R40_416 s_0_104 s_0_103 0.108
R40_417 s_0_105 s_0_104 0.108
R40_418 s_0_106 s_0_105 0.108
R40_419 s_0_107 s_0_106 0.108
R40_420 s_0_108 s_0_107 0.108
R40_421 s_0_109 s_0_108 0.108
R40_422 s_0_110 s_0_109 0.108
R40_423 s_0_111 s_0_110 0.108
R40_424 s_0_112 s_0_111 0.108
R40_425 s_0_113 s_0_112 0.001
R40_426 s_0_114 s_0_349 1.296
R40_427 s_0_115 s_0_114 0.108
R40_428 s_0_116 s_0_115 0.108
R40_429 s_0_117 s_0_116 0.108
R40_430 s_0_118 s_0_117 0.108
R40_431 s_0_119 s_0_118 0.108
R40_432 s_0_120 s_0_119 0.108
R40_433 s_0_121 s_0_120 0.108
R40_434 s_0_122 s_0_121 0.864
R40_435 s_0_123 s_0_122 0.108
R40_436 s_0_124 s_0_123 0.108
R40_437 s_0_125 s_0_124 0.108
R40_438 s_0_126 s_0_125 0.108
R40_439 s_0_127 s_0_126 0.108
R40_440 s_0_128 s_0_127 0.108
R40_441 s_0_129 s_0_128 0.108
R40_442 s_0_130 s_0_129 0.108
R40_443 s_0_131 s_0_130 0.108
R40_444 s_0_132 s_0_131 0.108
R40_445 s_0_133 s_0_132 0.108
R40_446 s_0_134 s_0_133 0.108
R40_447 s_0_135 s_0_134 0.108
R40_448 s_0_136 s_0_135 0.108
R40_449 s_0_137 s_0_136 0.108
R40_450 s_0_138 s_0_137 0.108
R40_451 s_0_139 s_0_138 0.108
R40_452 s_0_140 s_0_139 0.108
R40_453 s_0_141 s_0_140 0.108
R40_454 s_0_142 s_0_141 0.001
R40_455 s_0_143 s_0_349 1.296
R40_456 s_0_144 s_0_143 0.108
R40_457 s_0_145 s_0_144 0.108
R40_458 s_0_146 s_0_145 0.108
R40_459 s_0_147 s_0_146 0.108
R40_460 s_0_148 s_0_147 0.108
R40_461 s_0_149 s_0_148 0.108
R40_462 s_0_150 s_0_149 0.108
R40_463 s_0_151 s_0_150 0.864
R40_464 s_0_152 s_0_151 0.108
R40_465 s_0_153 s_0_152 0.108
R40_466 s_0_154 s_0_153 0.108
R40_467 s_0_155 s_0_154 0.108
R40_468 s_0_156 s_0_155 0.108
R40_469 s_0_157 s_0_156 0.108
R40_470 s_0_158 s_0_157 0.108
R40_471 s_0_159 s_0_158 0.108
R40_472 s_0_160 s_0_159 0.108
R40_473 s_0_161 s_0_160 0.108
R40_474 s_0_162 s_0_161 0.108
R40_475 s_0_163 s_0_162 0.108
R40_476 s_0_164 s_0_163 0.108
R40_477 s_0_165 s_0_164 0.108
R40_478 s_0_166 s_0_165 0.108
R40_479 s_0_167 s_0_166 0.108
R40_480 s_0_168 s_0_167 0.108
R40_481 s_0_169 s_0_168 0.108
R40_482 s_0_170 s_0_169 0.108
R40_483 s_0_171 s_0_170 0.001
R40_484 s_0_172 s_0_349 1.296
R40_485 s_0_173 s_0_172 0.108
R40_486 s_0_174 s_0_173 0.108
R40_487 s_0_175 s_0_174 0.108
R40_488 s_0_176 s_0_175 0.108
R40_489 s_0_177 s_0_176 0.108
R40_490 s_0_178 s_0_177 0.108
R40_491 s_0_179 s_0_178 0.108
R40_492 s_0_180 s_0_179 0.864
R40_493 s_0_181 s_0_180 0.108
R40_494 s_0_182 s_0_181 0.108
R40_495 s_0_183 s_0_182 0.108
R40_496 s_0_184 s_0_183 0.108
R40_497 s_0_185 s_0_184 0.108
R40_498 s_0_186 s_0_185 0.108
R40_499 s_0_187 s_0_186 0.108
R40_500 s_0_188 s_0_187 0.108
R40_501 s_0_189 s_0_188 0.108
R40_502 s_0_190 s_0_189 0.108
R40_503 s_0_191 s_0_190 0.108
R40_504 s_0_192 s_0_191 0.108
R40_505 s_0_193 s_0_192 0.108
R40_506 s_0_194 s_0_193 0.108
R40_507 s_0_195 s_0_194 0.108
R40_508 s_0_196 s_0_195 0.108
R40_509 s_0_197 s_0_196 0.108
R40_510 s_0_198 s_0_197 0.108
R40_511 s_0_199 s_0_198 0.108
R40_512 s_0_200 s_0_199 0.001
R40_513 s_0_201 s_0_349 1.296
R40_514 s_0_202 s_0_201 0.108
R40_515 s_0_203 s_0_202 0.108
R40_516 s_0_204 s_0_203 0.108
R40_517 s_0_205 s_0_204 0.108
R40_518 s_0_206 s_0_205 0.108
R40_519 s_0_207 s_0_206 0.108
R40_520 s_0_208 s_0_207 0.108
R40_521 s_0_209 s_0_208 0.864
R40_522 s_0_210 s_0_209 0.108
R40_523 s_0_211 s_0_210 0.108
R40_524 s_0_212 s_0_211 0.108
R40_525 s_0_213 s_0_212 0.108
R40_526 s_0_214 s_0_213 0.108
R40_527 s_0_215 s_0_214 0.108
R40_528 s_0_216 s_0_215 0.108
R40_529 s_0_217 s_0_216 0.108
R40_530 s_0_218 s_0_217 0.108
R40_531 s_0_219 s_0_218 0.108
R40_532 s_0_220 s_0_219 0.108
R40_533 s_0_221 s_0_220 0.108
R40_534 s_0_222 s_0_221 0.108
R40_535 s_0_223 s_0_222 0.108
R40_536 s_0_224 s_0_223 0.108
R40_537 s_0_225 s_0_224 0.108
R40_538 s_0_226 s_0_225 0.108
R40_539 s_0_227 s_0_226 0.108
R40_540 s_0_228 s_0_227 0.108
R40_541 s_0_229 s_0_228 0.001
R40_542 s_0_230 s_0_349 1.296
R40_543 s_0_231 s_0_230 0.108
R40_544 s_0_232 s_0_231 0.108
R40_545 s_0_233 s_0_232 0.108
R40_546 s_0_234 s_0_233 0.108
R40_547 s_0_235 s_0_234 0.108
R40_548 s_0_236 s_0_235 0.108
R40_549 s_0_237 s_0_236 0.108
R40_550 s_0_238 s_0_237 0.864
R40_551 s_0_239 s_0_238 0.108
R40_552 s_0_240 s_0_239 0.108
R40_553 s_0_241 s_0_240 0.108
R40_554 s_0_242 s_0_241 0.108
R40_555 s_0_243 s_0_242 0.108
R40_556 s_0_244 s_0_243 0.108
R40_557 s_0_245 s_0_244 0.108
R40_558 s_0_246 s_0_245 0.108
R40_559 s_0_247 s_0_246 0.108
R40_560 s_0_248 s_0_247 0.108
R40_561 s_0_249 s_0_248 0.108
R40_562 s_0_250 s_0_249 0.108
R40_563 s_0_251 s_0_250 0.108
R40_564 s_0_252 s_0_251 0.108
R40_565 s_0_253 s_0_252 0.108
R40_566 s_0_254 s_0_253 0.108
R40_567 s_0_255 s_0_254 0.108
R40_568 s_0_256 s_0_255 0.108
R40_569 s_0_257 s_0_256 0.108
R40_570 s_0_258 s_0_257 0.001
R40_571 s_0_259 s_0_349 1.296
R40_572 s_0_260 s_0_259 0.108
R40_573 s_0_261 s_0_260 0.108
R40_574 s_0_262 s_0_261 0.108
R40_575 s_0_263 s_0_262 0.108
R40_576 s_0_264 s_0_263 0.108
R40_577 s_0_265 s_0_264 0.108
R40_578 s_0_266 s_0_265 0.108
R40_579 s_0_267 s_0_266 0.864
R40_580 s_0_268 s_0_267 0.108
R40_581 s_0_269 s_0_268 0.108
R40_582 s_0_270 s_0_269 0.108
R40_583 s_0_271 s_0_270 0.108
R40_584 s_0_272 s_0_271 0.108
R40_585 s_0_273 s_0_272 0.108
R40_586 s_0_274 s_0_273 0.108
R40_587 s_0_275 s_0_274 0.108
R40_588 s_0_276 s_0_275 0.108
R40_589 s_0_277 s_0_276 0.108
R40_590 s_0_278 s_0_277 0.108
R40_591 s_0_279 s_0_278 0.108
R40_592 s_0_280 s_0_279 0.108
R40_593 s_0_281 s_0_280 0.108
R40_594 s_0_282 s_0_281 0.108
R40_595 s_0_283 s_0_282 0.108
R40_596 s_0_284 s_0_283 0.108
R40_597 s_0_285 s_0_284 0.108
R40_598 s_0_286 s_0_285 0.108
R40_599 s_0_287 s_0_286 0.001
R40_600 s_0_288 s_0_348 0.54
R40_601 s_0_289 s_0_288 0.108
R40_602 s_0_290 s_0_289 0.108
R40_603 s_0_291 s_0_290 0.108
R40_604 s_0_292 s_0_291 0.108
R40_605 s_0_293 s_0_292 0.108
R40_606 s_0_294 s_0_293 0.108
R40_607 s_0_295 s_0_294 0.108
R40_608 s_0_296 s_0_295 0.864
R40_609 s_0_297 s_0_296 0.108
R40_610 s_0_298 s_0_297 0.108
R40_611 s_0_299 s_0_298 0.108
R40_612 s_0_300 s_0_299 0.108
R40_613 s_0_301 s_0_300 0.108
R40_614 s_0_302 s_0_301 0.108
R40_615 s_0_303 s_0_302 0.108
R40_616 s_0_304 s_0_303 0.108
R40_617 s_0_305 s_0_304 0.108
R40_618 s_0_306 s_0_305 0.108
R40_619 s_0_307 s_0_306 0.108
R40_620 s_0_308 s_0_307 0.108
R40_621 s_0_309 s_0_308 0.108
R40_622 s_0_310 s_0_309 0.108
R40_623 s_0_311 s_0_310 0.108
R40_624 s_0_312 s_0_311 0.108
R40_625 s_0_313 s_0_312 0.108
R40_626 s_0_314 s_0_313 0.108
R40_627 s_0_315 s_0_314 0.108
R40_628 s_0_316 s_0_315 0.001
R40_629 s_0_317 s_0_346 0.54
R40_630 s_0_318 s_0_317 0.108
R40_631 s_0_319 s_0_318 0.108
R40_632 s_0_320 s_0_319 0.108
R40_633 s_0_321 s_0_320 0.108
R40_634 s_0_322 s_0_321 0.108
R40_635 s_0_323 s_0_322 0.108
R40_636 s_0_324 s_0_323 0.108
R40_637 s_0_325 s_0_324 0.864
R40_638 s_0_326 s_0_325 0.108
R40_639 s_0_327 s_0_326 0.108
R40_640 s_0_328 s_0_327 0.108
R40_641 s_0_329 s_0_328 0.108
R40_642 s_0_330 s_0_329 0.108
R40_643 s_0_331 s_0_330 0.108
R40_644 s_0_332 s_0_331 0.108
R40_645 s_0_333 s_0_332 0.108
R40_646 s_0_334 s_0_333 0.108
R40_647 s_0_335 s_0_334 0.108
R40_648 s_0_336 s_0_335 0.108
R40_649 s_0_337 s_0_336 0.108
R40_650 s_0_338 s_0_337 0.108
R40_651 s_0_339 s_0_338 0.108
R40_652 s_0_340 s_0_339 0.108
R40_653 s_0_341 s_0_340 0.108
R40_654 s_0_342 s_0_341 0.108
R40_655 s_0_343 s_0_342 0.108
R40_656 s_0_344 s_0_343 0.108
R40_657 s_0_345 s_0_344 0.001
R40_658 s_0_347 s_0_346 0.001
R40_659 s_0_348 s_0_347 0.001
R40_660 s_0_349 s_0_348 0.001
R40_661 s_0_350 s_0_349 0.001
R40_662 s_0_351 s_0_350 0.001
R40_663 s_0_352 s_0_351 0.001
R40_664 s_0_353 s_0_352 0.54
R40_665 s_0_354 s_0_353 0.108
R40_666 s_0_355 s_0_354 0.108
R40_667 s_0_356 s_0_355 0.108
R40_668 s_0_357 s_0_356 0.108
R40_669 s_0_358 s_0_357 0.108
R40_670 s_0_359 s_0_358 0.108
R40_671 s_0_360 s_0_359 0.108
R40_672 s_0_361 s_0_360 0.864
R40_673 s_0_362 s_0_361 0.108
R40_674 s_0_363 s_0_362 0.108
R40_675 s_0_364 s_0_363 0.108
R40_676 s_0_365 s_0_364 0.108
R40_677 s_0_366 s_0_365 0.108
R40_678 s_0_367 s_0_366 0.108
R40_679 s_0_368 s_0_367 0.108
R40_680 s_0_369 s_0_368 0.108
R40_681 s_0_370 s_0_369 0.108
R40_682 s_0_371 s_0_370 0.108
R40_683 s_0_372 s_0_371 0.108
R40_684 s_0_373 s_0_372 0.108
R40_685 s_0_374 s_0_373 0.108
R40_686 s_0_375 s_0_374 0.108
R40_687 s_0_376 s_0_375 0.108
R40_688 s_0_377 s_0_376 0.108
R40_689 s_0_378 s_0_377 0.108
R40_690 s_0_379 s_0_378 0.108
R40_691 s_0_380 s_0_379 0.108
R40_692 s_0_381 s_0_380 0.001

C710 s_0_349 vss 6.29069e-15
C711 s_0 vss 6.29069e-15
C712 s_0_27 vss 1.40901e-16
C713 s_0_350 vss 1.40901e-16
C714 s_0_28 vss 3.13114e-17
C715 s_0_27 vss 3.13114e-17
C716 s_0_29 vss 3.13114e-17
C717 s_0_28 vss 3.13114e-17
C718 s_0_30 vss 3.13114e-17
C719 s_0_29 vss 3.13114e-17
C720 s_0_31 vss 3.13114e-17
C721 s_0_30 vss 3.13114e-17
C722 s_0_32 vss 3.13114e-17
C723 s_0_31 vss 3.13114e-17
C724 s_0_33 vss 3.13114e-17
C725 s_0_32 vss 3.13114e-17
C726 s_0_34 vss 3.13114e-17
C727 s_0_33 vss 3.13114e-17
C728 s_0_35 vss 2.42663e-16
C729 s_0_34 vss 2.42663e-16
C730 s_0_36 vss 3.13114e-17
C731 s_0_35 vss 3.13114e-17
C732 s_0_37 vss 3.13114e-17
C733 s_0_36 vss 3.13114e-17
C734 s_0_38 vss 3.13114e-17
C735 s_0_37 vss 3.13114e-17
C736 s_0_39 vss 3.13114e-17
C737 s_0_38 vss 3.13114e-17
C738 s_0_40 vss 3.13114e-17
C739 s_0_39 vss 3.13114e-17
C740 s_0_41 vss 3.13114e-17
C741 s_0_40 vss 3.13114e-17
C742 s_0_42 vss 3.13114e-17
C743 s_0_41 vss 3.13114e-17
C744 s_0_43 vss 3.13114e-17
C745 s_0_42 vss 3.13114e-17
C746 s_0_44 vss 3.13114e-17
C747 s_0_43 vss 3.13114e-17
C748 s_0_45 vss 3.13114e-17
C749 s_0_44 vss 3.13114e-17
C750 s_0_46 vss 3.13114e-17
C751 s_0_45 vss 3.13114e-17
C752 s_0_47 vss 3.13114e-17
C753 s_0_46 vss 3.13114e-17
C754 s_0_48 vss 3.13114e-17
C755 s_0_47 vss 3.13114e-17
C756 s_0_49 vss 3.13114e-17
C757 s_0_48 vss 3.13114e-17
C758 s_0_50 vss 3.13114e-17
C759 s_0_49 vss 3.13114e-17
C760 s_0_51 vss 3.13114e-17
C761 s_0_50 vss 3.13114e-17
C762 s_0_52 vss 3.13114e-17
C763 s_0_51 vss 3.13114e-17
C764 s_0_53 vss 3.13114e-17
C765 s_0_52 vss 3.13114e-17
C766 s_0_54 vss 3.13114e-17
C767 s_0_53 vss 3.13114e-17
C768 s_0_55 vss 1.40901e-17
C769 s_0_54 vss 1.40901e-17
C770 s_0_56 vss 3.60081e-16
C771 s_0_349 vss 3.60081e-16
C772 s_0_57 vss 3.13114e-17
C773 s_0_56 vss 3.13114e-17
C774 s_0_58 vss 3.13114e-17
C775 s_0_57 vss 3.13114e-17
C776 s_0_59 vss 3.13114e-17
C777 s_0_58 vss 3.13114e-17
C778 s_0_60 vss 3.13114e-17
C779 s_0_59 vss 3.13114e-17
C780 s_0_61 vss 3.13114e-17
C781 s_0_60 vss 3.13114e-17
C782 s_0_62 vss 3.13114e-17
C783 s_0_61 vss 3.13114e-17
C784 s_0_63 vss 3.13114e-17
C785 s_0_62 vss 3.13114e-17
C786 s_0_64 vss 2.42663e-16
C787 s_0_63 vss 2.42663e-16
C788 s_0_65 vss 3.13114e-17
C789 s_0_64 vss 3.13114e-17
C790 s_0_66 vss 3.13114e-17
C791 s_0_65 vss 3.13114e-17
C792 s_0_67 vss 3.13114e-17
C793 s_0_66 vss 3.13114e-17
C794 s_0_68 vss 3.13114e-17
C795 s_0_67 vss 3.13114e-17
C796 s_0_69 vss 3.13114e-17
C797 s_0_68 vss 3.13114e-17
C798 s_0_70 vss 3.13114e-17
C799 s_0_69 vss 3.13114e-17
C800 s_0_71 vss 3.13114e-17
C801 s_0_70 vss 3.13114e-17
C802 s_0_72 vss 3.13114e-17
C803 s_0_71 vss 3.13114e-17
C804 s_0_73 vss 3.13114e-17
C805 s_0_72 vss 3.13114e-17
C806 s_0_74 vss 3.13114e-17
C807 s_0_73 vss 3.13114e-17
C808 s_0_75 vss 3.13114e-17
C809 s_0_74 vss 3.13114e-17
C810 s_0_76 vss 3.13114e-17
C811 s_0_75 vss 3.13114e-17
C812 s_0_77 vss 3.13114e-17
C813 s_0_76 vss 3.13114e-17
C814 s_0_78 vss 3.13114e-17
C815 s_0_77 vss 3.13114e-17
C816 s_0_79 vss 3.13114e-17
C817 s_0_78 vss 3.13114e-17
C818 s_0_80 vss 3.13114e-17
C819 s_0_79 vss 3.13114e-17
C820 s_0_81 vss 3.13114e-17
C821 s_0_80 vss 3.13114e-17
C822 s_0_82 vss 3.13114e-17
C823 s_0_81 vss 3.13114e-17
C824 s_0_83 vss 3.13114e-17
C825 s_0_82 vss 3.13114e-17
C826 s_0_84 vss 1.40901e-17
C827 s_0_83 vss 1.40901e-17
C828 s_0_85 vss 3.60081e-16
C829 s_0_349 vss 3.60081e-16
C830 s_0_86 vss 3.13114e-17
C831 s_0_85 vss 3.13114e-17
C832 s_0_87 vss 3.13114e-17
C833 s_0_86 vss 3.13114e-17
C834 s_0_88 vss 3.13114e-17
C835 s_0_87 vss 3.13114e-17
C836 s_0_89 vss 3.13114e-17
C837 s_0_88 vss 3.13114e-17
C838 s_0_90 vss 3.13114e-17
C839 s_0_89 vss 3.13114e-17
C840 s_0_91 vss 3.13114e-17
C841 s_0_90 vss 3.13114e-17
C842 s_0_92 vss 3.13114e-17
C843 s_0_91 vss 3.13114e-17
C844 s_0_93 vss 2.42663e-16
C845 s_0_92 vss 2.42663e-16
C846 s_0_94 vss 3.13114e-17
C847 s_0_93 vss 3.13114e-17
C848 s_0_95 vss 3.13114e-17
C849 s_0_94 vss 3.13114e-17
C850 s_0_96 vss 3.13114e-17
C851 s_0_95 vss 3.13114e-17
C852 s_0_97 vss 3.13114e-17
C853 s_0_96 vss 3.13114e-17
C854 s_0_98 vss 3.13114e-17
C855 s_0_97 vss 3.13114e-17
C856 s_0_99 vss 3.13114e-17
C857 s_0_98 vss 3.13114e-17
C858 s_0_100 vss 3.13114e-17
C859 s_0_99 vss 3.13114e-17
C860 s_0_101 vss 3.13114e-17
C861 s_0_100 vss 3.13114e-17
C862 s_0_102 vss 3.13114e-17
C863 s_0_101 vss 3.13114e-17
C864 s_0_103 vss 3.13114e-17
C865 s_0_102 vss 3.13114e-17
C866 s_0_104 vss 3.13114e-17
C867 s_0_103 vss 3.13114e-17
C868 s_0_105 vss 3.13114e-17
C869 s_0_104 vss 3.13114e-17
C870 s_0_106 vss 3.13114e-17
C871 s_0_105 vss 3.13114e-17
C872 s_0_107 vss 3.13114e-17
C873 s_0_106 vss 3.13114e-17
C874 s_0_108 vss 3.13114e-17
C875 s_0_107 vss 3.13114e-17
C876 s_0_109 vss 3.13114e-17
C877 s_0_108 vss 3.13114e-17
C878 s_0_110 vss 3.13114e-17
C879 s_0_109 vss 3.13114e-17
C880 s_0_111 vss 3.13114e-17
C881 s_0_110 vss 3.13114e-17
C882 s_0_112 vss 3.13114e-17
C883 s_0_111 vss 3.13114e-17
C884 s_0_113 vss 1.40901e-17
C885 s_0_112 vss 1.40901e-17
C886 s_0_114 vss 3.60081e-16
C887 s_0_349 vss 3.60081e-16
C888 s_0_115 vss 3.13114e-17
C889 s_0_114 vss 3.13114e-17
C890 s_0_116 vss 3.13114e-17
C891 s_0_115 vss 3.13114e-17
C892 s_0_117 vss 3.13114e-17
C893 s_0_116 vss 3.13114e-17
C894 s_0_118 vss 3.13114e-17
C895 s_0_117 vss 3.13114e-17
C896 s_0_119 vss 3.13114e-17
C897 s_0_118 vss 3.13114e-17
C898 s_0_120 vss 3.13114e-17
C899 s_0_119 vss 3.13114e-17
C900 s_0_121 vss 3.13114e-17
C901 s_0_120 vss 3.13114e-17
C902 s_0_122 vss 2.42663e-16
C903 s_0_121 vss 2.42663e-16
C904 s_0_123 vss 3.13114e-17
C905 s_0_122 vss 3.13114e-17
C906 s_0_124 vss 3.13114e-17
C907 s_0_123 vss 3.13114e-17
C908 s_0_125 vss 3.13114e-17
C909 s_0_124 vss 3.13114e-17
C910 s_0_126 vss 3.13114e-17
C911 s_0_125 vss 3.13114e-17
C912 s_0_127 vss 3.13114e-17
C913 s_0_126 vss 3.13114e-17
C914 s_0_128 vss 3.13114e-17
C915 s_0_127 vss 3.13114e-17
C916 s_0_129 vss 3.13114e-17
C917 s_0_128 vss 3.13114e-17
C918 s_0_130 vss 3.13114e-17
C919 s_0_129 vss 3.13114e-17
C920 s_0_131 vss 3.13114e-17
C921 s_0_130 vss 3.13114e-17
C922 s_0_132 vss 3.13114e-17
C923 s_0_131 vss 3.13114e-17
C924 s_0_133 vss 3.13114e-17
C925 s_0_132 vss 3.13114e-17
C926 s_0_134 vss 3.13114e-17
C927 s_0_133 vss 3.13114e-17
C928 s_0_135 vss 3.13114e-17
C929 s_0_134 vss 3.13114e-17
C930 s_0_136 vss 3.13114e-17
C931 s_0_135 vss 3.13114e-17
C932 s_0_137 vss 3.13114e-17
C933 s_0_136 vss 3.13114e-17
C934 s_0_138 vss 3.13114e-17
C935 s_0_137 vss 3.13114e-17
C936 s_0_139 vss 3.13114e-17
C937 s_0_138 vss 3.13114e-17
C938 s_0_140 vss 3.13114e-17
C939 s_0_139 vss 3.13114e-17
C940 s_0_141 vss 3.13114e-17
C941 s_0_140 vss 3.13114e-17
C942 s_0_142 vss 1.40901e-17
C943 s_0_141 vss 1.40901e-17
C944 s_0_143 vss 3.60081e-16
C945 s_0_349 vss 3.60081e-16
C946 s_0_144 vss 3.13114e-17
C947 s_0_143 vss 3.13114e-17
C948 s_0_145 vss 3.13114e-17
C949 s_0_144 vss 3.13114e-17
C950 s_0_146 vss 3.13114e-17
C951 s_0_145 vss 3.13114e-17
C952 s_0_147 vss 3.13114e-17
C953 s_0_146 vss 3.13114e-17
C954 s_0_148 vss 3.13114e-17
C955 s_0_147 vss 3.13114e-17
C956 s_0_149 vss 3.13114e-17
C957 s_0_148 vss 3.13114e-17
C958 s_0_150 vss 3.13114e-17
C959 s_0_149 vss 3.13114e-17
C960 s_0_151 vss 2.42663e-16
C961 s_0_150 vss 2.42663e-16
C962 s_0_152 vss 3.13114e-17
C963 s_0_151 vss 3.13114e-17
C964 s_0_153 vss 3.13114e-17
C965 s_0_152 vss 3.13114e-17
C966 s_0_154 vss 3.13114e-17
C967 s_0_153 vss 3.13114e-17
C968 s_0_155 vss 3.13114e-17
C969 s_0_154 vss 3.13114e-17
C970 s_0_156 vss 3.13114e-17
C971 s_0_155 vss 3.13114e-17
C972 s_0_157 vss 3.13114e-17
C973 s_0_156 vss 3.13114e-17
C974 s_0_158 vss 3.13114e-17
C975 s_0_157 vss 3.13114e-17
C976 s_0_159 vss 3.13114e-17
C977 s_0_158 vss 3.13114e-17
C978 s_0_160 vss 3.13114e-17
C979 s_0_159 vss 3.13114e-17
C980 s_0_161 vss 3.13114e-17
C981 s_0_160 vss 3.13114e-17
C982 s_0_162 vss 3.13114e-17
C983 s_0_161 vss 3.13114e-17
C984 s_0_163 vss 3.13114e-17
C985 s_0_162 vss 3.13114e-17
C986 s_0_164 vss 3.13114e-17
C987 s_0_163 vss 3.13114e-17
C988 s_0_165 vss 3.13114e-17
C989 s_0_164 vss 3.13114e-17
C990 s_0_166 vss 3.13114e-17
C991 s_0_165 vss 3.13114e-17
C992 s_0_167 vss 3.13114e-17
C993 s_0_166 vss 3.13114e-17
C994 s_0_168 vss 3.13114e-17
C995 s_0_167 vss 3.13114e-17
C996 s_0_169 vss 3.13114e-17
C997 s_0_168 vss 3.13114e-17
C998 s_0_170 vss 3.13114e-17
C999 s_0_169 vss 3.13114e-17
C1000 s_0_171 vss 1.40901e-17
C1001 s_0_170 vss 1.40901e-17
C1002 s_0_172 vss 3.60081e-16
C1003 s_0_349 vss 3.60081e-16
C1004 s_0_173 vss 3.13114e-17
C1005 s_0_172 vss 3.13114e-17
C1006 s_0_174 vss 3.13114e-17
C1007 s_0_173 vss 3.13114e-17
C1008 s_0_175 vss 3.13114e-17
C1009 s_0_174 vss 3.13114e-17
C1010 s_0_176 vss 3.13114e-17
C1011 s_0_175 vss 3.13114e-17
C1012 s_0_177 vss 3.13114e-17
C1013 s_0_176 vss 3.13114e-17
C1014 s_0_178 vss 3.13114e-17
C1015 s_0_177 vss 3.13114e-17
C1016 s_0_179 vss 3.13114e-17
C1017 s_0_178 vss 3.13114e-17
C1018 s_0_180 vss 2.42663e-16
C1019 s_0_179 vss 2.42663e-16
C1020 s_0_181 vss 3.13114e-17
C1021 s_0_180 vss 3.13114e-17
C1022 s_0_182 vss 3.13114e-17
C1023 s_0_181 vss 3.13114e-17
C1024 s_0_183 vss 3.13114e-17
C1025 s_0_182 vss 3.13114e-17
C1026 s_0_184 vss 3.13114e-17
C1027 s_0_183 vss 3.13114e-17
C1028 s_0_185 vss 3.13114e-17
C1029 s_0_184 vss 3.13114e-17
C1030 s_0_186 vss 3.13114e-17
C1031 s_0_185 vss 3.13114e-17
C1032 s_0_187 vss 3.13114e-17
C1033 s_0_186 vss 3.13114e-17
C1034 s_0_188 vss 3.13114e-17
C1035 s_0_187 vss 3.13114e-17
C1036 s_0_189 vss 3.13114e-17
C1037 s_0_188 vss 3.13114e-17
C1038 s_0_190 vss 3.13114e-17
C1039 s_0_189 vss 3.13114e-17
C1040 s_0_191 vss 3.13114e-17
C1041 s_0_190 vss 3.13114e-17
C1042 s_0_192 vss 3.13114e-17
C1043 s_0_191 vss 3.13114e-17
C1044 s_0_193 vss 3.13114e-17
C1045 s_0_192 vss 3.13114e-17
C1046 s_0_194 vss 3.13114e-17
C1047 s_0_193 vss 3.13114e-17
C1048 s_0_195 vss 3.13114e-17
C1049 s_0_194 vss 3.13114e-17
C1050 s_0_196 vss 3.13114e-17
C1051 s_0_195 vss 3.13114e-17
C1052 s_0_197 vss 3.13114e-17
C1053 s_0_196 vss 3.13114e-17
C1054 s_0_198 vss 3.13114e-17
C1055 s_0_197 vss 3.13114e-17
C1056 s_0_199 vss 3.13114e-17
C1057 s_0_198 vss 3.13114e-17
C1058 s_0_200 vss 1.40901e-17
C1059 s_0_199 vss 1.40901e-17
C1060 s_0_201 vss 3.60081e-16
C1061 s_0_349 vss 3.60081e-16
C1062 s_0_202 vss 3.13114e-17
C1063 s_0_201 vss 3.13114e-17
C1064 s_0_203 vss 3.13114e-17
C1065 s_0_202 vss 3.13114e-17
C1066 s_0_204 vss 3.13114e-17
C1067 s_0_203 vss 3.13114e-17
C1068 s_0_205 vss 3.13114e-17
C1069 s_0_204 vss 3.13114e-17
C1070 s_0_206 vss 3.13114e-17
C1071 s_0_205 vss 3.13114e-17
C1072 s_0_207 vss 3.13114e-17
C1073 s_0_206 vss 3.13114e-17
C1074 s_0_208 vss 3.13114e-17
C1075 s_0_207 vss 3.13114e-17
C1076 s_0_209 vss 2.42663e-16
C1077 s_0_208 vss 2.42663e-16
C1078 s_0_210 vss 3.13114e-17
C1079 s_0_209 vss 3.13114e-17
C1080 s_0_211 vss 3.13114e-17
C1081 s_0_210 vss 3.13114e-17
C1082 s_0_212 vss 3.13114e-17
C1083 s_0_211 vss 3.13114e-17
C1084 s_0_213 vss 3.13114e-17
C1085 s_0_212 vss 3.13114e-17
C1086 s_0_214 vss 3.13114e-17
C1087 s_0_213 vss 3.13114e-17
C1088 s_0_215 vss 3.13114e-17
C1089 s_0_214 vss 3.13114e-17
C1090 s_0_216 vss 3.13114e-17
C1091 s_0_215 vss 3.13114e-17
C1092 s_0_217 vss 3.13114e-17
C1093 s_0_216 vss 3.13114e-17
C1094 s_0_218 vss 3.13114e-17
C1095 s_0_217 vss 3.13114e-17
C1096 s_0_219 vss 3.13114e-17
C1097 s_0_218 vss 3.13114e-17
C1098 s_0_220 vss 3.13114e-17
C1099 s_0_219 vss 3.13114e-17
C1100 s_0_221 vss 3.13114e-17
C1101 s_0_220 vss 3.13114e-17
C1102 s_0_222 vss 3.13114e-17
C1103 s_0_221 vss 3.13114e-17
C1104 s_0_223 vss 3.13114e-17
C1105 s_0_222 vss 3.13114e-17
C1106 s_0_224 vss 3.13114e-17
C1107 s_0_223 vss 3.13114e-17
C1108 s_0_225 vss 3.13114e-17
C1109 s_0_224 vss 3.13114e-17
C1110 s_0_226 vss 3.13114e-17
C1111 s_0_225 vss 3.13114e-17
C1112 s_0_227 vss 3.13114e-17
C1113 s_0_226 vss 3.13114e-17
C1114 s_0_228 vss 3.13114e-17
C1115 s_0_227 vss 3.13114e-17
C1116 s_0_229 vss 1.40901e-17
C1117 s_0_228 vss 1.40901e-17
C1118 s_0_230 vss 3.60081e-16
C1119 s_0_349 vss 3.60081e-16
C1120 s_0_231 vss 3.13114e-17
C1121 s_0_230 vss 3.13114e-17
C1122 s_0_232 vss 3.13114e-17
C1123 s_0_231 vss 3.13114e-17
C1124 s_0_233 vss 3.13114e-17
C1125 s_0_232 vss 3.13114e-17
C1126 s_0_234 vss 3.13114e-17
C1127 s_0_233 vss 3.13114e-17
C1128 s_0_235 vss 3.13114e-17
C1129 s_0_234 vss 3.13114e-17
C1130 s_0_236 vss 3.13114e-17
C1131 s_0_235 vss 3.13114e-17
C1132 s_0_237 vss 3.13114e-17
C1133 s_0_236 vss 3.13114e-17
C1134 s_0_238 vss 2.42663e-16
C1135 s_0_237 vss 2.42663e-16
C1136 s_0_239 vss 3.13114e-17
C1137 s_0_238 vss 3.13114e-17
C1138 s_0_240 vss 3.13114e-17
C1139 s_0_239 vss 3.13114e-17
C1140 s_0_241 vss 3.13114e-17
C1141 s_0_240 vss 3.13114e-17
C1142 s_0_242 vss 3.13114e-17
C1143 s_0_241 vss 3.13114e-17
C1144 s_0_243 vss 3.13114e-17
C1145 s_0_242 vss 3.13114e-17
C1146 s_0_244 vss 3.13114e-17
C1147 s_0_243 vss 3.13114e-17
C1148 s_0_245 vss 3.13114e-17
C1149 s_0_244 vss 3.13114e-17
C1150 s_0_246 vss 3.13114e-17
C1151 s_0_245 vss 3.13114e-17
C1152 s_0_247 vss 3.13114e-17
C1153 s_0_246 vss 3.13114e-17
C1154 s_0_248 vss 3.13114e-17
C1155 s_0_247 vss 3.13114e-17
C1156 s_0_249 vss 3.13114e-17
C1157 s_0_248 vss 3.13114e-17
C1158 s_0_250 vss 3.13114e-17
C1159 s_0_249 vss 3.13114e-17
C1160 s_0_251 vss 3.13114e-17
C1161 s_0_250 vss 3.13114e-17
C1162 s_0_252 vss 3.13114e-17
C1163 s_0_251 vss 3.13114e-17
C1164 s_0_253 vss 3.13114e-17
C1165 s_0_252 vss 3.13114e-17
C1166 s_0_254 vss 3.13114e-17
C1167 s_0_253 vss 3.13114e-17
C1168 s_0_255 vss 3.13114e-17
C1169 s_0_254 vss 3.13114e-17
C1170 s_0_256 vss 3.13114e-17
C1171 s_0_255 vss 3.13114e-17
C1172 s_0_257 vss 3.13114e-17
C1173 s_0_256 vss 3.13114e-17
C1174 s_0_258 vss 1.40901e-17
C1175 s_0_257 vss 1.40901e-17
C1176 s_0_259 vss 3.60081e-16
C1177 s_0_349 vss 3.60081e-16
C1178 s_0_260 vss 3.13114e-17
C1179 s_0_259 vss 3.13114e-17
C1180 s_0_261 vss 3.13114e-17
C1181 s_0_260 vss 3.13114e-17
C1182 s_0_262 vss 3.13114e-17
C1183 s_0_261 vss 3.13114e-17
C1184 s_0_263 vss 3.13114e-17
C1185 s_0_262 vss 3.13114e-17
C1186 s_0_264 vss 3.13114e-17
C1187 s_0_263 vss 3.13114e-17
C1188 s_0_265 vss 3.13114e-17
C1189 s_0_264 vss 3.13114e-17
C1190 s_0_266 vss 3.13114e-17
C1191 s_0_265 vss 3.13114e-17
C1192 s_0_267 vss 2.42663e-16
C1193 s_0_266 vss 2.42663e-16
C1194 s_0_268 vss 3.13114e-17
C1195 s_0_267 vss 3.13114e-17
C1196 s_0_269 vss 3.13114e-17
C1197 s_0_268 vss 3.13114e-17
C1198 s_0_270 vss 3.13114e-17
C1199 s_0_269 vss 3.13114e-17
C1200 s_0_271 vss 3.13114e-17
C1201 s_0_270 vss 3.13114e-17
C1202 s_0_272 vss 3.13114e-17
C1203 s_0_271 vss 3.13114e-17
C1204 s_0_273 vss 3.13114e-17
C1205 s_0_272 vss 3.13114e-17
C1206 s_0_274 vss 3.13114e-17
C1207 s_0_273 vss 3.13114e-17
C1208 s_0_275 vss 3.13114e-17
C1209 s_0_274 vss 3.13114e-17
C1210 s_0_276 vss 3.13114e-17
C1211 s_0_275 vss 3.13114e-17
C1212 s_0_277 vss 3.13114e-17
C1213 s_0_276 vss 3.13114e-17
C1214 s_0_278 vss 3.13114e-17
C1215 s_0_277 vss 3.13114e-17
C1216 s_0_279 vss 3.13114e-17
C1217 s_0_278 vss 3.13114e-17
C1218 s_0_280 vss 3.13114e-17
C1219 s_0_279 vss 3.13114e-17
C1220 s_0_281 vss 3.13114e-17
C1221 s_0_280 vss 3.13114e-17
C1222 s_0_282 vss 3.13114e-17
C1223 s_0_281 vss 3.13114e-17
C1224 s_0_283 vss 3.13114e-17
C1225 s_0_282 vss 3.13114e-17
C1226 s_0_284 vss 3.13114e-17
C1227 s_0_283 vss 3.13114e-17
C1228 s_0_285 vss 3.13114e-17
C1229 s_0_284 vss 3.13114e-17
C1230 s_0_286 vss 3.13114e-17
C1231 s_0_285 vss 3.13114e-17
C1232 s_0_287 vss 1.40901e-17
C1233 s_0_286 vss 1.40901e-17
C1234 s_0_288 vss 1.40901e-16
C1235 s_0_348 vss 1.40901e-16
C1236 s_0_289 vss 3.13114e-17
C1237 s_0_288 vss 3.13114e-17
C1238 s_0_290 vss 3.13114e-17
C1239 s_0_289 vss 3.13114e-17
C1240 s_0_291 vss 3.13114e-17
C1241 s_0_290 vss 3.13114e-17
C1242 s_0_292 vss 3.13114e-17
C1243 s_0_291 vss 3.13114e-17
C1244 s_0_293 vss 3.13114e-17
C1245 s_0_292 vss 3.13114e-17
C1246 s_0_294 vss 3.13114e-17
C1247 s_0_293 vss 3.13114e-17
C1248 s_0_295 vss 3.13114e-17
C1249 s_0_294 vss 3.13114e-17
C1250 s_0_296 vss 2.42663e-16
C1251 s_0_295 vss 2.42663e-16
C1252 s_0_297 vss 3.13114e-17
C1253 s_0_296 vss 3.13114e-17
C1254 s_0_298 vss 3.13114e-17
C1255 s_0_297 vss 3.13114e-17
C1256 s_0_299 vss 3.13114e-17
C1257 s_0_298 vss 3.13114e-17
C1258 s_0_300 vss 3.13114e-17
C1259 s_0_299 vss 3.13114e-17
C1260 s_0_301 vss 3.13114e-17
C1261 s_0_300 vss 3.13114e-17
C1262 s_0_302 vss 3.13114e-17
C1263 s_0_301 vss 3.13114e-17
C1264 s_0_303 vss 3.13114e-17
C1265 s_0_302 vss 3.13114e-17
C1266 s_0_304 vss 3.13114e-17
C1267 s_0_303 vss 3.13114e-17
C1268 s_0_305 vss 3.13114e-17
C1269 s_0_304 vss 3.13114e-17
C1270 s_0_306 vss 3.13114e-17
C1271 s_0_305 vss 3.13114e-17
C1272 s_0_307 vss 3.13114e-17
C1273 s_0_306 vss 3.13114e-17
C1274 s_0_308 vss 3.13114e-17
C1275 s_0_307 vss 3.13114e-17
C1276 s_0_309 vss 3.13114e-17
C1277 s_0_308 vss 3.13114e-17
C1278 s_0_310 vss 3.13114e-17
C1279 s_0_309 vss 3.13114e-17
C1280 s_0_311 vss 3.13114e-17
C1281 s_0_310 vss 3.13114e-17
C1282 s_0_312 vss 3.13114e-17
C1283 s_0_311 vss 3.13114e-17
C1284 s_0_313 vss 3.13114e-17
C1285 s_0_312 vss 3.13114e-17
C1286 s_0_314 vss 3.13114e-17
C1287 s_0_313 vss 3.13114e-17
C1288 s_0_315 vss 3.13114e-17
C1289 s_0_314 vss 3.13114e-17
C1290 s_0_316 vss 1.40901e-17
C1291 s_0_315 vss 1.40901e-17
C1292 s_0_317 vss 1.40901e-16
C1293 s_0_346 vss 1.40901e-16
C1294 s_0_318 vss 3.13114e-17
C1295 s_0_317 vss 3.13114e-17
C1296 s_0_319 vss 3.13114e-17
C1297 s_0_318 vss 3.13114e-17
C1298 s_0_320 vss 3.13114e-17
C1299 s_0_319 vss 3.13114e-17
C1300 s_0_321 vss 3.13114e-17
C1301 s_0_320 vss 3.13114e-17
C1302 s_0_322 vss 3.13114e-17
C1303 s_0_321 vss 3.13114e-17
C1304 s_0_323 vss 3.13114e-17
C1305 s_0_322 vss 3.13114e-17
C1306 s_0_324 vss 3.13114e-17
C1307 s_0_323 vss 3.13114e-17
C1308 s_0_325 vss 2.42663e-16
C1309 s_0_324 vss 2.42663e-16
C1310 s_0_326 vss 3.13114e-17
C1311 s_0_325 vss 3.13114e-17
C1312 s_0_327 vss 3.13114e-17
C1313 s_0_326 vss 3.13114e-17
C1314 s_0_328 vss 3.13114e-17
C1315 s_0_327 vss 3.13114e-17
C1316 s_0_329 vss 3.13114e-17
C1317 s_0_328 vss 3.13114e-17
C1318 s_0_330 vss 3.13114e-17
C1319 s_0_329 vss 3.13114e-17
C1320 s_0_331 vss 3.13114e-17
C1321 s_0_330 vss 3.13114e-17
C1322 s_0_332 vss 3.13114e-17
C1323 s_0_331 vss 3.13114e-17
C1324 s_0_333 vss 3.13114e-17
C1325 s_0_332 vss 3.13114e-17
C1326 s_0_334 vss 3.13114e-17
C1327 s_0_333 vss 3.13114e-17
C1328 s_0_335 vss 3.13114e-17
C1329 s_0_334 vss 3.13114e-17
C1330 s_0_336 vss 3.13114e-17
C1331 s_0_335 vss 3.13114e-17
C1332 s_0_337 vss 3.13114e-17
C1333 s_0_336 vss 3.13114e-17
C1334 s_0_338 vss 3.13114e-17
C1335 s_0_337 vss 3.13114e-17
C1336 s_0_339 vss 3.13114e-17
C1337 s_0_338 vss 3.13114e-17
C1338 s_0_340 vss 3.13114e-17
C1339 s_0_339 vss 3.13114e-17
C1340 s_0_341 vss 3.13114e-17
C1341 s_0_340 vss 3.13114e-17
C1342 s_0_342 vss 3.13114e-17
C1343 s_0_341 vss 3.13114e-17
C1344 s_0_343 vss 3.13114e-17
C1345 s_0_342 vss 3.13114e-17
C1346 s_0_344 vss 3.13114e-17
C1347 s_0_343 vss 3.13114e-17
C1348 s_0_345 vss 1.40901e-17
C1349 s_0_344 vss 1.40901e-17
C1350 s_0_347 vss 2.95333e-17
C1351 s_0_346 vss 2.95333e-17
C1352 s_0_348 vss 3.71708e-16
C1353 s_0_347 vss 3.71708e-16
C1354 s_0_349 vss 2.15831e-15
C1355 s_0_348 vss 2.15831e-15
C1356 s_0_350 vss 2.15831e-15
C1357 s_0_349 vss 2.15831e-15
C1358 s_0_351 vss 3.71708e-16
C1359 s_0_350 vss 3.71708e-16
C1360 s_0_352 vss 2.95333e-17
C1361 s_0_351 vss 2.95333e-17
C1362 s_0_353 vss 1.40901e-16
C1363 s_0_352 vss 1.40901e-16
C1364 s_0_354 vss 3.13114e-17
C1365 s_0_353 vss 3.13114e-17
C1366 s_0_355 vss 3.13114e-17
C1367 s_0_354 vss 3.13114e-17
C1368 s_0_356 vss 3.13114e-17
C1369 s_0_355 vss 3.13114e-17
C1370 s_0_357 vss 3.13114e-17
C1371 s_0_356 vss 3.13114e-17
C1372 s_0_358 vss 3.13114e-17
C1373 s_0_357 vss 3.13114e-17
C1374 s_0_359 vss 3.13114e-17
C1375 s_0_358 vss 3.13114e-17
C1376 s_0_360 vss 3.13114e-17
C1377 s_0_359 vss 3.13114e-17
C1378 s_0_361 vss 2.42663e-16
C1379 s_0_360 vss 2.42663e-16
C1380 s_0_362 vss 3.13114e-17
C1381 s_0_361 vss 3.13114e-17
C1382 s_0_363 vss 3.13114e-17
C1383 s_0_362 vss 3.13114e-17
C1384 s_0_364 vss 3.13114e-17
C1385 s_0_363 vss 3.13114e-17
C1386 s_0_365 vss 3.13114e-17
C1387 s_0_364 vss 3.13114e-17
C1388 s_0_366 vss 3.13114e-17
C1389 s_0_365 vss 3.13114e-17
C1390 s_0_367 vss 3.13114e-17
C1391 s_0_366 vss 3.13114e-17
C1392 s_0_368 vss 3.13114e-17
C1393 s_0_367 vss 3.13114e-17
C1394 s_0_369 vss 3.13114e-17
C1395 s_0_368 vss 3.13114e-17
C1396 s_0_370 vss 3.13114e-17
C1397 s_0_369 vss 3.13114e-17
C1398 s_0_371 vss 3.13114e-17
C1399 s_0_370 vss 3.13114e-17
C1400 s_0_372 vss 3.13114e-17
C1401 s_0_371 vss 3.13114e-17
C1402 s_0_373 vss 3.13114e-17
C1403 s_0_372 vss 3.13114e-17
C1404 s_0_374 vss 3.13114e-17
C1405 s_0_373 vss 3.13114e-17
C1406 s_0_375 vss 3.13114e-17
C1407 s_0_374 vss 3.13114e-17
C1408 s_0_376 vss 3.13114e-17
C1409 s_0_375 vss 3.13114e-17
C1410 s_0_377 vss 3.13114e-17
C1411 s_0_376 vss 3.13114e-17
C1412 s_0_378 vss 3.13114e-17
C1413 s_0_377 vss 3.13114e-17
C1414 s_0_379 vss 3.13114e-17
C1415 s_0_378 vss 3.13114e-17
C1416 s_0_380 vss 3.13114e-17
C1417 s_0_379 vss 3.13114e-17
C1418 s_0_381 vss 1.40901e-17
C1419 s_0_380 vss 1.40901e-17

R41_1 n780 n780_27 0.001
R41_2 n780 n780_28 0.001
R41_3 n780 n780_26 0.001
R41_4 n780 n780_23 0.001
R41_5 n780 n780_22 0.001
R41_6 n780 n780_24 0.001
R41_7 n780 n780_25 0.001
R41_8 n780_20 n780_5 0.001
R41_9 n780_21 n780_4 0.001
R41_10 n780_18 n780_5 0.001
R41_11 n780_19 n780_5 0.001
R41_12 n780_16 n780_5 0.001
R41_13 n780_17 n780_5 0.001
R41_14 n780_13 n780_5 0.001
R41_15 n780_14 n780_5 0.001
R41_16 n780_15 n780_5 0.001
R41_17 n780_11 n780_5 0.001
R41_18 n780_10 n780_5 0.001
R41_19 n780_12 n780_5 0.001
R41_20 n780_9 n780_5 0.001
R41_21 n780_7 n780_5 0.001
R41_22 n780_8 n780_5 0.001
R41_23 n780_6 n780_5 0.001
R41_24 n780_2 n780_3 453.6
R41_25 n780_4 n780_3 14.4
R41_26 n780_7 n780_6 0.108
R41_27 n780_8 n780_7 0.108
R41_28 n780_9 n780_8 0.108
R41_29 n780_10 n780_9 0.108
R41_30 n780_11 n780_10 0.108
R41_31 n780_12 n780_11 0.108
R41_32 n780_13 n780_12 0.108
R41_33 n780_14 n780_13 0.108
R41_34 n780_15 n780_14 0.108
R41_35 n780_16 n780_15 0.108
R41_36 n780_17 n780_16 0.108
R41_37 n780_18 n780_17 0.108
R41_38 n780_19 n780_18 0.108
R41_39 n780_20 n780_19 0.108
R41_40 n780_21 n780_20 0.108
R41_41 n780_22 n780_21 0.756
R41_42 n780_23 n780_22 0.108
R41_43 n780_24 n780_23 0.108
R41_44 n780_25 n780_24 0.108
R41_45 n780_26 n780_25 0.108
R41_46 n780_27 n780_26 0.108
R41_47 n780_28 n780_27 0.108

C1420 n780_2 vss 4.98819e-16
C1421 n780_3 vss 4.98819e-16
C1422 n780_4 vss 8.41104e-17
C1423 n780_3 vss 8.41104e-17
C1424 n780_7 vss 2.92378e-17
C1425 n780_6 vss 2.92378e-17
C1426 n780_8 vss 2.92378e-17
C1427 n780_7 vss 2.92378e-17
C1428 n780_9 vss 2.92378e-17
C1429 n780_8 vss 2.92378e-17
C1430 n780_10 vss 2.92378e-17
C1431 n780_9 vss 2.92378e-17
C1432 n780_11 vss 2.92378e-17
C1433 n780_10 vss 2.92378e-17
C1434 n780_12 vss 2.92378e-17
C1435 n780_11 vss 2.92378e-17
C1436 n780_13 vss 2.92378e-17
C1437 n780_12 vss 2.92378e-17
C1438 n780_14 vss 2.92378e-17
C1439 n780_13 vss 2.92378e-17
C1440 n780_15 vss 2.92378e-17
C1441 n780_14 vss 2.92378e-17
C1442 n780_16 vss 2.92378e-17
C1443 n780_15 vss 2.92378e-17
C1444 n780_17 vss 2.92378e-17
C1445 n780_16 vss 2.92378e-17
C1446 n780_18 vss 2.92378e-17
C1447 n780_17 vss 2.92378e-17
C1448 n780_19 vss 2.92378e-17
C1449 n780_18 vss 2.92378e-17
C1450 n780_20 vss 2.92378e-17
C1451 n780_19 vss 2.92378e-17
C1452 n780_21 vss 3.65472e-17
C1453 n780_20 vss 3.65472e-17
C1454 n780_22 vss 1.46189e-16
C1455 n780_21 vss 1.46189e-16
C1456 n780_23 vss 2.92378e-17
C1457 n780_22 vss 2.92378e-17
C1458 n780_24 vss 2.92378e-17
C1459 n780_23 vss 2.92378e-17
C1460 n780_25 vss 2.92378e-17
C1461 n780_24 vss 2.92378e-17
C1462 n780_26 vss 2.92378e-17
C1463 n780_25 vss 2.92378e-17
C1464 n780_27 vss 2.92378e-17
C1465 n780_26 vss 2.92378e-17
C1466 n780_28 vss 2.92378e-17
C1467 n780_27 vss 2.92378e-17

R42_1 n817 n817_35 0.001
R42_2 n817 n817_36 0.001
R42_3 n817 n817_37 0.001
R42_4 n817 n817_33 0.001
R42_5 n817 n817_32 0.001
R42_6 n817 n817_31 0.001
R42_7 n817 n817_34 0.001
R42_8 n817_14 n817_11 0.001
R42_9 n817_29 n817_13 0.001
R42_10 n817_28 n817_13 0.001
R42_11 n817_25 n817_13 0.001
R42_12 n817_26 n817_13 0.001
R42_13 n817_27 n817_13 0.001
R42_14 n817_22 n817_13 0.001
R42_15 n817_23 n817_13 0.001
R42_16 n817_24 n817_13 0.001
R42_17 n817_21 n817_13 0.001
R42_18 n817_19 n817_13 0.001
R42_19 n817_20 n817_13 0.001
R42_20 n817_16 n817_13 0.001
R42_21 n817_15 n817_13 0.001
R42_22 n817_18 n817_13 0.001
R42_23 n817_17 n817_13 0.001
R42_24 n817_3 n817_2 43.2
R42_25 n817_12 n817_3 21.6
R42_26 n817_4 n817_12 21.6
R42_27 n817_5 n817_4 43.2
R42_28 n817_7 n817_6 43.2
R42_29 n817_10 n817_7 21.6
R42_30 n817_8 n817_10 21.6
R42_31 n817_9 n817_8 43.2
R42_32 n817_11 n817_10 28.8
R42_33 n817_12 n817_11 28.8
R42_34 n817_30 n817_14 0.648
R42_35 n817_16 n817_15 0.108
R42_36 n817_17 n817_16 0.108
R42_37 n817_18 n817_17 0.108
R42_38 n817_19 n817_18 0.108
R42_39 n817_20 n817_19 0.108
R42_40 n817_21 n817_20 0.108
R42_41 n817_22 n817_21 0.108
R42_42 n817_23 n817_22 0.108
R42_43 n817_24 n817_23 0.108
R42_44 n817_25 n817_24 0.108
R42_45 n817_26 n817_25 0.108
R42_46 n817_27 n817_26 0.108
R42_47 n817_28 n817_27 0.108
R42_48 n817_29 n817_28 0.108
R42_49 n817_30 n817_29 0.432
R42_50 n817_31 n817_30 0.54
R42_51 n817_32 n817_31 0.108
R42_52 n817_33 n817_32 0.108
R42_53 n817_34 n817_33 0.108
R42_54 n817_35 n817_34 0.108
R42_55 n817_36 n817_35 0.108
R42_56 n817_37 n817_36 0.108

C1468 n817_3 vss 4.69476e-17
C1469 n817_2 vss 4.69476e-17
C1470 n817_12 vss 2.34738e-17
C1471 n817_3 vss 2.34738e-17
C1472 n817_4 vss 2.34738e-17
C1473 n817_12 vss 2.34738e-17
C1474 n817_5 vss 4.69476e-17
C1475 n817_4 vss 4.69476e-17
C1476 n817_7 vss 4.69476e-17
C1477 n817_6 vss 4.69476e-17
C1478 n817_10 vss 2.34738e-17
C1479 n817_7 vss 2.34738e-17
C1480 n817_8 vss 2.34738e-17
C1481 n817_10 vss 2.34738e-17
C1482 n817_9 vss 4.69476e-17
C1483 n817_8 vss 4.69476e-17
C1484 n817_11 vss 7.33536e-17
C1485 n817_10 vss 7.33536e-17
C1486 n817_12 vss 8.25228e-17
C1487 n817_11 vss 8.25228e-17
C1488 n817_30 vss 1.3157e-16
C1489 n817_14 vss 1.3157e-16
C1490 n817_16 vss 2.92378e-17
C1491 n817_15 vss 2.92378e-17
C1492 n817_17 vss 2.92378e-17
C1493 n817_16 vss 2.92378e-17
C1494 n817_18 vss 2.92378e-17
C1495 n817_17 vss 2.92378e-17
C1496 n817_19 vss 2.92378e-17
C1497 n817_18 vss 2.92378e-17
C1498 n817_20 vss 2.92378e-17
C1499 n817_19 vss 2.92378e-17
C1500 n817_21 vss 2.92378e-17
C1501 n817_20 vss 2.92378e-17
C1502 n817_22 vss 2.92378e-17
C1503 n817_21 vss 2.92378e-17
C1504 n817_23 vss 2.92378e-17
C1505 n817_22 vss 2.92378e-17
C1506 n817_24 vss 2.92378e-17
C1507 n817_23 vss 2.92378e-17
C1508 n817_25 vss 2.92378e-17
C1509 n817_24 vss 2.92378e-17
C1510 n817_26 vss 2.92378e-17
C1511 n817_25 vss 2.92378e-17
C1512 n817_27 vss 2.92378e-17
C1513 n817_26 vss 2.92378e-17
C1514 n817_28 vss 2.92378e-17
C1515 n817_27 vss 2.92378e-17
C1516 n817_29 vss 2.92378e-17
C1517 n817_28 vss 2.92378e-17
C1518 n817_30 vss 8.77133e-17
C1519 n817_29 vss 8.77133e-17
C1520 n817_31 vss 9.50227e-17
C1521 n817_30 vss 9.50227e-17
C1522 n817_32 vss 2.92378e-17
C1523 n817_31 vss 2.92378e-17
C1524 n817_33 vss 2.92378e-17
C1525 n817_32 vss 2.92378e-17
C1526 n817_34 vss 2.92378e-17
C1527 n817_33 vss 2.92378e-17
C1528 n817_35 vss 2.92378e-17
C1529 n817_34 vss 2.92378e-17
C1530 n817_36 vss 2.92378e-17
C1531 n817_35 vss 2.92378e-17
C1532 n817_37 vss 2.92378e-17
C1533 n817_36 vss 2.92378e-17

R43_1 n939 n939_5 0.001
R43_2 n939 n939_8 0.001
R43_3 n939 n939_7 0.001
R43_4 n939_6 n939_23 0.001
R43_5 n939_22 n939_15 0.001
R43_6 n939_16 n939_10 0.001
R43_7 n939_17 n939_10 0.001
R43_8 n939_14 n939_10 0.001
R43_9 n939_19 n939_158 0.001
R43_10 n939_20 n939_159 0.001
R43_11 n939_21 n939_160 0.001
R43_12 n939 n939_2 0.001
R43_13 n939 n939_4 0.001
R43_14 n939 n939_3 0.001
R43_15 n939_12 n939_10 0.001
R43_16 n939_11 n939_10 0.001
R43_17 n939_13 n939_10 0.001
R43_18 n939_138 n939_24 0.001
R43_19 n939_137 n939_24 0.001
R43_20 n939_135 n939_24 0.001
R43_21 n939_136 n939_24 0.001
R43_22 n939_153 n939_25 0.001
R43_23 n939_150 n939_25 0.001
R43_24 n939_151 n939_25 0.001
R43_25 n939_152 n939_25 0.001
R43_26 n939_131 n939_24 0.001
R43_27 n939_132 n939_24 0.001
R43_28 n939_133 n939_24 0.001
R43_29 n939_134 n939_24 0.001
R43_30 n939_146 n939_25 0.001
R43_31 n939_149 n939_25 0.001
R43_32 n939_147 n939_25 0.001
R43_33 n939_148 n939_25 0.001
R43_34 n939_130 n939_24 0.001
R43_35 n939_127 n939_24 0.001
R43_36 n939_128 n939_24 0.001
R43_37 n939_129 n939_24 0.001
R43_38 n939_145 n939_25 0.001
R43_39 n939_142 n939_25 0.001
R43_40 n939_143 n939_25 0.001
R43_41 n939_144 n939_25 0.001
R43_42 n939_124 n939_24 0.001
R43_43 n939_125 n939_24 0.001
R43_44 n939_126 n939_24 0.001
R43_45 n939_140 n939_25 0.001
R43_46 n939_141 n939_25 0.001
R43_47 n939_139 n939_25 0.001
R43_48 n939_168 n939_28 0.001
R43_49 n939_167 n939_34 0.001
R43_50 n939_165 n939_40 0.001
R43_51 n939_164 n939_46 0.001
R43_52 n939_163 n939_52 0.001
R43_53 n939_162 n939_58 0.001
R43_54 n939_123 n939_63 0.001
R43_55 n939_62 n939_66 0.001
R43_56 n939_122 n939_72 0.001
R43_57 n939_71 n939_75 0.001
R43_58 n939_121 n939_81 0.001
R43_59 n939_80 n939_84 0.001
R43_60 n939_120 n939_90 0.001
R43_61 n939_89 n939_93 0.001
R43_62 n939_119 n939_99 0.001
R43_63 n939_98 n939_102 0.001
R43_64 n939_118 n939_108 0.001
R43_65 n939_107 n939_111 0.001
R43_66 n939_156 n939_116 0.001
R43_67 n939_154 n939_117 0.001
R43_68 n939_65 n939_64 21.6
R43_69 n939_68 n939_65 21.6
R43_70 n939_69 n939_68 43.2
R43_71 n939_70 n939_69 43.2
R43_72 n939_74 n939_73 21.6
R43_73 n939_77 n939_74 21.6
R43_74 n939_78 n939_77 43.2
R43_75 n939_79 n939_78 43.2
R43_76 n939_83 n939_82 21.6
R43_77 n939_86 n939_83 21.6
R43_78 n939_87 n939_86 43.2
R43_79 n939_88 n939_87 43.2
R43_80 n939_101 n939_100 21.6
R43_81 n939_104 n939_101 21.6
R43_82 n939_105 n939_104 43.2
R43_83 n939_106 n939_105 43.2
R43_84 n939_92 n939_91 21.6
R43_85 n939_95 n939_92 21.6
R43_86 n939_96 n939_95 43.2
R43_87 n939_97 n939_96 43.2
R43_88 n939_110 n939_109 21.6
R43_89 n939_113 n939_110 21.6
R43_90 n939_114 n939_113 43.2
R43_91 n939_115 n939_114 43.2
R43_92 n939_67 n939_65 28.8
R43_93 n939_76 n939_74 28.8
R43_94 n939_85 n939_83 28.8
R43_95 n939_103 n939_101 28.8
R43_96 n939_94 n939_92 28.8
R43_97 n939_112 n939_110 28.8
R43_98 n939_67 n939_66 7.2
R43_99 n939_76 n939_75 7.2
R43_100 n939_85 n939_84 7.2
R43_101 n939_103 n939_102 7.2
R43_102 n939_94 n939_93 7.2
R43_103 n939_112 n939_111 7.2
R43_104 n939_27 n939_26 21.6
R43_105 n939_29 n939_27 21.6
R43_106 n939_30 n939_29 43.2
R43_107 n939_31 n939_30 43.2
R43_108 n939_33 n939_32 21.6
R43_109 n939_35 n939_33 21.6
R43_110 n939_36 n939_35 43.2
R43_111 n939_37 n939_36 43.2
R43_112 n939_39 n939_38 21.6
R43_113 n939_41 n939_39 21.6
R43_114 n939_42 n939_41 43.2
R43_115 n939_43 n939_42 43.2
R43_116 n939_45 n939_44 21.6
R43_117 n939_47 n939_45 21.6
R43_118 n939_48 n939_47 43.2
R43_119 n939_49 n939_48 43.2
R43_120 n939_51 n939_50 21.6
R43_121 n939_53 n939_51 21.6
R43_122 n939_54 n939_53 43.2
R43_123 n939_55 n939_54 43.2
R43_124 n939_57 n939_56 21.6
R43_125 n939_59 n939_57 21.6
R43_126 n939_60 n939_59 43.2
R43_127 n939_61 n939_60 43.2
R43_128 n939_28 n939_27 28.8
R43_129 n939_34 n939_33 28.8
R43_130 n939_40 n939_39 28.8
R43_131 n939_46 n939_45 28.8
R43_132 n939_52 n939_51 28.8
R43_133 n939_58 n939_57 28.8
R43_134 n939_63 n939_62 0.216
R43_135 n939_72 n939_71 0.216
R43_136 n939_81 n939_80 0.216
R43_137 n939_99 n939_98 0.216
R43_138 n939_90 n939_89 0.216
R43_139 n939_108 n939_107 0.216
R43_140 n939_124 n939_166 0.648
R43_141 n939_125 n939_124 0.108
R43_142 n939_126 n939_125 0.108
R43_143 n939_127 n939_126 0.108
R43_144 n939_128 n939_127 0.108
R43_145 n939_129 n939_128 0.108
R43_146 n939_130 n939_129 0.108
R43_147 n939_131 n939_130 0.108
R43_148 n939_132 n939_131 0.108
R43_149 n939_133 n939_132 0.108
R43_150 n939_134 n939_133 0.108
R43_151 n939_135 n939_134 0.108
R43_152 n939_136 n939_135 0.108
R43_153 n939_137 n939_136 0.108
R43_154 n939_138 n939_137 0.108
R43_155 n939_139 n939_165 0.648
R43_156 n939_140 n939_139 0.108
R43_157 n939_141 n939_140 0.108
R43_158 n939_142 n939_141 0.108
R43_159 n939_143 n939_142 0.108
R43_160 n939_144 n939_143 0.108
R43_161 n939_145 n939_144 0.108
R43_162 n939_146 n939_145 0.108
R43_163 n939_147 n939_146 0.108
R43_164 n939_148 n939_147 0.108
R43_165 n939_149 n939_148 0.108
R43_166 n939_150 n939_149 0.108
R43_167 n939_151 n939_150 0.108
R43_168 n939_152 n939_151 0.108
R43_169 n939_153 n939_152 0.108
R43_170 n939_117 n939_116 0.054
R43_171 n939_118 n939_117 0.108
R43_172 n939_119 n939_118 0.432
R43_173 n939_120 n939_119 0.432
R43_174 n939_121 n939_120 0.432
R43_175 n939_122 n939_121 0.432
R43_176 n939_123 n939_122 0.432
R43_177 n939_162 n939_157 0.432
R43_178 n939_163 n939_162 0.648
R43_179 n939_164 n939_163 0.648
R43_180 n939_165 n939_164 0.648
R43_181 n939_166 n939_165 0.324
R43_182 n939_167 n939_166 0.216
R43_183 n939_168 n939_167 0.648
R43_184 n939_169 n939_168 0.001
R43_185 n939_154 n939_156 0.108
R43_186 n939_155 n939_154 0.001
R43_187 n939_12 n939_11 0.108
R43_188 n939_13 n939_12 0.108
R43_189 n939_14 n939_13 0.108
R43_190 n939_15 n939_14 0.108
R43_191 n939_16 n939_15 0.108
R43_192 n939_17 n939_16 0.108
R43_193 n939_18 n939_17 0.001
R43_194 n939_157 n939_156 3.024
R43_195 n939_158 n939_157 3.348
R43_196 n939_159 n939_158 0.108
R43_197 n939_160 n939_159 0.108
R43_198 n939_161 n939_160 0.001
R43_199 n939_20 n939_19 0.054
R43_200 n939_21 n939_20 0.054
R43_201 n939_22 n939_21 1.458
R43_202 n939_23 n939_22 0.216
R43_203 n939_3 n939_2 0.108
R43_204 n939_4 n939_3 0.108
R43_205 n939_5 n939_4 0.108
R43_206 n939_6 n939_5 0.108
R43_207 n939_7 n939_6 0.108
R43_208 n939_8 n939_7 0.108
R43_209 n939_9 n939_8 0.001

C1534 n939_65 vss 2.34738e-17
C1535 n939_64 vss 2.34738e-17
C1536 n939_68 vss 2.34738e-17
C1537 n939_65 vss 2.34738e-17
C1538 n939_69 vss 4.69476e-17
C1539 n939_68 vss 4.69476e-17
C1540 n939_70 vss 4.69476e-17
C1541 n939_69 vss 4.69476e-17
C1542 n939_74 vss 2.34738e-17
C1543 n939_73 vss 2.34738e-17
C1544 n939_77 vss 2.34738e-17
C1545 n939_74 vss 2.34738e-17
C1546 n939_78 vss 4.69476e-17
C1547 n939_77 vss 4.69476e-17
C1548 n939_79 vss 4.69476e-17
C1549 n939_78 vss 4.69476e-17
C1550 n939_83 vss 2.34738e-17
C1551 n939_82 vss 2.34738e-17
C1552 n939_86 vss 2.34738e-17
C1553 n939_83 vss 2.34738e-17
C1554 n939_87 vss 4.69476e-17
C1555 n939_86 vss 4.69476e-17
C1556 n939_88 vss 4.69476e-17
C1557 n939_87 vss 4.69476e-17
C1558 n939_101 vss 2.34738e-17
C1559 n939_100 vss 2.34738e-17
C1560 n939_104 vss 2.34738e-17
C1561 n939_101 vss 2.34738e-17
C1562 n939_105 vss 4.69476e-17
C1563 n939_104 vss 4.69476e-17
C1564 n939_106 vss 4.69476e-17
C1565 n939_105 vss 4.69476e-17
C1566 n939_92 vss 2.34738e-17
C1567 n939_91 vss 2.34738e-17
C1568 n939_95 vss 2.34738e-17
C1569 n939_92 vss 2.34738e-17
C1570 n939_96 vss 4.69476e-17
C1571 n939_95 vss 4.69476e-17
C1572 n939_97 vss 4.69476e-17
C1573 n939_96 vss 4.69476e-17
C1574 n939_110 vss 2.34738e-17
C1575 n939_109 vss 2.34738e-17
C1576 n939_113 vss 2.34738e-17
C1577 n939_110 vss 2.34738e-17
C1578 n939_114 vss 4.69476e-17
C1579 n939_113 vss 4.69476e-17
C1580 n939_115 vss 4.69476e-17
C1581 n939_114 vss 4.69476e-17
C1582 n939_67 vss 7.33536e-17
C1583 n939_65 vss 7.33536e-17
C1584 n939_76 vss 7.33536e-17
C1585 n939_74 vss 7.33536e-17
C1586 n939_85 vss 7.33536e-17
C1587 n939_83 vss 7.33536e-17
C1588 n939_103 vss 7.33536e-17
C1589 n939_101 vss 7.33536e-17
C1590 n939_94 vss 7.33536e-17
C1591 n939_92 vss 7.33536e-17
C1592 n939_112 vss 7.33536e-17
C1593 n939_110 vss 7.33536e-17
C1594 n939_67 vss 5.2569e-17
C1595 n939_66 vss 5.2569e-17
C1596 n939_76 vss 5.2569e-17
C1597 n939_75 vss 5.2569e-17
C1598 n939_85 vss 5.2569e-17
C1599 n939_84 vss 5.2569e-17
C1600 n939_103 vss 5.2569e-17
C1601 n939_102 vss 5.2569e-17
C1602 n939_94 vss 5.2569e-17
C1603 n939_93 vss 5.2569e-17
C1604 n939_112 vss 5.2569e-17
C1605 n939_111 vss 5.2569e-17
C1606 n939_27 vss 2.34738e-17
C1607 n939_26 vss 2.34738e-17
C1608 n939_29 vss 2.34738e-17
C1609 n939_27 vss 2.34738e-17
C1610 n939_30 vss 4.69476e-17
C1611 n939_29 vss 4.69476e-17
C1612 n939_31 vss 4.69476e-17
C1613 n939_30 vss 4.69476e-17
C1614 n939_33 vss 2.34738e-17
C1615 n939_32 vss 2.34738e-17
C1616 n939_35 vss 2.34738e-17
C1617 n939_33 vss 2.34738e-17
C1618 n939_36 vss 4.69476e-17
C1619 n939_35 vss 4.69476e-17
C1620 n939_37 vss 4.69476e-17
C1621 n939_36 vss 4.69476e-17
C1622 n939_39 vss 2.34738e-17
C1623 n939_38 vss 2.34738e-17
C1624 n939_41 vss 2.34738e-17
C1625 n939_39 vss 2.34738e-17
C1626 n939_42 vss 4.69476e-17
C1627 n939_41 vss 4.69476e-17
C1628 n939_43 vss 4.69476e-17
C1629 n939_42 vss 4.69476e-17
C1630 n939_45 vss 2.34738e-17
C1631 n939_44 vss 2.34738e-17
C1632 n939_47 vss 2.34738e-17
C1633 n939_45 vss 2.34738e-17
C1634 n939_48 vss 4.69476e-17
C1635 n939_47 vss 4.69476e-17
C1636 n939_49 vss 4.69476e-17
C1637 n939_48 vss 4.69476e-17
C1638 n939_51 vss 2.34738e-17
C1639 n939_50 vss 2.34738e-17
C1640 n939_53 vss 2.34738e-17
C1641 n939_51 vss 2.34738e-17
C1642 n939_54 vss 4.69476e-17
C1643 n939_53 vss 4.69476e-17
C1644 n939_55 vss 4.69476e-17
C1645 n939_54 vss 4.69476e-17
C1646 n939_57 vss 2.34738e-17
C1647 n939_56 vss 2.34738e-17
C1648 n939_59 vss 2.34738e-17
C1649 n939_57 vss 2.34738e-17
C1650 n939_60 vss 4.69476e-17
C1651 n939_59 vss 4.69476e-17
C1652 n939_61 vss 4.69476e-17
C1653 n939_60 vss 4.69476e-17
C1654 n939_28 vss 7.33536e-17
C1655 n939_27 vss 7.33536e-17
C1656 n939_34 vss 7.33536e-17
C1657 n939_33 vss 7.33536e-17
C1658 n939_40 vss 7.33536e-17
C1659 n939_39 vss 7.33536e-17
C1660 n939_46 vss 7.33536e-17
C1661 n939_45 vss 7.33536e-17
C1662 n939_52 vss 7.33536e-17
C1663 n939_51 vss 7.33536e-17
C1664 n939_58 vss 7.33536e-17
C1665 n939_57 vss 7.33536e-17
C1666 n939_63 vss 4.38566e-17
C1667 n939_62 vss 4.38566e-17
C1668 n939_72 vss 4.38566e-17
C1669 n939_71 vss 4.38566e-17
C1670 n939_81 vss 4.38566e-17
C1671 n939_80 vss 4.38566e-17
C1672 n939_99 vss 4.38566e-17
C1673 n939_98 vss 4.38566e-17
C1674 n939_90 vss 4.38566e-17
C1675 n939_89 vss 4.38566e-17
C1676 n939_108 vss 4.38566e-17
C1677 n939_107 vss 4.38566e-17
C1678 n939_124 vss 1.20606e-16
C1679 n939_166 vss 1.20606e-16
C1680 n939_125 vss 2.92378e-17
C1681 n939_124 vss 2.92378e-17
C1682 n939_126 vss 2.92378e-17
C1683 n939_125 vss 2.92378e-17
C1684 n939_127 vss 2.92378e-17
C1685 n939_126 vss 2.92378e-17
C1686 n939_128 vss 2.92378e-17
C1687 n939_127 vss 2.92378e-17
C1688 n939_129 vss 2.92378e-17
C1689 n939_128 vss 2.92378e-17
C1690 n939_130 vss 2.92378e-17
C1691 n939_129 vss 2.92378e-17
C1692 n939_131 vss 2.92378e-17
C1693 n939_130 vss 2.92378e-17
C1694 n939_132 vss 2.92378e-17
C1695 n939_131 vss 2.92378e-17
C1696 n939_133 vss 2.92378e-17
C1697 n939_132 vss 2.92378e-17
C1698 n939_134 vss 2.92378e-17
C1699 n939_133 vss 2.92378e-17
C1700 n939_135 vss 2.92378e-17
C1701 n939_134 vss 2.92378e-17
C1702 n939_136 vss 2.92378e-17
C1703 n939_135 vss 2.92378e-17
C1704 n939_137 vss 2.92378e-17
C1705 n939_136 vss 2.92378e-17
C1706 n939_138 vss 2.92378e-17
C1707 n939_137 vss 2.92378e-17
C1708 n939_139 vss 1.20606e-16
C1709 n939_165 vss 1.20606e-16
C1710 n939_140 vss 2.92378e-17
C1711 n939_139 vss 2.92378e-17
C1712 n939_141 vss 2.92378e-17
C1713 n939_140 vss 2.92378e-17
C1714 n939_142 vss 2.92378e-17
C1715 n939_141 vss 2.92378e-17
C1716 n939_143 vss 2.92378e-17
C1717 n939_142 vss 2.92378e-17
C1718 n939_144 vss 2.92378e-17
C1719 n939_143 vss 2.92378e-17
C1720 n939_145 vss 2.92378e-17
C1721 n939_144 vss 2.92378e-17
C1722 n939_146 vss 2.92378e-17
C1723 n939_145 vss 2.92378e-17
C1724 n939_147 vss 2.92378e-17
C1725 n939_146 vss 2.92378e-17
C1726 n939_148 vss 2.92378e-17
C1727 n939_147 vss 2.92378e-17
C1728 n939_149 vss 2.92378e-17
C1729 n939_148 vss 2.92378e-17
C1730 n939_150 vss 2.92378e-17
C1731 n939_149 vss 2.92378e-17
C1732 n939_151 vss 2.92378e-17
C1733 n939_150 vss 2.92378e-17
C1734 n939_152 vss 2.92378e-17
C1735 n939_151 vss 2.92378e-17
C1736 n939_153 vss 2.92378e-17
C1737 n939_152 vss 2.92378e-17
C1738 n939_117 vss 3.2562e-17
C1739 n939_116 vss 3.2562e-17
C1740 n939_118 vss 4.55868e-17
C1741 n939_117 vss 4.55868e-17
C1742 n939_119 vss 1.56298e-16
C1743 n939_118 vss 1.56298e-16
C1744 n939_120 vss 1.56298e-16
C1745 n939_119 vss 1.56298e-16
C1746 n939_121 vss 1.56298e-16
C1747 n939_120 vss 1.56298e-16
C1748 n939_122 vss 1.56298e-16
C1749 n939_121 vss 1.56298e-16
C1750 n939_123 vss 1.56298e-16
C1751 n939_122 vss 1.56298e-16
C1752 n939_162 vss 1.33073e-16
C1753 n939_157 vss 1.33073e-16
C1754 n939_163 vss 1.87868e-16
C1755 n939_162 vss 1.87868e-16
C1756 n939_164 vss 1.87868e-16
C1757 n939_163 vss 1.87868e-16
C1758 n939_165 vss 1.95696e-16
C1759 n939_164 vss 1.95696e-16
C1760 n939_166 vss 1.01762e-16
C1761 n939_165 vss 1.01762e-16
C1762 n939_167 vss 7.82784e-17
C1763 n939_166 vss 7.82784e-17
C1764 n939_168 vss 1.87868e-16
C1765 n939_167 vss 1.87868e-16
C1766 n939_169 vss 1.40901e-17
C1767 n939_168 vss 1.40901e-17
C1768 n939_154 vss 3.91392e-17
C1769 n939_156 vss 3.91392e-17
C1770 n939_155 vss 1.40901e-17
C1771 n939_154 vss 1.40901e-17
C1772 n939_12 vss 2.92378e-17
C1773 n939_11 vss 2.92378e-17
C1774 n939_13 vss 2.92378e-17
C1775 n939_12 vss 2.92378e-17
C1776 n939_14 vss 2.92378e-17
C1777 n939_13 vss 2.92378e-17
C1778 n939_15 vss 3.65472e-17
C1779 n939_14 vss 3.65472e-17
C1780 n939_16 vss 2.92378e-17
C1781 n939_15 vss 2.92378e-17
C1782 n939_17 vss 3.65472e-17
C1783 n939_16 vss 3.65472e-17
C1784 n939_18 vss 1.3157e-17
C1785 n939_17 vss 1.3157e-17
C1786 n939_157 vss 7.94526e-16
C1787 n939_156 vss 7.94526e-16
C1788 n939_158 vss 8.96288e-16
C1789 n939_157 vss 8.96288e-16
C1790 n939_159 vss 3.13114e-17
C1791 n939_158 vss 3.13114e-17
C1792 n939_160 vss 3.13114e-17
C1793 n939_159 vss 3.13114e-17
C1794 n939_161 vss 1.40901e-17
C1795 n939_160 vss 1.40901e-17
C1796 n939_20 vss 2.60496e-17
C1797 n939_19 vss 2.60496e-17
C1798 n939_21 vss 2.60496e-17
C1799 n939_20 vss 2.60496e-17
C1800 n939_22 vss 5.40529e-16
C1801 n939_21 vss 5.40529e-16
C1802 n939_23 vss 7.81488e-17
C1803 n939_22 vss 7.81488e-17
C1804 n939_3 vss 2.92378e-17
C1805 n939_2 vss 2.92378e-17
C1806 n939_4 vss 2.92378e-17
C1807 n939_3 vss 2.92378e-17
C1808 n939_5 vss 2.92378e-17
C1809 n939_4 vss 2.92378e-17
C1810 n939_6 vss 3.65472e-17
C1811 n939_5 vss 3.65472e-17
C1812 n939_7 vss 2.92378e-17
C1813 n939_6 vss 2.92378e-17
C1814 n939_8 vss 3.65472e-17
C1815 n939_7 vss 3.65472e-17
C1816 n939_9 vss 1.3157e-17
C1817 n939_8 vss 1.3157e-17

R44_1 n1110_23 n1110_6 0.001
R44_2 n1110_5 n1110 0.001
R44_3 n1110_8 n1110 0.001
R44_4 n1110_7 n1110 0.001
R44_5 n1110_10 n1110_14 0.001
R44_6 n1110_10 n1110_16 0.001
R44_7 n1110_10 n1110_17 0.001
R44_8 n1110_15 n1110_22 0.001
R44_9 n1110_19 n1110_158 0.001
R44_10 n1110_20 n1110_159 0.001
R44_11 n1110_21 n1110_160 0.001
R44_12 n1110_3 n1110 0.001
R44_13 n1110_2 n1110 0.001
R44_14 n1110_4 n1110 0.001
R44_15 n1110_10 n1110_12 0.001
R44_16 n1110_10 n1110_11 0.001
R44_17 n1110_10 n1110_13 0.001
R44_18 n1110_152 n1110_24 0.001
R44_19 n1110_150 n1110_24 0.001
R44_20 n1110_151 n1110_24 0.001
R44_21 n1110_153 n1110_24 0.001
R44_22 n1110_138 n1110_25 0.001
R44_23 n1110_135 n1110_25 0.001
R44_24 n1110_136 n1110_25 0.001
R44_25 n1110_137 n1110_25 0.001
R44_26 n1110_146 n1110_24 0.001
R44_27 n1110_148 n1110_24 0.001
R44_28 n1110_149 n1110_24 0.001
R44_29 n1110_147 n1110_24 0.001
R44_30 n1110_131 n1110_25 0.001
R44_31 n1110_132 n1110_25 0.001
R44_32 n1110_133 n1110_25 0.001
R44_33 n1110_134 n1110_25 0.001
R44_34 n1110_145 n1110_24 0.001
R44_35 n1110_142 n1110_24 0.001
R44_36 n1110_143 n1110_24 0.001
R44_37 n1110_144 n1110_24 0.001
R44_38 n1110_130 n1110_25 0.001
R44_39 n1110_127 n1110_25 0.001
R44_40 n1110_128 n1110_25 0.001
R44_41 n1110_129 n1110_25 0.001
R44_42 n1110_140 n1110_24 0.001
R44_43 n1110_141 n1110_24 0.001
R44_44 n1110_139 n1110_24 0.001
R44_45 n1110_126 n1110_25 0.001
R44_46 n1110_124 n1110_25 0.001
R44_47 n1110_125 n1110_25 0.001
R44_48 n1110_168 n1110_28 0.001
R44_49 n1110_167 n1110_34 0.001
R44_50 n1110_165 n1110_40 0.001
R44_51 n1110_164 n1110_46 0.001
R44_52 n1110_163 n1110_52 0.001
R44_53 n1110_162 n1110_58 0.001
R44_54 n1110_123 n1110_63 0.001
R44_55 n1110_62 n1110_66 0.001
R44_56 n1110_122 n1110_72 0.001
R44_57 n1110_71 n1110_75 0.001
R44_58 n1110_121 n1110_81 0.001
R44_59 n1110_80 n1110_84 0.001
R44_60 n1110_120 n1110_90 0.001
R44_61 n1110_89 n1110_93 0.001
R44_62 n1110_119 n1110_99 0.001
R44_63 n1110_98 n1110_102 0.001
R44_64 n1110_118 n1110_108 0.001
R44_65 n1110_107 n1110_111 0.001
R44_66 n1110_156 n1110_116 0.001
R44_67 n1110_154 n1110_117 0.001
R44_68 n1110_65 n1110_64 21.6
R44_69 n1110_68 n1110_65 21.6
R44_70 n1110_69 n1110_68 43.2
R44_71 n1110_70 n1110_69 43.2
R44_72 n1110_83 n1110_82 21.6
R44_73 n1110_86 n1110_83 21.6
R44_74 n1110_87 n1110_86 43.2
R44_75 n1110_88 n1110_87 43.2
R44_76 n1110_74 n1110_73 21.6
R44_77 n1110_77 n1110_74 21.6
R44_78 n1110_78 n1110_77 43.2
R44_79 n1110_79 n1110_78 43.2
R44_80 n1110_92 n1110_91 21.6
R44_81 n1110_95 n1110_92 21.6
R44_82 n1110_96 n1110_95 43.2
R44_83 n1110_97 n1110_96 43.2
R44_84 n1110_101 n1110_100 21.6
R44_85 n1110_104 n1110_101 21.6
R44_86 n1110_105 n1110_104 43.2
R44_87 n1110_106 n1110_105 43.2
R44_88 n1110_110 n1110_109 21.6
R44_89 n1110_113 n1110_110 21.6
R44_90 n1110_114 n1110_113 43.2
R44_91 n1110_115 n1110_114 43.2
R44_92 n1110_67 n1110_65 28.8
R44_93 n1110_85 n1110_83 28.8
R44_94 n1110_76 n1110_74 28.8
R44_95 n1110_94 n1110_92 28.8
R44_96 n1110_103 n1110_101 28.8
R44_97 n1110_112 n1110_110 28.8
R44_98 n1110_67 n1110_66 7.2
R44_99 n1110_85 n1110_84 7.2
R44_100 n1110_76 n1110_75 7.2
R44_101 n1110_94 n1110_93 7.2
R44_102 n1110_103 n1110_102 7.2
R44_103 n1110_112 n1110_111 7.2
R44_104 n1110_27 n1110_26 21.6
R44_105 n1110_29 n1110_27 21.6
R44_106 n1110_30 n1110_29 43.2
R44_107 n1110_31 n1110_30 43.2
R44_108 n1110_33 n1110_32 21.6
R44_109 n1110_35 n1110_33 21.6
R44_110 n1110_36 n1110_35 43.2
R44_111 n1110_37 n1110_36 43.2
R44_112 n1110_39 n1110_38 21.6
R44_113 n1110_41 n1110_39 21.6
R44_114 n1110_42 n1110_41 43.2
R44_115 n1110_43 n1110_42 43.2
R44_116 n1110_45 n1110_44 21.6
R44_117 n1110_47 n1110_45 21.6
R44_118 n1110_48 n1110_47 43.2
R44_119 n1110_49 n1110_48 43.2
R44_120 n1110_51 n1110_50 21.6
R44_121 n1110_53 n1110_51 21.6
R44_122 n1110_54 n1110_53 43.2
R44_123 n1110_55 n1110_54 43.2
R44_124 n1110_57 n1110_56 21.6
R44_125 n1110_59 n1110_57 21.6
R44_126 n1110_60 n1110_59 43.2
R44_127 n1110_61 n1110_60 43.2
R44_128 n1110_28 n1110_27 28.8
R44_129 n1110_34 n1110_33 28.8
R44_130 n1110_40 n1110_39 28.8
R44_131 n1110_46 n1110_45 28.8
R44_132 n1110_52 n1110_51 28.8
R44_133 n1110_58 n1110_57 28.8
R44_134 n1110_63 n1110_62 0.216
R44_135 n1110_81 n1110_80 0.216
R44_136 n1110_72 n1110_71 0.216
R44_137 n1110_90 n1110_89 0.216
R44_138 n1110_99 n1110_98 0.216
R44_139 n1110_108 n1110_107 0.216
R44_140 n1110_124 n1110_165 0.648
R44_141 n1110_125 n1110_124 0.108
R44_142 n1110_126 n1110_125 0.108
R44_143 n1110_127 n1110_126 0.108
R44_144 n1110_128 n1110_127 0.108
R44_145 n1110_129 n1110_128 0.108
R44_146 n1110_130 n1110_129 0.108
R44_147 n1110_131 n1110_130 0.108
R44_148 n1110_132 n1110_131 0.108
R44_149 n1110_133 n1110_132 0.108
R44_150 n1110_134 n1110_133 0.108
R44_151 n1110_135 n1110_134 0.108
R44_152 n1110_136 n1110_135 0.108
R44_153 n1110_137 n1110_136 0.108
R44_154 n1110_138 n1110_137 0.108
R44_155 n1110_139 n1110_166 0.648
R44_156 n1110_140 n1110_139 0.108
R44_157 n1110_141 n1110_140 0.108
R44_158 n1110_142 n1110_141 0.108
R44_159 n1110_143 n1110_142 0.108
R44_160 n1110_144 n1110_143 0.108
R44_161 n1110_145 n1110_144 0.108
R44_162 n1110_146 n1110_145 0.108
R44_163 n1110_147 n1110_146 0.108
R44_164 n1110_148 n1110_147 0.108
R44_165 n1110_149 n1110_148 0.108
R44_166 n1110_150 n1110_149 0.108
R44_167 n1110_151 n1110_150 0.108
R44_168 n1110_152 n1110_151 0.108
R44_169 n1110_153 n1110_152 0.108
R44_170 n1110_117 n1110_116 0.054
R44_171 n1110_118 n1110_117 0.108
R44_172 n1110_119 n1110_118 0.432
R44_173 n1110_120 n1110_119 0.432
R44_174 n1110_121 n1110_120 0.432
R44_175 n1110_122 n1110_121 0.432
R44_176 n1110_123 n1110_122 0.432
R44_177 n1110_162 n1110_157 0.432
R44_178 n1110_163 n1110_162 0.648
R44_179 n1110_164 n1110_163 0.648
R44_180 n1110_165 n1110_164 0.648
R44_181 n1110_166 n1110_165 0.324
R44_182 n1110_167 n1110_166 0.216
R44_183 n1110_168 n1110_167 0.648
R44_184 n1110_169 n1110_168 0.001
R44_185 n1110_154 n1110_156 0.108
R44_186 n1110_155 n1110_154 0.001
R44_187 n1110_3 n1110_2 0.108
R44_188 n1110_4 n1110_3 0.108
R44_189 n1110_5 n1110_4 0.108
R44_190 n1110_6 n1110_5 0.108
R44_191 n1110_7 n1110_6 0.108
R44_192 n1110_8 n1110_7 0.108
R44_193 n1110_9 n1110_8 0.001
R44_194 n1110_157 n1110_156 3.024
R44_195 n1110_158 n1110_157 3.348
R44_196 n1110_159 n1110_158 0.108
R44_197 n1110_160 n1110_159 0.108
R44_198 n1110_161 n1110_160 0.001
R44_199 n1110_20 n1110_19 0.054
R44_200 n1110_21 n1110_20 0.054
R44_201 n1110_22 n1110_21 1.458
R44_202 n1110_23 n1110_22 0.216
R44_203 n1110_12 n1110_11 0.108
R44_204 n1110_13 n1110_12 0.108
R44_205 n1110_14 n1110_13 0.108
R44_206 n1110_15 n1110_14 0.108
R44_207 n1110_16 n1110_15 0.108
R44_208 n1110_17 n1110_16 0.108
R44_209 n1110_18 n1110_17 0.001

C1818 n1110_65 vss 2.34738e-17
C1819 n1110_64 vss 2.34738e-17
C1820 n1110_68 vss 2.34738e-17
C1821 n1110_65 vss 2.34738e-17
C1822 n1110_69 vss 4.69476e-17
C1823 n1110_68 vss 4.69476e-17
C1824 n1110_70 vss 4.69476e-17
C1825 n1110_69 vss 4.69476e-17
C1826 n1110_83 vss 2.34738e-17
C1827 n1110_82 vss 2.34738e-17
C1828 n1110_86 vss 2.34738e-17
C1829 n1110_83 vss 2.34738e-17
C1830 n1110_87 vss 4.69476e-17
C1831 n1110_86 vss 4.69476e-17
C1832 n1110_88 vss 4.69476e-17
C1833 n1110_87 vss 4.69476e-17
C1834 n1110_74 vss 2.34738e-17
C1835 n1110_73 vss 2.34738e-17
C1836 n1110_77 vss 2.34738e-17
C1837 n1110_74 vss 2.34738e-17
C1838 n1110_78 vss 4.69476e-17
C1839 n1110_77 vss 4.69476e-17
C1840 n1110_79 vss 4.69476e-17
C1841 n1110_78 vss 4.69476e-17
C1842 n1110_92 vss 2.34738e-17
C1843 n1110_91 vss 2.34738e-17
C1844 n1110_95 vss 2.34738e-17
C1845 n1110_92 vss 2.34738e-17
C1846 n1110_96 vss 4.69476e-17
C1847 n1110_95 vss 4.69476e-17
C1848 n1110_97 vss 4.69476e-17
C1849 n1110_96 vss 4.69476e-17
C1850 n1110_101 vss 2.34738e-17
C1851 n1110_100 vss 2.34738e-17
C1852 n1110_104 vss 2.34738e-17
C1853 n1110_101 vss 2.34738e-17
C1854 n1110_105 vss 4.69476e-17
C1855 n1110_104 vss 4.69476e-17
C1856 n1110_106 vss 4.69476e-17
C1857 n1110_105 vss 4.69476e-17
C1858 n1110_110 vss 2.34738e-17
C1859 n1110_109 vss 2.34738e-17
C1860 n1110_113 vss 2.34738e-17
C1861 n1110_110 vss 2.34738e-17
C1862 n1110_114 vss 4.69476e-17
C1863 n1110_113 vss 4.69476e-17
C1864 n1110_115 vss 4.69476e-17
C1865 n1110_114 vss 4.69476e-17
C1866 n1110_67 vss 7.33536e-17
C1867 n1110_65 vss 7.33536e-17
C1868 n1110_85 vss 7.33536e-17
C1869 n1110_83 vss 7.33536e-17
C1870 n1110_76 vss 7.33536e-17
C1871 n1110_74 vss 7.33536e-17
C1872 n1110_94 vss 7.33536e-17
C1873 n1110_92 vss 7.33536e-17
C1874 n1110_103 vss 7.33536e-17
C1875 n1110_101 vss 7.33536e-17
C1876 n1110_112 vss 7.33536e-17
C1877 n1110_110 vss 7.33536e-17
C1878 n1110_67 vss 5.2569e-17
C1879 n1110_66 vss 5.2569e-17
C1880 n1110_85 vss 5.2569e-17
C1881 n1110_84 vss 5.2569e-17
C1882 n1110_76 vss 5.2569e-17
C1883 n1110_75 vss 5.2569e-17
C1884 n1110_94 vss 5.2569e-17
C1885 n1110_93 vss 5.2569e-17
C1886 n1110_103 vss 5.2569e-17
C1887 n1110_102 vss 5.2569e-17
C1888 n1110_112 vss 5.2569e-17
C1889 n1110_111 vss 5.2569e-17
C1890 n1110_27 vss 2.34738e-17
C1891 n1110_26 vss 2.34738e-17
C1892 n1110_29 vss 2.34738e-17
C1893 n1110_27 vss 2.34738e-17
C1894 n1110_30 vss 4.69476e-17
C1895 n1110_29 vss 4.69476e-17
C1896 n1110_31 vss 4.69476e-17
C1897 n1110_30 vss 4.69476e-17
C1898 n1110_33 vss 2.34738e-17
C1899 n1110_32 vss 2.34738e-17
C1900 n1110_35 vss 2.34738e-17
C1901 n1110_33 vss 2.34738e-17
C1902 n1110_36 vss 4.69476e-17
C1903 n1110_35 vss 4.69476e-17
C1904 n1110_37 vss 4.69476e-17
C1905 n1110_36 vss 4.69476e-17
C1906 n1110_39 vss 2.34738e-17
C1907 n1110_38 vss 2.34738e-17
C1908 n1110_41 vss 2.34738e-17
C1909 n1110_39 vss 2.34738e-17
C1910 n1110_42 vss 4.69476e-17
C1911 n1110_41 vss 4.69476e-17
C1912 n1110_43 vss 4.69476e-17
C1913 n1110_42 vss 4.69476e-17
C1914 n1110_45 vss 2.34738e-17
C1915 n1110_44 vss 2.34738e-17
C1916 n1110_47 vss 2.34738e-17
C1917 n1110_45 vss 2.34738e-17
C1918 n1110_48 vss 4.69476e-17
C1919 n1110_47 vss 4.69476e-17
C1920 n1110_49 vss 4.69476e-17
C1921 n1110_48 vss 4.69476e-17
C1922 n1110_51 vss 2.34738e-17
C1923 n1110_50 vss 2.34738e-17
C1924 n1110_53 vss 2.34738e-17
C1925 n1110_51 vss 2.34738e-17
C1926 n1110_54 vss 4.69476e-17
C1927 n1110_53 vss 4.69476e-17
C1928 n1110_55 vss 4.69476e-17
C1929 n1110_54 vss 4.69476e-17
C1930 n1110_57 vss 2.34738e-17
C1931 n1110_56 vss 2.34738e-17
C1932 n1110_59 vss 2.34738e-17
C1933 n1110_57 vss 2.34738e-17
C1934 n1110_60 vss 4.69476e-17
C1935 n1110_59 vss 4.69476e-17
C1936 n1110_61 vss 4.69476e-17
C1937 n1110_60 vss 4.69476e-17
C1938 n1110_28 vss 7.33536e-17
C1939 n1110_27 vss 7.33536e-17
C1940 n1110_34 vss 7.33536e-17
C1941 n1110_33 vss 7.33536e-17
C1942 n1110_40 vss 7.33536e-17
C1943 n1110_39 vss 7.33536e-17
C1944 n1110_46 vss 7.33536e-17
C1945 n1110_45 vss 7.33536e-17
C1946 n1110_52 vss 7.33536e-17
C1947 n1110_51 vss 7.33536e-17
C1948 n1110_58 vss 7.33536e-17
C1949 n1110_57 vss 7.33536e-17
C1950 n1110_63 vss 4.38566e-17
C1951 n1110_62 vss 4.38566e-17
C1952 n1110_81 vss 4.38566e-17
C1953 n1110_80 vss 4.38566e-17
C1954 n1110_72 vss 4.38566e-17
C1955 n1110_71 vss 4.38566e-17
C1956 n1110_90 vss 4.38566e-17
C1957 n1110_89 vss 4.38566e-17
C1958 n1110_99 vss 4.38566e-17
C1959 n1110_98 vss 4.38566e-17
C1960 n1110_108 vss 4.38566e-17
C1961 n1110_107 vss 4.38566e-17
C1962 n1110_124 vss 1.20606e-16
C1963 n1110_165 vss 1.20606e-16
C1964 n1110_125 vss 2.92378e-17
C1965 n1110_124 vss 2.92378e-17
C1966 n1110_126 vss 2.92378e-17
C1967 n1110_125 vss 2.92378e-17
C1968 n1110_127 vss 2.92378e-17
C1969 n1110_126 vss 2.92378e-17
C1970 n1110_128 vss 2.92378e-17
C1971 n1110_127 vss 2.92378e-17
C1972 n1110_129 vss 2.92378e-17
C1973 n1110_128 vss 2.92378e-17
C1974 n1110_130 vss 2.92378e-17
C1975 n1110_129 vss 2.92378e-17
C1976 n1110_131 vss 2.92378e-17
C1977 n1110_130 vss 2.92378e-17
C1978 n1110_132 vss 2.92378e-17
C1979 n1110_131 vss 2.92378e-17
C1980 n1110_133 vss 2.92378e-17
C1981 n1110_132 vss 2.92378e-17
C1982 n1110_134 vss 2.92378e-17
C1983 n1110_133 vss 2.92378e-17
C1984 n1110_135 vss 2.92378e-17
C1985 n1110_134 vss 2.92378e-17
C1986 n1110_136 vss 2.92378e-17
C1987 n1110_135 vss 2.92378e-17
C1988 n1110_137 vss 2.92378e-17
C1989 n1110_136 vss 2.92378e-17
C1990 n1110_138 vss 2.92378e-17
C1991 n1110_137 vss 2.92378e-17
C1992 n1110_139 vss 1.20606e-16
C1993 n1110_166 vss 1.20606e-16
C1994 n1110_140 vss 2.92378e-17
C1995 n1110_139 vss 2.92378e-17
C1996 n1110_141 vss 2.92378e-17
C1997 n1110_140 vss 2.92378e-17
C1998 n1110_142 vss 2.92378e-17
C1999 n1110_141 vss 2.92378e-17
C2000 n1110_143 vss 2.92378e-17
C2001 n1110_142 vss 2.92378e-17
C2002 n1110_144 vss 2.92378e-17
C2003 n1110_143 vss 2.92378e-17
C2004 n1110_145 vss 2.92378e-17
C2005 n1110_144 vss 2.92378e-17
C2006 n1110_146 vss 2.92378e-17
C2007 n1110_145 vss 2.92378e-17
C2008 n1110_147 vss 2.92378e-17
C2009 n1110_146 vss 2.92378e-17
C2010 n1110_148 vss 2.92378e-17
C2011 n1110_147 vss 2.92378e-17
C2012 n1110_149 vss 2.92378e-17
C2013 n1110_148 vss 2.92378e-17
C2014 n1110_150 vss 2.92378e-17
C2015 n1110_149 vss 2.92378e-17
C2016 n1110_151 vss 2.92378e-17
C2017 n1110_150 vss 2.92378e-17
C2018 n1110_152 vss 2.92378e-17
C2019 n1110_151 vss 2.92378e-17
C2020 n1110_153 vss 2.92378e-17
C2021 n1110_152 vss 2.92378e-17
C2022 n1110_117 vss 3.2562e-17
C2023 n1110_116 vss 3.2562e-17
C2024 n1110_118 vss 4.55868e-17
C2025 n1110_117 vss 4.55868e-17
C2026 n1110_119 vss 1.56298e-16
C2027 n1110_118 vss 1.56298e-16
C2028 n1110_120 vss 1.56298e-16
C2029 n1110_119 vss 1.56298e-16
C2030 n1110_121 vss 1.56298e-16
C2031 n1110_120 vss 1.56298e-16
C2032 n1110_122 vss 1.56298e-16
C2033 n1110_121 vss 1.56298e-16
C2034 n1110_123 vss 1.56298e-16
C2035 n1110_122 vss 1.56298e-16
C2036 n1110_162 vss 1.33073e-16
C2037 n1110_157 vss 1.33073e-16
C2038 n1110_163 vss 1.87868e-16
C2039 n1110_162 vss 1.87868e-16
C2040 n1110_164 vss 1.87868e-16
C2041 n1110_163 vss 1.87868e-16
C2042 n1110_165 vss 1.95696e-16
C2043 n1110_164 vss 1.95696e-16
C2044 n1110_166 vss 1.01762e-16
C2045 n1110_165 vss 1.01762e-16
C2046 n1110_167 vss 7.82784e-17
C2047 n1110_166 vss 7.82784e-17
C2048 n1110_168 vss 1.87868e-16
C2049 n1110_167 vss 1.87868e-16
C2050 n1110_169 vss 1.40901e-17
C2051 n1110_168 vss 1.40901e-17
C2052 n1110_154 vss 3.91392e-17
C2053 n1110_156 vss 3.91392e-17
C2054 n1110_155 vss 1.40901e-17
C2055 n1110_154 vss 1.40901e-17
C2056 n1110_3 vss 2.92378e-17
C2057 n1110_2 vss 2.92378e-17
C2058 n1110_4 vss 2.92378e-17
C2059 n1110_3 vss 2.92378e-17
C2060 n1110_5 vss 2.92378e-17
C2061 n1110_4 vss 2.92378e-17
C2062 n1110_6 vss 3.65472e-17
C2063 n1110_5 vss 3.65472e-17
C2064 n1110_7 vss 2.92378e-17
C2065 n1110_6 vss 2.92378e-17
C2066 n1110_8 vss 3.65472e-17
C2067 n1110_7 vss 3.65472e-17
C2068 n1110_9 vss 1.3157e-17
C2069 n1110_8 vss 1.3157e-17
C2070 n1110_157 vss 7.94526e-16
C2071 n1110_156 vss 7.94526e-16
C2072 n1110_158 vss 8.96288e-16
C2073 n1110_157 vss 8.96288e-16
C2074 n1110_159 vss 3.13114e-17
C2075 n1110_158 vss 3.13114e-17
C2076 n1110_160 vss 3.13114e-17
C2077 n1110_159 vss 3.13114e-17
C2078 n1110_161 vss 1.40901e-17
C2079 n1110_160 vss 1.40901e-17
C2080 n1110_20 vss 2.60496e-17
C2081 n1110_19 vss 2.60496e-17
C2082 n1110_21 vss 2.60496e-17
C2083 n1110_20 vss 2.60496e-17
C2084 n1110_22 vss 5.40529e-16
C2085 n1110_21 vss 5.40529e-16
C2086 n1110_23 vss 7.81488e-17
C2087 n1110_22 vss 7.81488e-17
C2088 n1110_12 vss 2.92378e-17
C2089 n1110_11 vss 2.92378e-17
C2090 n1110_13 vss 2.92378e-17
C2091 n1110_12 vss 2.92378e-17
C2092 n1110_14 vss 2.92378e-17
C2093 n1110_13 vss 2.92378e-17
C2094 n1110_15 vss 3.65472e-17
C2095 n1110_14 vss 3.65472e-17
C2096 n1110_16 vss 2.92378e-17
C2097 n1110_15 vss 2.92378e-17
C2098 n1110_17 vss 3.65472e-17
C2099 n1110_16 vss 3.65472e-17
C2100 n1110_18 vss 1.3157e-17
C2101 n1110_17 vss 1.3157e-17

R45_1 n1191 n1191_27 0.001
R45_2 n1191 n1191_28 0.001
R45_3 n1191 n1191_26 0.001
R45_4 n1191 n1191_23 0.001
R45_5 n1191 n1191_22 0.001
R45_6 n1191 n1191_24 0.001
R45_7 n1191 n1191_25 0.001
R45_8 n1191_20 n1191_5 0.001
R45_9 n1191_21 n1191_4 0.001
R45_10 n1191_18 n1191_5 0.001
R45_11 n1191_19 n1191_5 0.001
R45_12 n1191_16 n1191_5 0.001
R45_13 n1191_17 n1191_5 0.001
R45_14 n1191_13 n1191_5 0.001
R45_15 n1191_15 n1191_5 0.001
R45_16 n1191_14 n1191_5 0.001
R45_17 n1191_10 n1191_5 0.001
R45_18 n1191_12 n1191_5 0.001
R45_19 n1191_11 n1191_5 0.001
R45_20 n1191_7 n1191_5 0.001
R45_21 n1191_8 n1191_5 0.001
R45_22 n1191_6 n1191_5 0.001
R45_23 n1191_9 n1191_5 0.001
R45_24 n1191_2 n1191_3 453.6
R45_25 n1191_4 n1191_3 14.4
R45_26 n1191_7 n1191_6 0.108
R45_27 n1191_8 n1191_7 0.108
R45_28 n1191_9 n1191_8 0.108
R45_29 n1191_10 n1191_9 0.108
R45_30 n1191_11 n1191_10 0.108
R45_31 n1191_12 n1191_11 0.108
R45_32 n1191_13 n1191_12 0.108
R45_33 n1191_14 n1191_13 0.108
R45_34 n1191_15 n1191_14 0.108
R45_35 n1191_16 n1191_15 0.108
R45_36 n1191_17 n1191_16 0.108
R45_37 n1191_18 n1191_17 0.108
R45_38 n1191_19 n1191_18 0.108
R45_39 n1191_20 n1191_19 0.108
R45_40 n1191_21 n1191_20 0.108
R45_41 n1191_22 n1191_21 0.756
R45_42 n1191_23 n1191_22 0.108
R45_43 n1191_24 n1191_23 0.108
R45_44 n1191_25 n1191_24 0.108
R45_45 n1191_26 n1191_25 0.108
R45_46 n1191_27 n1191_26 0.108
R45_47 n1191_28 n1191_27 0.108

C2102 n1191_2 vss 4.98819e-16
C2103 n1191_3 vss 4.98819e-16
C2104 n1191_4 vss 8.41104e-17
C2105 n1191_3 vss 8.41104e-17
C2106 n1191_7 vss 2.92378e-17
C2107 n1191_6 vss 2.92378e-17
C2108 n1191_8 vss 2.92378e-17
C2109 n1191_7 vss 2.92378e-17
C2110 n1191_9 vss 2.92378e-17
C2111 n1191_8 vss 2.92378e-17
C2112 n1191_10 vss 2.92378e-17
C2113 n1191_9 vss 2.92378e-17
C2114 n1191_11 vss 2.92378e-17
C2115 n1191_10 vss 2.92378e-17
C2116 n1191_12 vss 2.92378e-17
C2117 n1191_11 vss 2.92378e-17
C2118 n1191_13 vss 2.92378e-17
C2119 n1191_12 vss 2.92378e-17
C2120 n1191_14 vss 2.92378e-17
C2121 n1191_13 vss 2.92378e-17
C2122 n1191_15 vss 2.92378e-17
C2123 n1191_14 vss 2.92378e-17
C2124 n1191_16 vss 2.92378e-17
C2125 n1191_15 vss 2.92378e-17
C2126 n1191_17 vss 2.92378e-17
C2127 n1191_16 vss 2.92378e-17
C2128 n1191_18 vss 2.92378e-17
C2129 n1191_17 vss 2.92378e-17
C2130 n1191_19 vss 2.92378e-17
C2131 n1191_18 vss 2.92378e-17
C2132 n1191_20 vss 2.92378e-17
C2133 n1191_19 vss 2.92378e-17
C2134 n1191_21 vss 3.65472e-17
C2135 n1191_20 vss 3.65472e-17
C2136 n1191_22 vss 1.46189e-16
C2137 n1191_21 vss 1.46189e-16
C2138 n1191_23 vss 2.92378e-17
C2139 n1191_22 vss 2.92378e-17
C2140 n1191_24 vss 2.92378e-17
C2141 n1191_23 vss 2.92378e-17
C2142 n1191_25 vss 2.92378e-17
C2143 n1191_24 vss 2.92378e-17
C2144 n1191_26 vss 2.92378e-17
C2145 n1191_25 vss 2.92378e-17
C2146 n1191_27 vss 2.92378e-17
C2147 n1191_26 vss 2.92378e-17
C2148 n1191_28 vss 2.92378e-17
C2149 n1191_27 vss 2.92378e-17

R46_1 n1228 n1228_35 0.001
R46_2 n1228 n1228_36 0.001
R46_3 n1228 n1228_37 0.001
R46_4 n1228 n1228_32 0.001
R46_5 n1228 n1228_31 0.001
R46_6 n1228 n1228_33 0.001
R46_7 n1228 n1228_34 0.001
R46_8 n1228_14 n1228_11 0.001
R46_9 n1228_29 n1228_13 0.001
R46_10 n1228_26 n1228_13 0.001
R46_11 n1228_27 n1228_13 0.001
R46_12 n1228_28 n1228_13 0.001
R46_13 n1228_25 n1228_13 0.001
R46_14 n1228_22 n1228_13 0.001
R46_15 n1228_23 n1228_13 0.001
R46_16 n1228_24 n1228_13 0.001
R46_17 n1228_21 n1228_13 0.001
R46_18 n1228_19 n1228_13 0.001
R46_19 n1228_20 n1228_13 0.001
R46_20 n1228_18 n1228_13 0.001
R46_21 n1228_17 n1228_13 0.001
R46_22 n1228_16 n1228_13 0.001
R46_23 n1228_15 n1228_13 0.001
R46_24 n1228_3 n1228_2 43.2
R46_25 n1228_12 n1228_3 21.6
R46_26 n1228_4 n1228_12 21.6
R46_27 n1228_5 n1228_4 43.2
R46_28 n1228_7 n1228_6 43.2
R46_29 n1228_10 n1228_7 21.6
R46_30 n1228_8 n1228_10 21.6
R46_31 n1228_9 n1228_8 43.2
R46_32 n1228_11 n1228_10 28.8
R46_33 n1228_12 n1228_11 28.8
R46_34 n1228_30 n1228_14 0.648
R46_35 n1228_16 n1228_15 0.108
R46_36 n1228_17 n1228_16 0.108
R46_37 n1228_18 n1228_17 0.108
R46_38 n1228_19 n1228_18 0.108
R46_39 n1228_20 n1228_19 0.108
R46_40 n1228_21 n1228_20 0.108
R46_41 n1228_22 n1228_21 0.108
R46_42 n1228_23 n1228_22 0.108
R46_43 n1228_24 n1228_23 0.108
R46_44 n1228_25 n1228_24 0.108
R46_45 n1228_26 n1228_25 0.108
R46_46 n1228_27 n1228_26 0.108
R46_47 n1228_28 n1228_27 0.108
R46_48 n1228_29 n1228_28 0.108
R46_49 n1228_30 n1228_29 0.432
R46_50 n1228_31 n1228_30 0.54
R46_51 n1228_32 n1228_31 0.108
R46_52 n1228_33 n1228_32 0.108
R46_53 n1228_34 n1228_33 0.108
R46_54 n1228_35 n1228_34 0.108
R46_55 n1228_36 n1228_35 0.108
R46_56 n1228_37 n1228_36 0.108

C2150 n1228_3 vss 4.69476e-17
C2151 n1228_2 vss 4.69476e-17
C2152 n1228_12 vss 2.34738e-17
C2153 n1228_3 vss 2.34738e-17
C2154 n1228_4 vss 2.34738e-17
C2155 n1228_12 vss 2.34738e-17
C2156 n1228_5 vss 4.69476e-17
C2157 n1228_4 vss 4.69476e-17
C2158 n1228_7 vss 4.69476e-17
C2159 n1228_6 vss 4.69476e-17
C2160 n1228_10 vss 2.34738e-17
C2161 n1228_7 vss 2.34738e-17
C2162 n1228_8 vss 2.34738e-17
C2163 n1228_10 vss 2.34738e-17
C2164 n1228_9 vss 4.69476e-17
C2165 n1228_8 vss 4.69476e-17
C2166 n1228_11 vss 7.33536e-17
C2167 n1228_10 vss 7.33536e-17
C2168 n1228_12 vss 8.25228e-17
C2169 n1228_11 vss 8.25228e-17
C2170 n1228_30 vss 1.3157e-16
C2171 n1228_14 vss 1.3157e-16
C2172 n1228_16 vss 2.92378e-17
C2173 n1228_15 vss 2.92378e-17
C2174 n1228_17 vss 2.92378e-17
C2175 n1228_16 vss 2.92378e-17
C2176 n1228_18 vss 2.92378e-17
C2177 n1228_17 vss 2.92378e-17
C2178 n1228_19 vss 2.92378e-17
C2179 n1228_18 vss 2.92378e-17
C2180 n1228_20 vss 2.92378e-17
C2181 n1228_19 vss 2.92378e-17
C2182 n1228_21 vss 2.92378e-17
C2183 n1228_20 vss 2.92378e-17
C2184 n1228_22 vss 2.92378e-17
C2185 n1228_21 vss 2.92378e-17
C2186 n1228_23 vss 2.92378e-17
C2187 n1228_22 vss 2.92378e-17
C2188 n1228_24 vss 2.92378e-17
C2189 n1228_23 vss 2.92378e-17
C2190 n1228_25 vss 2.92378e-17
C2191 n1228_24 vss 2.92378e-17
C2192 n1228_26 vss 2.92378e-17
C2193 n1228_25 vss 2.92378e-17
C2194 n1228_27 vss 2.92378e-17
C2195 n1228_26 vss 2.92378e-17
C2196 n1228_28 vss 2.92378e-17
C2197 n1228_27 vss 2.92378e-17
C2198 n1228_29 vss 2.92378e-17
C2199 n1228_28 vss 2.92378e-17
C2200 n1228_30 vss 8.77133e-17
C2201 n1228_29 vss 8.77133e-17
C2202 n1228_31 vss 9.50227e-17
C2203 n1228_30 vss 9.50227e-17
C2204 n1228_32 vss 2.92378e-17
C2205 n1228_31 vss 2.92378e-17
C2206 n1228_33 vss 2.92378e-17
C2207 n1228_32 vss 2.92378e-17
C2208 n1228_34 vss 2.92378e-17
C2209 n1228_33 vss 2.92378e-17
C2210 n1228_35 vss 2.92378e-17
C2211 n1228_34 vss 2.92378e-17
C2212 n1228_36 vss 2.92378e-17
C2213 n1228_35 vss 2.92378e-17
C2214 n1228_37 vss 2.92378e-17
C2215 n1228_36 vss 2.92378e-17

R47_1 b_3_2 b_3_84 0.001
R47_2 b_3_82 b_3_5 0.001
R47_3 b_3_42 b_3_7 0.001
R47_4 b_3_74 b_3_8 0.001
R47_5 b_3_40 b_3_7 0.001
R47_6 b_3_41 b_3_7 0.001
R47_7 b_3_72 b_3_8 0.001
R47_8 b_3_73 b_3_8 0.001
R47_9 b_3_38 b_3_7 0.001
R47_10 b_3_39 b_3_7 0.001
R47_11 b_3_71 b_3_8 0.001
R47_12 b_3_70 b_3_8 0.001
R47_13 b_3_37 b_3_7 0.001
R47_14 b_3_36 b_3_7 0.001
R47_15 b_3_68 b_3_8 0.001
R47_16 b_3_69 b_3_8 0.001
R47_17 b_3_34 b_3_7 0.001
R47_18 b_3_35 b_3_7 0.001
R47_19 b_3_67 b_3_8 0.001
R47_20 b_3_66 b_3_8 0.001
R47_21 b_3_32 b_3_7 0.001
R47_22 b_3_33 b_3_7 0.001
R47_23 b_3_64 b_3_8 0.001
R47_24 b_3_65 b_3_8 0.001
R47_25 b_3_30 b_3_7 0.001
R47_26 b_3_31 b_3_7 0.001
R47_27 b_3_63 b_3_8 0.001
R47_28 b_3_62 b_3_8 0.001
R47_29 b_3_29 b_3_7 0.001
R47_30 b_3_28 b_3_7 0.001
R47_31 b_3_60 b_3_8 0.001
R47_32 b_3_61 b_3_8 0.001
R47_33 b_3_27 b_3_7 0.001
R47_34 b_3_26 b_3_7 0.001
R47_35 b_3_59 b_3_8 0.001
R47_36 b_3_58 b_3_8 0.001
R47_37 b_3_24 b_3_7 0.001
R47_38 b_3_25 b_3_7 0.001
R47_39 b_3_57 b_3_8 0.001
R47_40 b_3_56 b_3_8 0.001
R47_41 b_3_23 b_3_7 0.001
R47_42 b_3_55 b_3_8 0.001
R47_43 b_3_22 b_3_9 0.001
R47_44 b_3_54 b_3_10 0.001
R47_45 b_3_21 b_3_9 0.001
R47_46 b_3_20 b_3_9 0.001
R47_47 b_3_53 b_3_10 0.001
R47_48 b_3_52 b_3_10 0.001
R47_49 b_3_18 b_3_9 0.001
R47_50 b_3_19 b_3_9 0.001
R47_51 b_3_51 b_3_10 0.001
R47_52 b_3_50 b_3_10 0.001
R47_53 b_3_16 b_3_9 0.001
R47_54 b_3_17 b_3_9 0.001
R47_55 b_3_48 b_3_10 0.001
R47_56 b_3_49 b_3_10 0.001
R47_57 b_3_15 b_3_9 0.001
R47_58 b_3_47 b_3_10 0.001
R47_59 b_3 b_3_11 0.001
R47_60 b_3 b_3_13 0.001
R47_61 b_3_14 b_3_13 0.001
R47_62 b_3_46 b_3_14 0.54
R47_63 b_3_15 b_3_45 0.54
R47_64 b_3_16 b_3_15 0.108
R47_65 b_3_17 b_3_16 0.108
R47_66 b_3_18 b_3_17 0.108
R47_67 b_3_19 b_3_18 0.108
R47_68 b_3_20 b_3_19 0.108
R47_69 b_3_21 b_3_20 0.108
R47_70 b_3_22 b_3_21 0.108
R47_71 b_3_23 b_3_22 0.864
R47_72 b_3_24 b_3_23 0.108
R47_73 b_3_25 b_3_24 0.108
R47_74 b_3_26 b_3_25 0.108
R47_75 b_3_27 b_3_26 0.108
R47_76 b_3_28 b_3_27 0.108
R47_77 b_3_29 b_3_28 0.108
R47_78 b_3_30 b_3_29 0.108
R47_79 b_3_31 b_3_30 0.108
R47_80 b_3_32 b_3_31 0.108
R47_81 b_3_33 b_3_32 0.108
R47_82 b_3_34 b_3_33 0.108
R47_83 b_3_35 b_3_34 0.108
R47_84 b_3_36 b_3_35 0.108
R47_85 b_3_37 b_3_36 0.108
R47_86 b_3_38 b_3_37 0.108
R47_87 b_3_39 b_3_38 0.108
R47_88 b_3_40 b_3_39 0.108
R47_89 b_3_41 b_3_40 0.108
R47_90 b_3_42 b_3_41 0.108
R47_91 b_3_43 b_3_42 0.001
R47_92 b_3_46 b_3_44 0.001
R47_93 b_3_45 b_3_46 0.108
R47_94 b_3_47 b_3_46 0.54
R47_95 b_3_48 b_3_47 0.108
R47_96 b_3_49 b_3_48 0.108
R47_97 b_3_50 b_3_49 0.108
R47_98 b_3_51 b_3_50 0.108
R47_99 b_3_52 b_3_51 0.108
R47_100 b_3_53 b_3_52 0.108
R47_101 b_3_54 b_3_53 0.108
R47_102 b_3_55 b_3_54 0.864
R47_103 b_3_56 b_3_55 0.108
R47_104 b_3_57 b_3_56 0.108
R47_105 b_3_58 b_3_57 0.108
R47_106 b_3_59 b_3_58 0.108
R47_107 b_3_60 b_3_59 0.108
R47_108 b_3_61 b_3_60 0.108
R47_109 b_3_62 b_3_61 0.108
R47_110 b_3_63 b_3_62 0.108
R47_111 b_3_64 b_3_63 0.108
R47_112 b_3_65 b_3_64 0.108
R47_113 b_3_66 b_3_65 0.108
R47_114 b_3_67 b_3_66 0.108
R47_115 b_3_68 b_3_67 0.108
R47_116 b_3_69 b_3_68 0.108
R47_117 b_3_70 b_3_69 0.108
R47_118 b_3_71 b_3_70 0.108
R47_119 b_3_72 b_3_71 0.108
R47_120 b_3_73 b_3_72 0.108
R47_121 b_3_74 b_3_73 0.108
R47_122 b_3_75 b_3_74 0.001
R47_123 b_3_76 b_3_75 0.216
R47_124 b_3_77 b_3_76 0.001
R47_125 b_3_78 b_3_77 0.001
R47_126 b_3_78 b_3_79 1.08
R47_127 b_3_80 b_3_79 2.268
R47_128 b_3_6 b_3_5 21.6
R47_129 b_3_83 b_3_80 0.324
R47_130 b_3_82 b_3_81 0.001
R47_131 b_3_83 b_3_82 0.216
R47_132 b_3_84 b_3_83 0.216
R47_133 b_3_85 b_3_84 0.001
R47_134 b_3_1 b_3_2 7.2
R47_135 b_3_3 b_3_2 7.2
R47_136 b_3_4 b_3_3 14.4

C2216 b_3 vss 4.3846e-15
C2217 b_3_13 vss 4.3846e-15
C2218 b_3_14 vss 3.48676e-17
C2219 b_3_13 vss 3.48676e-17
C2220 b_3_46 vss 6.8969e-16
C2221 b_3_14 vss 6.8969e-16
C2222 b_3_15 vss 1.40901e-16
C2223 b_3_45 vss 1.40901e-16
C2224 b_3_16 vss 3.13114e-17
C2225 b_3_15 vss 3.13114e-17
C2226 b_3_17 vss 3.13114e-17
C2227 b_3_16 vss 3.13114e-17
C2228 b_3_18 vss 3.13114e-17
C2229 b_3_17 vss 3.13114e-17
C2230 b_3_19 vss 3.13114e-17
C2231 b_3_18 vss 3.13114e-17
C2232 b_3_20 vss 3.13114e-17
C2233 b_3_19 vss 3.13114e-17
C2234 b_3_21 vss 3.13114e-17
C2235 b_3_20 vss 3.13114e-17
C2236 b_3_22 vss 3.13114e-17
C2237 b_3_21 vss 3.13114e-17
C2238 b_3_23 vss 2.42663e-16
C2239 b_3_22 vss 2.42663e-16
C2240 b_3_24 vss 3.13114e-17
C2241 b_3_23 vss 3.13114e-17
C2242 b_3_25 vss 3.13114e-17
C2243 b_3_24 vss 3.13114e-17
C2244 b_3_26 vss 3.13114e-17
C2245 b_3_25 vss 3.13114e-17
C2246 b_3_27 vss 3.13114e-17
C2247 b_3_26 vss 3.13114e-17
C2248 b_3_28 vss 3.13114e-17
C2249 b_3_27 vss 3.13114e-17
C2250 b_3_29 vss 3.13114e-17
C2251 b_3_28 vss 3.13114e-17
C2252 b_3_30 vss 3.13114e-17
C2253 b_3_29 vss 3.13114e-17
C2254 b_3_31 vss 3.13114e-17
C2255 b_3_30 vss 3.13114e-17
C2256 b_3_32 vss 3.13114e-17
C2257 b_3_31 vss 3.13114e-17
C2258 b_3_33 vss 3.13114e-17
C2259 b_3_32 vss 3.13114e-17
C2260 b_3_34 vss 3.13114e-17
C2261 b_3_33 vss 3.13114e-17
C2262 b_3_35 vss 3.13114e-17
C2263 b_3_34 vss 3.13114e-17
C2264 b_3_36 vss 3.13114e-17
C2265 b_3_35 vss 3.13114e-17
C2266 b_3_37 vss 3.13114e-17
C2267 b_3_36 vss 3.13114e-17
C2268 b_3_38 vss 3.13114e-17
C2269 b_3_37 vss 3.13114e-17
C2270 b_3_39 vss 3.13114e-17
C2271 b_3_38 vss 3.13114e-17
C2272 b_3_40 vss 3.13114e-17
C2273 b_3_39 vss 3.13114e-17
C2274 b_3_41 vss 3.13114e-17
C2275 b_3_40 vss 3.13114e-17
C2276 b_3_42 vss 3.13114e-17
C2277 b_3_41 vss 3.13114e-17
C2278 b_3_43 vss 1.40901e-17
C2279 b_3_42 vss 1.40901e-17
C2280 b_3_46 vss 6.34418e-17
C2281 b_3_44 vss 6.34418e-17
C2282 b_3_45 vss 1.42197e-16
C2283 b_3_46 vss 1.42197e-16
C2284 b_3_47 vss 1.40901e-16
C2285 b_3_46 vss 1.40901e-16
C2286 b_3_48 vss 3.13114e-17
C2287 b_3_47 vss 3.13114e-17
C2288 b_3_49 vss 3.13114e-17
C2289 b_3_48 vss 3.13114e-17
C2290 b_3_50 vss 3.13114e-17
C2291 b_3_49 vss 3.13114e-17
C2292 b_3_51 vss 3.13114e-17
C2293 b_3_50 vss 3.13114e-17
C2294 b_3_52 vss 3.13114e-17
C2295 b_3_51 vss 3.13114e-17
C2296 b_3_53 vss 3.13114e-17
C2297 b_3_52 vss 3.13114e-17
C2298 b_3_54 vss 3.13114e-17
C2299 b_3_53 vss 3.13114e-17
C2300 b_3_55 vss 2.42663e-16
C2301 b_3_54 vss 2.42663e-16
C2302 b_3_56 vss 3.13114e-17
C2303 b_3_55 vss 3.13114e-17
C2304 b_3_57 vss 3.13114e-17
C2305 b_3_56 vss 3.13114e-17
C2306 b_3_58 vss 3.13114e-17
C2307 b_3_57 vss 3.13114e-17
C2308 b_3_59 vss 3.13114e-17
C2309 b_3_58 vss 3.13114e-17
C2310 b_3_60 vss 3.13114e-17
C2311 b_3_59 vss 3.13114e-17
C2312 b_3_61 vss 3.13114e-17
C2313 b_3_60 vss 3.13114e-17
C2314 b_3_62 vss 3.13114e-17
C2315 b_3_61 vss 3.13114e-17
C2316 b_3_63 vss 3.13114e-17
C2317 b_3_62 vss 3.13114e-17
C2318 b_3_64 vss 3.13114e-17
C2319 b_3_63 vss 3.13114e-17
C2320 b_3_65 vss 3.13114e-17
C2321 b_3_64 vss 3.13114e-17
C2322 b_3_66 vss 3.13114e-17
C2323 b_3_65 vss 3.13114e-17
C2324 b_3_67 vss 3.13114e-17
C2325 b_3_66 vss 3.13114e-17
C2326 b_3_68 vss 3.13114e-17
C2327 b_3_67 vss 3.13114e-17
C2328 b_3_69 vss 3.13114e-17
C2329 b_3_68 vss 3.13114e-17
C2330 b_3_70 vss 3.13114e-17
C2331 b_3_69 vss 3.13114e-17
C2332 b_3_71 vss 3.13114e-17
C2333 b_3_70 vss 3.13114e-17
C2334 b_3_72 vss 3.13114e-17
C2335 b_3_71 vss 3.13114e-17
C2336 b_3_73 vss 3.13114e-17
C2337 b_3_72 vss 3.13114e-17
C2338 b_3_74 vss 3.13114e-17
C2339 b_3_73 vss 3.13114e-17
C2340 b_3_75 vss 1.40901e-17
C2341 b_3_74 vss 1.40901e-17
C2342 b_3_76 vss 8.14095e-17
C2343 b_3_75 vss 8.14095e-17
C2344 b_3_77 vss 1.25245e-17
C2345 b_3_76 vss 1.25245e-17
C2346 b_3_78 vss 2.50491e-17
C2347 b_3_77 vss 2.50491e-17
C2348 b_3_78 vss 2.97458e-16
C2349 b_3_79 vss 2.97458e-16
C2350 b_3_80 vss 6.18399e-16
C2351 b_3_79 vss 6.18399e-16
C2352 b_3_6 vss 9.46242e-17
C2353 b_3_5 vss 9.46242e-17
C2354 b_3_83 vss 9.39341e-17
C2355 b_3_80 vss 9.39341e-17
C2356 b_3_82 vss 1.40901e-17
C2357 b_3_81 vss 1.40901e-17
C2358 b_3_83 vss 7.04506e-17
C2359 b_3_82 vss 7.04506e-17
C2360 b_3_84 vss 7.82784e-17
C2361 b_3_83 vss 7.82784e-17
C2362 b_3_85 vss 1.40901e-17
C2363 b_3_84 vss 1.40901e-17
C2364 b_3_1 vss 3.15414e-17
C2365 b_3_2 vss 3.15414e-17
C2366 b_3_3 vss 3.15414e-17
C2367 b_3_2 vss 3.15414e-17
C2368 b_3_4 vss 6.30828e-17
C2369 b_3_3 vss 6.30828e-17

R48_1 n1367_7 n1367_39 0.001
R48_2 n1367_38 n1367_2 0.001
R48_3 n1367_1 n1367_18 0.001
R48_4 n1367_19 n1367_8 0.001
R48_5 n1367_7 n1367_36 0.001
R48_6 n1367_7 n1367_37 0.001
R48_7 n1367_16 n1367_8 0.001
R48_8 n1367_17 n1367_8 0.001
R48_9 n1367_23 n1367_4 0.001
R48_10 n1367_34 n1367_3 0.001
R48_11 n1367_7 n1367_35 0.001
R48_12 n1367_15 n1367_8 0.001
R48_13 n1367_20 n1367_10 0.001
R48_14 n1367_31 n1367_9 0.001
R48_15 n1367_30 n1367_13 0.001
R48_16 n1367_29 n1367_13 0.001
R48_17 n1367_28 n1367_13 0.001
R48_18 n1367_27 n1367_13 0.001
R48_19 n1367_26 n1367_13 0.001
R48_20 n1367_10 n1367_9 7.2
R48_21 n1367_11 n1367_10 21.6
R48_22 n1367_12 n1367_11 0.001
R48_23 n1367_15 n1367_14 0.001
R48_24 n1367_16 n1367_15 0.108
R48_25 n1367_17 n1367_16 0.108
R48_26 n1367_18 n1367_17 0.108
R48_27 n1367_19 n1367_18 0.108
R48_28 n1367_22 n1367_19 0.324
R48_29 n1367_2 n1367_1 0.216
R48_30 n1367_20 n1367_31 0.108
R48_31 n1367_21 n1367_20 0.001
R48_32 n1367_4 n1367_3 7.2
R48_33 n1367_5 n1367_4 21.6
R48_34 n1367 n1367_5 0.001
R48_35 n1367_40 n1367_22 0.324
R48_36 n1367_23 n1367_34 0.108
R48_37 n1367_24 n1367_23 0.001
R48_38 n1367_26 n1367_25 0.001
R48_39 n1367_27 n1367_26 0.108
R48_40 n1367_28 n1367_27 0.108
R48_41 n1367_29 n1367_28 0.108
R48_42 n1367_30 n1367_29 0.108
R48_43 n1367_31 n1367_30 0.108
R48_44 n1367_32 n1367_31 0.216
R48_45 n1367_33 n1367_32 0.108
R48_46 n1367_34 n1367_33 0.216
R48_47 n1367_35 n1367_34 0.108
R48_48 n1367_36 n1367_35 0.108
R48_49 n1367_37 n1367_36 0.108
R48_50 n1367_38 n1367_37 0.108
R48_51 n1367_39 n1367_38 0.108
R48_52 n1367_40 n1367_39 0.324

C2370 n1367_10 vss 4.20552e-17
C2371 n1367_9 vss 4.20552e-17
C2372 n1367_11 vss 9.46242e-17
C2373 n1367_10 vss 9.46242e-17
C2374 n1367_12 vss 5.47139e-16
C2375 n1367_11 vss 5.47139e-16
C2376 n1367_15 vss 1.40901e-17
C2377 n1367_14 vss 1.40901e-17
C2378 n1367_16 vss 3.91392e-17
C2379 n1367_15 vss 3.91392e-17
C2380 n1367_17 vss 3.91392e-17
C2381 n1367_16 vss 3.91392e-17
C2382 n1367_18 vss 3.91392e-17
C2383 n1367_17 vss 3.91392e-17
C2384 n1367_19 vss 3.91392e-17
C2385 n1367_18 vss 3.91392e-17
C2386 n1367_22 vss 1.0959e-16
C2387 n1367_19 vss 1.0959e-16
C2388 n1367_2 vss 7.81488e-17
C2389 n1367_1 vss 7.81488e-17
C2390 n1367_20 vss 3.71822e-17
C2391 n1367_31 vss 3.71822e-17
C2392 n1367_21 vss 1.40901e-17
C2393 n1367_20 vss 1.40901e-17
C2394 n1367_4 vss 4.20552e-17
C2395 n1367_3 vss 4.20552e-17
C2396 n1367_5 vss 9.46242e-17
C2397 n1367_4 vss 9.46242e-17
C2398 n1367 vss 3.05111e-16
C2399 n1367_5 vss 3.05111e-16
C2400 n1367_40 vss 9.39341e-17
C2401 n1367_22 vss 9.39341e-17
C2402 n1367_23 vss 3.71822e-17
C2403 n1367_34 vss 3.71822e-17
C2404 n1367_24 vss 1.40901e-17
C2405 n1367_23 vss 1.40901e-17
C2406 n1367_26 vss 1.40901e-17
C2407 n1367_25 vss 1.40901e-17
C2408 n1367_27 vss 3.91392e-17
C2409 n1367_26 vss 3.91392e-17
C2410 n1367_28 vss 3.91392e-17
C2411 n1367_27 vss 3.91392e-17
C2412 n1367_29 vss 4.6967e-17
C2413 n1367_28 vss 4.6967e-17
C2414 n1367_30 vss 3.91392e-17
C2415 n1367_29 vss 3.91392e-17
C2416 n1367_31 vss 4.6967e-17
C2417 n1367_30 vss 4.6967e-17
C2418 n1367_32 vss 6.41883e-17
C2419 n1367_31 vss 6.41883e-17
C2420 n1367_33 vss 2.81802e-17
C2421 n1367_32 vss 2.81802e-17
C2422 n1367_34 vss 5.63604e-17
C2423 n1367_33 vss 5.63604e-17
C2424 n1367_35 vss 4.6967e-17
C2425 n1367_34 vss 4.6967e-17
C2426 n1367_36 vss 3.91392e-17
C2427 n1367_35 vss 3.91392e-17
C2428 n1367_37 vss 3.91392e-17
C2429 n1367_36 vss 3.91392e-17
C2430 n1367_38 vss 3.91392e-17
C2431 n1367_37 vss 3.91392e-17
C2432 n1367_39 vss 3.91392e-17
C2433 n1367_38 vss 3.91392e-17
C2434 n1367_40 vss 1.0959e-16
C2435 n1367_39 vss 1.0959e-16

R49_1 b_2_2 b_2_84 0.001
R49_2 b_2_82 b_2_5 0.001
R49_3 b_2_40 b_2_7 0.001
R49_4 b_2_74 b_2_8 0.001
R49_5 b_2_38 b_2_7 0.001
R49_6 b_2_39 b_2_7 0.001
R49_7 b_2_72 b_2_8 0.001
R49_8 b_2_73 b_2_8 0.001
R49_9 b_2_37 b_2_7 0.001
R49_10 b_2_36 b_2_7 0.001
R49_11 b_2_71 b_2_8 0.001
R49_12 b_2_70 b_2_8 0.001
R49_13 b_2_34 b_2_7 0.001
R49_14 b_2_35 b_2_7 0.001
R49_15 b_2_68 b_2_8 0.001
R49_16 b_2_69 b_2_8 0.001
R49_17 b_2_33 b_2_7 0.001
R49_18 b_2_32 b_2_7 0.001
R49_19 b_2_67 b_2_8 0.001
R49_20 b_2_66 b_2_8 0.001
R49_21 b_2_30 b_2_7 0.001
R49_22 b_2_31 b_2_7 0.001
R49_23 b_2_64 b_2_8 0.001
R49_24 b_2_65 b_2_8 0.001
R49_25 b_2_28 b_2_7 0.001
R49_26 b_2_29 b_2_7 0.001
R49_27 b_2_62 b_2_8 0.001
R49_28 b_2_63 b_2_8 0.001
R49_29 b_2_27 b_2_7 0.001
R49_30 b_2_26 b_2_7 0.001
R49_31 b_2_60 b_2_8 0.001
R49_32 b_2_61 b_2_8 0.001
R49_33 b_2_25 b_2_7 0.001
R49_34 b_2_24 b_2_7 0.001
R49_35 b_2_58 b_2_8 0.001
R49_36 b_2_59 b_2_8 0.001
R49_37 b_2_22 b_2_7 0.001
R49_38 b_2_23 b_2_7 0.001
R49_39 b_2_56 b_2_8 0.001
R49_40 b_2_57 b_2_8 0.001
R49_41 b_2_21 b_2_7 0.001
R49_42 b_2_55 b_2_8 0.001
R49_43 b_2_20 b_2_9 0.001
R49_44 b_2_54 b_2_10 0.001
R49_45 b_2_18 b_2_9 0.001
R49_46 b_2_19 b_2_9 0.001
R49_47 b_2_53 b_2_10 0.001
R49_48 b_2_52 b_2_10 0.001
R49_49 b_2_17 b_2_9 0.001
R49_50 b_2_16 b_2_9 0.001
R49_51 b_2_51 b_2_10 0.001
R49_52 b_2_50 b_2_10 0.001
R49_53 b_2_14 b_2_9 0.001
R49_54 b_2_15 b_2_9 0.001
R49_55 b_2_48 b_2_10 0.001
R49_56 b_2_49 b_2_10 0.001
R49_57 b_2_13 b_2_9 0.001
R49_58 b_2_47 b_2_10 0.001
R49_59 b_2 b_2_11 0.001
R49_60 b_2 b_2_42 0.001
R49_61 b_2_13 b_2_45 0.54
R49_62 b_2_14 b_2_13 0.108
R49_63 b_2_15 b_2_14 0.108
R49_64 b_2_16 b_2_15 0.108
R49_65 b_2_17 b_2_16 0.108
R49_66 b_2_18 b_2_17 0.108
R49_67 b_2_19 b_2_18 0.108
R49_68 b_2_20 b_2_19 0.108
R49_69 b_2_21 b_2_20 0.864
R49_70 b_2_22 b_2_21 0.108
R49_71 b_2_23 b_2_22 0.108
R49_72 b_2_24 b_2_23 0.108
R49_73 b_2_25 b_2_24 0.108
R49_74 b_2_26 b_2_25 0.108
R49_75 b_2_27 b_2_26 0.108
R49_76 b_2_28 b_2_27 0.108
R49_77 b_2_29 b_2_28 0.108
R49_78 b_2_30 b_2_29 0.108
R49_79 b_2_31 b_2_30 0.108
R49_80 b_2_32 b_2_31 0.108
R49_81 b_2_33 b_2_32 0.108
R49_82 b_2_34 b_2_33 0.108
R49_83 b_2_35 b_2_34 0.108
R49_84 b_2_36 b_2_35 0.108
R49_85 b_2_37 b_2_36 0.108
R49_86 b_2_38 b_2_37 0.108
R49_87 b_2_39 b_2_38 0.108
R49_88 b_2_40 b_2_39 0.108
R49_89 b_2_41 b_2_40 0.001
R49_90 b_2_43 b_2_42 0.001
R49_91 b_2_46 b_2_43 0.54
R49_92 b_2_46 b_2_44 0.001
R49_93 b_2_45 b_2_46 0.108
R49_94 b_2_47 b_2_46 0.54
R49_95 b_2_48 b_2_47 0.108
R49_96 b_2_49 b_2_48 0.108
R49_97 b_2_50 b_2_49 0.108
R49_98 b_2_51 b_2_50 0.108
R49_99 b_2_52 b_2_51 0.108
R49_100 b_2_53 b_2_52 0.108
R49_101 b_2_54 b_2_53 0.108
R49_102 b_2_55 b_2_54 0.864
R49_103 b_2_56 b_2_55 0.108
R49_104 b_2_57 b_2_56 0.108
R49_105 b_2_58 b_2_57 0.108
R49_106 b_2_59 b_2_58 0.108
R49_107 b_2_60 b_2_59 0.108
R49_108 b_2_61 b_2_60 0.108
R49_109 b_2_62 b_2_61 0.108
R49_110 b_2_63 b_2_62 0.108
R49_111 b_2_64 b_2_63 0.108
R49_112 b_2_65 b_2_64 0.108
R49_113 b_2_66 b_2_65 0.108
R49_114 b_2_67 b_2_66 0.108
R49_115 b_2_68 b_2_67 0.108
R49_116 b_2_69 b_2_68 0.108
R49_117 b_2_70 b_2_69 0.108
R49_118 b_2_71 b_2_70 0.108
R49_119 b_2_72 b_2_71 0.108
R49_120 b_2_73 b_2_72 0.108
R49_121 b_2_74 b_2_73 0.108
R49_122 b_2_75 b_2_74 0.001
R49_123 b_2_76 b_2_75 0.216
R49_124 b_2_77 b_2_76 0.001
R49_125 b_2_78 b_2_77 0.001
R49_126 b_2_78 b_2_79 1.08
R49_127 b_2_80 b_2_79 2.268
R49_128 b_2_6 b_2_5 21.6
R49_129 b_2_83 b_2_80 0.324
R49_130 b_2_82 b_2_81 0.001
R49_131 b_2_83 b_2_82 0.216
R49_132 b_2_84 b_2_83 0.216
R49_133 b_2_85 b_2_84 0.001
R49_134 b_2_1 b_2_2 7.2
R49_135 b_2_3 b_2_2 7.2
R49_136 b_2_4 b_2_3 14.4

C2436 b_2 vss 4.3846e-15
C2437 b_2_42 vss 4.3846e-15
C2438 b_2_13 vss 1.40901e-16
C2439 b_2_45 vss 1.40901e-16
C2440 b_2_14 vss 3.13114e-17
C2441 b_2_13 vss 3.13114e-17
C2442 b_2_15 vss 3.13114e-17
C2443 b_2_14 vss 3.13114e-17
C2444 b_2_16 vss 3.13114e-17
C2445 b_2_15 vss 3.13114e-17
C2446 b_2_17 vss 3.13114e-17
C2447 b_2_16 vss 3.13114e-17
C2448 b_2_18 vss 3.13114e-17
C2449 b_2_17 vss 3.13114e-17
C2450 b_2_19 vss 3.13114e-17
C2451 b_2_18 vss 3.13114e-17
C2452 b_2_20 vss 3.13114e-17
C2453 b_2_19 vss 3.13114e-17
C2454 b_2_21 vss 2.42663e-16
C2455 b_2_20 vss 2.42663e-16
C2456 b_2_22 vss 3.13114e-17
C2457 b_2_21 vss 3.13114e-17
C2458 b_2_23 vss 3.13114e-17
C2459 b_2_22 vss 3.13114e-17
C2460 b_2_24 vss 3.13114e-17
C2461 b_2_23 vss 3.13114e-17
C2462 b_2_25 vss 3.13114e-17
C2463 b_2_24 vss 3.13114e-17
C2464 b_2_26 vss 3.13114e-17
C2465 b_2_25 vss 3.13114e-17
C2466 b_2_27 vss 3.13114e-17
C2467 b_2_26 vss 3.13114e-17
C2468 b_2_28 vss 3.13114e-17
C2469 b_2_27 vss 3.13114e-17
C2470 b_2_29 vss 3.13114e-17
C2471 b_2_28 vss 3.13114e-17
C2472 b_2_30 vss 3.13114e-17
C2473 b_2_29 vss 3.13114e-17
C2474 b_2_31 vss 3.13114e-17
C2475 b_2_30 vss 3.13114e-17
C2476 b_2_32 vss 3.13114e-17
C2477 b_2_31 vss 3.13114e-17
C2478 b_2_33 vss 3.13114e-17
C2479 b_2_32 vss 3.13114e-17
C2480 b_2_34 vss 3.13114e-17
C2481 b_2_33 vss 3.13114e-17
C2482 b_2_35 vss 3.13114e-17
C2483 b_2_34 vss 3.13114e-17
C2484 b_2_36 vss 3.13114e-17
C2485 b_2_35 vss 3.13114e-17
C2486 b_2_37 vss 3.13114e-17
C2487 b_2_36 vss 3.13114e-17
C2488 b_2_38 vss 3.13114e-17
C2489 b_2_37 vss 3.13114e-17
C2490 b_2_39 vss 3.13114e-17
C2491 b_2_38 vss 3.13114e-17
C2492 b_2_40 vss 3.13114e-17
C2493 b_2_39 vss 3.13114e-17
C2494 b_2_41 vss 1.40901e-17
C2495 b_2_40 vss 1.40901e-17
C2496 b_2_43 vss 3.48676e-17
C2497 b_2_42 vss 3.48676e-17
C2498 b_2_46 vss 6.8969e-16
C2499 b_2_43 vss 6.8969e-16
C2500 b_2_46 vss 6.34418e-17
C2501 b_2_44 vss 6.34418e-17
C2502 b_2_45 vss 1.42197e-16
C2503 b_2_46 vss 1.42197e-16
C2504 b_2_47 vss 1.40901e-16
C2505 b_2_46 vss 1.40901e-16
C2506 b_2_48 vss 3.13114e-17
C2507 b_2_47 vss 3.13114e-17
C2508 b_2_49 vss 3.13114e-17
C2509 b_2_48 vss 3.13114e-17
C2510 b_2_50 vss 3.13114e-17
C2511 b_2_49 vss 3.13114e-17
C2512 b_2_51 vss 3.13114e-17
C2513 b_2_50 vss 3.13114e-17
C2514 b_2_52 vss 3.13114e-17
C2515 b_2_51 vss 3.13114e-17
C2516 b_2_53 vss 3.13114e-17
C2517 b_2_52 vss 3.13114e-17
C2518 b_2_54 vss 3.13114e-17
C2519 b_2_53 vss 3.13114e-17
C2520 b_2_55 vss 2.42663e-16
C2521 b_2_54 vss 2.42663e-16
C2522 b_2_56 vss 3.13114e-17
C2523 b_2_55 vss 3.13114e-17
C2524 b_2_57 vss 3.13114e-17
C2525 b_2_56 vss 3.13114e-17
C2526 b_2_58 vss 3.13114e-17
C2527 b_2_57 vss 3.13114e-17
C2528 b_2_59 vss 3.13114e-17
C2529 b_2_58 vss 3.13114e-17
C2530 b_2_60 vss 3.13114e-17
C2531 b_2_59 vss 3.13114e-17
C2532 b_2_61 vss 3.13114e-17
C2533 b_2_60 vss 3.13114e-17
C2534 b_2_62 vss 3.13114e-17
C2535 b_2_61 vss 3.13114e-17
C2536 b_2_63 vss 3.13114e-17
C2537 b_2_62 vss 3.13114e-17
C2538 b_2_64 vss 3.13114e-17
C2539 b_2_63 vss 3.13114e-17
C2540 b_2_65 vss 3.13114e-17
C2541 b_2_64 vss 3.13114e-17
C2542 b_2_66 vss 3.13114e-17
C2543 b_2_65 vss 3.13114e-17
C2544 b_2_67 vss 3.13114e-17
C2545 b_2_66 vss 3.13114e-17
C2546 b_2_68 vss 3.13114e-17
C2547 b_2_67 vss 3.13114e-17
C2548 b_2_69 vss 3.13114e-17
C2549 b_2_68 vss 3.13114e-17
C2550 b_2_70 vss 3.13114e-17
C2551 b_2_69 vss 3.13114e-17
C2552 b_2_71 vss 3.13114e-17
C2553 b_2_70 vss 3.13114e-17
C2554 b_2_72 vss 3.13114e-17
C2555 b_2_71 vss 3.13114e-17
C2556 b_2_73 vss 3.13114e-17
C2557 b_2_72 vss 3.13114e-17
C2558 b_2_74 vss 3.13114e-17
C2559 b_2_73 vss 3.13114e-17
C2560 b_2_75 vss 1.40901e-17
C2561 b_2_74 vss 1.40901e-17
C2562 b_2_76 vss 8.14095e-17
C2563 b_2_75 vss 8.14095e-17
C2564 b_2_77 vss 1.25245e-17
C2565 b_2_76 vss 1.25245e-17
C2566 b_2_78 vss 2.50491e-17
C2567 b_2_77 vss 2.50491e-17
C2568 b_2_78 vss 2.97458e-16
C2569 b_2_79 vss 2.97458e-16
C2570 b_2_80 vss 6.18399e-16
C2571 b_2_79 vss 6.18399e-16
C2572 b_2_6 vss 9.46242e-17
C2573 b_2_5 vss 9.46242e-17
C2574 b_2_83 vss 9.39341e-17
C2575 b_2_80 vss 9.39341e-17
C2576 b_2_82 vss 1.40901e-17
C2577 b_2_81 vss 1.40901e-17
C2578 b_2_83 vss 7.04506e-17
C2579 b_2_82 vss 7.04506e-17
C2580 b_2_84 vss 7.82784e-17
C2581 b_2_83 vss 7.82784e-17
C2582 b_2_85 vss 1.40901e-17
C2583 b_2_84 vss 1.40901e-17
C2584 b_2_1 vss 3.15414e-17
C2585 b_2_2 vss 3.15414e-17
C2586 b_2_3 vss 3.15414e-17
C2587 b_2_2 vss 3.15414e-17
C2588 b_2_4 vss 6.30828e-17
C2589 b_2_3 vss 6.30828e-17

R50_1 n1496_39 n1496_7 0.001
R50_2 n1496_38 n1496_2 0.001
R50_3 n1496_1 n1496_18 0.001
R50_4 n1496_19 n1496_8 0.001
R50_5 n1496_36 n1496_7 0.001
R50_6 n1496_37 n1496_7 0.001
R50_7 n1496_16 n1496_8 0.001
R50_8 n1496_17 n1496_8 0.001
R50_9 n1496_4 n1496_30 0.001
R50_10 n1496_3 n1496_34 0.001
R50_11 n1496_35 n1496_7 0.001
R50_12 n1496_15 n1496_8 0.001
R50_13 n1496_20 n1496_10 0.001
R50_14 n1496_29 n1496_9 0.001
R50_15 n1496_28 n1496_13 0.001
R50_16 n1496_26 n1496_13 0.001
R50_17 n1496_27 n1496_13 0.001
R50_18 n1496_25 n1496_13 0.001
R50_19 n1496_24 n1496_13 0.001
R50_20 n1496_10 n1496_9 7.2
R50_21 n1496_11 n1496_10 21.6
R50_22 n1496_12 n1496_11 0.001
R50_23 n1496_15 n1496_14 0.001
R50_24 n1496_16 n1496_15 0.108
R50_25 n1496_17 n1496_16 0.108
R50_26 n1496_18 n1496_17 0.108
R50_27 n1496_19 n1496_18 0.108
R50_28 n1496_22 n1496_19 0.324
R50_29 n1496_2 n1496_1 0.216
R50_30 n1496_20 n1496_29 0.108
R50_31 n1496_21 n1496_20 0.001
R50_32 n1496_40 n1496_22 0.324
R50_33 n1496_24 n1496_23 0.001
R50_34 n1496_25 n1496_24 0.108
R50_35 n1496_26 n1496_25 0.108
R50_36 n1496_27 n1496_26 0.108
R50_37 n1496_28 n1496_27 0.108
R50_38 n1496_29 n1496_28 0.108
R50_39 n1496_32 n1496_29 0.216
R50_40 n1496_30 n1496_34 0.108
R50_41 n1496_31 n1496_30 0.001
R50_42 n1496_33 n1496_32 0.108
R50_43 n1496_34 n1496_33 0.216
R50_44 n1496_35 n1496_34 0.108
R50_45 n1496_36 n1496_35 0.108
R50_46 n1496_37 n1496_36 0.108
R50_47 n1496_38 n1496_37 0.108
R50_48 n1496_39 n1496_38 0.108
R50_49 n1496_40 n1496_39 0.324
R50_50 n1496_4 n1496_3 7.2
R50_51 n1496_5 n1496_4 21.6
R50_52 n1496 n1496_5 0.001

C2590 n1496_10 vss 4.20552e-17
C2591 n1496_9 vss 4.20552e-17
C2592 n1496_11 vss 9.46242e-17
C2593 n1496_10 vss 9.46242e-17
C2594 n1496_12 vss 5.47139e-16
C2595 n1496_11 vss 5.47139e-16
C2596 n1496_15 vss 1.40901e-17
C2597 n1496_14 vss 1.40901e-17
C2598 n1496_16 vss 3.91392e-17
C2599 n1496_15 vss 3.91392e-17
C2600 n1496_17 vss 3.91392e-17
C2601 n1496_16 vss 3.91392e-17
C2602 n1496_18 vss 3.91392e-17
C2603 n1496_17 vss 3.91392e-17
C2604 n1496_19 vss 3.91392e-17
C2605 n1496_18 vss 3.91392e-17
C2606 n1496_22 vss 1.0959e-16
C2607 n1496_19 vss 1.0959e-16
C2608 n1496_2 vss 7.81488e-17
C2609 n1496_1 vss 7.81488e-17
C2610 n1496_20 vss 3.71822e-17
C2611 n1496_29 vss 3.71822e-17
C2612 n1496_21 vss 1.40901e-17
C2613 n1496_20 vss 1.40901e-17
C2614 n1496_40 vss 9.39341e-17
C2615 n1496_22 vss 9.39341e-17
C2616 n1496_24 vss 1.40901e-17
C2617 n1496_23 vss 1.40901e-17
C2618 n1496_25 vss 3.91392e-17
C2619 n1496_24 vss 3.91392e-17
C2620 n1496_26 vss 3.91392e-17
C2621 n1496_25 vss 3.91392e-17
C2622 n1496_27 vss 4.6967e-17
C2623 n1496_26 vss 4.6967e-17
C2624 n1496_28 vss 3.91392e-17
C2625 n1496_27 vss 3.91392e-17
C2626 n1496_29 vss 4.6967e-17
C2627 n1496_28 vss 4.6967e-17
C2628 n1496_32 vss 6.41883e-17
C2629 n1496_29 vss 6.41883e-17
C2630 n1496_30 vss 3.71822e-17
C2631 n1496_34 vss 3.71822e-17
C2632 n1496_31 vss 1.40901e-17
C2633 n1496_30 vss 1.40901e-17
C2634 n1496_33 vss 2.81802e-17
C2635 n1496_32 vss 2.81802e-17
C2636 n1496_34 vss 5.63604e-17
C2637 n1496_33 vss 5.63604e-17
C2638 n1496_35 vss 4.6967e-17
C2639 n1496_34 vss 4.6967e-17
C2640 n1496_36 vss 3.91392e-17
C2641 n1496_35 vss 3.91392e-17
C2642 n1496_37 vss 3.91392e-17
C2643 n1496_36 vss 3.91392e-17
C2644 n1496_38 vss 3.91392e-17
C2645 n1496_37 vss 3.91392e-17
C2646 n1496_39 vss 3.91392e-17
C2647 n1496_38 vss 3.91392e-17
C2648 n1496_40 vss 1.0959e-16
C2649 n1496_39 vss 1.0959e-16
C2650 n1496_4 vss 4.20552e-17
C2651 n1496_3 vss 4.20552e-17
C2652 n1496_5 vss 9.46242e-17
C2653 n1496_4 vss 9.46242e-17
C2654 n1496 vss 3.05111e-16
C2655 n1496_5 vss 3.05111e-16

R51_1 b_1_2 b_1_84 0.001
R51_2 b_1_82 b_1_5 0.001
R51_3 b_1_42 b_1_7 0.001
R51_4 b_1_74 b_1_8 0.001
R51_5 b_1_40 b_1_7 0.001
R51_6 b_1_41 b_1_7 0.001
R51_7 b_1_72 b_1_8 0.001
R51_8 b_1_73 b_1_8 0.001
R51_9 b_1_38 b_1_7 0.001
R51_10 b_1_39 b_1_7 0.001
R51_11 b_1_71 b_1_8 0.001
R51_12 b_1_70 b_1_8 0.001
R51_13 b_1_37 b_1_7 0.001
R51_14 b_1_36 b_1_7 0.001
R51_15 b_1_68 b_1_8 0.001
R51_16 b_1_69 b_1_8 0.001
R51_17 b_1_34 b_1_7 0.001
R51_18 b_1_35 b_1_7 0.001
R51_19 b_1_67 b_1_8 0.001
R51_20 b_1_66 b_1_8 0.001
R51_21 b_1_32 b_1_7 0.001
R51_22 b_1_33 b_1_7 0.001
R51_23 b_1_64 b_1_8 0.001
R51_24 b_1_65 b_1_8 0.001
R51_25 b_1_30 b_1_7 0.001
R51_26 b_1_31 b_1_7 0.001
R51_27 b_1_63 b_1_8 0.001
R51_28 b_1_62 b_1_8 0.001
R51_29 b_1_29 b_1_7 0.001
R51_30 b_1_28 b_1_7 0.001
R51_31 b_1_60 b_1_8 0.001
R51_32 b_1_61 b_1_8 0.001
R51_33 b_1_27 b_1_7 0.001
R51_34 b_1_26 b_1_7 0.001
R51_35 b_1_59 b_1_8 0.001
R51_36 b_1_58 b_1_8 0.001
R51_37 b_1_24 b_1_7 0.001
R51_38 b_1_25 b_1_7 0.001
R51_39 b_1_56 b_1_8 0.001
R51_40 b_1_57 b_1_8 0.001
R51_41 b_1_23 b_1_7 0.001
R51_42 b_1_55 b_1_8 0.001
R51_43 b_1_22 b_1_9 0.001
R51_44 b_1_54 b_1_10 0.001
R51_45 b_1_21 b_1_9 0.001
R51_46 b_1_20 b_1_9 0.001
R51_47 b_1_53 b_1_10 0.001
R51_48 b_1_52 b_1_10 0.001
R51_49 b_1_18 b_1_9 0.001
R51_50 b_1_19 b_1_9 0.001
R51_51 b_1_51 b_1_10 0.001
R51_52 b_1_50 b_1_10 0.001
R51_53 b_1_16 b_1_9 0.001
R51_54 b_1_17 b_1_9 0.001
R51_55 b_1_48 b_1_10 0.001
R51_56 b_1_49 b_1_10 0.001
R51_57 b_1_15 b_1_9 0.001
R51_58 b_1_47 b_1_10 0.001
R51_59 b_1 b_1_11 0.001
R51_60 b_1 b_1_13 0.001
R51_61 b_1_14 b_1_13 0.001
R51_62 b_1_46 b_1_14 0.54
R51_63 b_1_15 b_1_45 0.54
R51_64 b_1_16 b_1_15 0.108
R51_65 b_1_17 b_1_16 0.108
R51_66 b_1_18 b_1_17 0.108
R51_67 b_1_19 b_1_18 0.108
R51_68 b_1_20 b_1_19 0.108
R51_69 b_1_21 b_1_20 0.108
R51_70 b_1_22 b_1_21 0.108
R51_71 b_1_23 b_1_22 0.864
R51_72 b_1_24 b_1_23 0.108
R51_73 b_1_25 b_1_24 0.108
R51_74 b_1_26 b_1_25 0.108
R51_75 b_1_27 b_1_26 0.108
R51_76 b_1_28 b_1_27 0.108
R51_77 b_1_29 b_1_28 0.108
R51_78 b_1_30 b_1_29 0.108
R51_79 b_1_31 b_1_30 0.108
R51_80 b_1_32 b_1_31 0.108
R51_81 b_1_33 b_1_32 0.108
R51_82 b_1_34 b_1_33 0.108
R51_83 b_1_35 b_1_34 0.108
R51_84 b_1_36 b_1_35 0.108
R51_85 b_1_37 b_1_36 0.108
R51_86 b_1_38 b_1_37 0.108
R51_87 b_1_39 b_1_38 0.108
R51_88 b_1_40 b_1_39 0.108
R51_89 b_1_41 b_1_40 0.108
R51_90 b_1_42 b_1_41 0.108
R51_91 b_1_43 b_1_42 0.001
R51_92 b_1_46 b_1_44 0.001
R51_93 b_1_45 b_1_46 0.108
R51_94 b_1_47 b_1_46 0.54
R51_95 b_1_48 b_1_47 0.108
R51_96 b_1_49 b_1_48 0.108
R51_97 b_1_50 b_1_49 0.108
R51_98 b_1_51 b_1_50 0.108
R51_99 b_1_52 b_1_51 0.108
R51_100 b_1_53 b_1_52 0.108
R51_101 b_1_54 b_1_53 0.108
R51_102 b_1_55 b_1_54 0.864
R51_103 b_1_56 b_1_55 0.108
R51_104 b_1_57 b_1_56 0.108
R51_105 b_1_58 b_1_57 0.108
R51_106 b_1_59 b_1_58 0.108
R51_107 b_1_60 b_1_59 0.108
R51_108 b_1_61 b_1_60 0.108
R51_109 b_1_62 b_1_61 0.108
R51_110 b_1_63 b_1_62 0.108
R51_111 b_1_64 b_1_63 0.108
R51_112 b_1_65 b_1_64 0.108
R51_113 b_1_66 b_1_65 0.108
R51_114 b_1_67 b_1_66 0.108
R51_115 b_1_68 b_1_67 0.108
R51_116 b_1_69 b_1_68 0.108
R51_117 b_1_70 b_1_69 0.108
R51_118 b_1_71 b_1_70 0.108
R51_119 b_1_72 b_1_71 0.108
R51_120 b_1_73 b_1_72 0.108
R51_121 b_1_74 b_1_73 0.108
R51_122 b_1_75 b_1_74 0.001
R51_123 b_1_76 b_1_75 0.216
R51_124 b_1_77 b_1_76 0.001
R51_125 b_1_78 b_1_77 0.001
R51_126 b_1_78 b_1_79 1.08
R51_127 b_1_80 b_1_79 2.268
R51_128 b_1_6 b_1_5 21.6
R51_129 b_1_83 b_1_80 0.324
R51_130 b_1_82 b_1_81 0.001
R51_131 b_1_83 b_1_82 0.216
R51_132 b_1_84 b_1_83 0.216
R51_133 b_1_85 b_1_84 0.001
R51_134 b_1_1 b_1_2 7.2
R51_135 b_1_3 b_1_2 7.2
R51_136 b_1_4 b_1_3 14.4

C2656 b_1 vss 4.3846e-15
C2657 b_1_13 vss 4.3846e-15
C2658 b_1_14 vss 3.48676e-17
C2659 b_1_13 vss 3.48676e-17
C2660 b_1_46 vss 6.8969e-16
C2661 b_1_14 vss 6.8969e-16
C2662 b_1_15 vss 1.40901e-16
C2663 b_1_45 vss 1.40901e-16
C2664 b_1_16 vss 3.13114e-17
C2665 b_1_15 vss 3.13114e-17
C2666 b_1_17 vss 3.13114e-17
C2667 b_1_16 vss 3.13114e-17
C2668 b_1_18 vss 3.13114e-17
C2669 b_1_17 vss 3.13114e-17
C2670 b_1_19 vss 3.13114e-17
C2671 b_1_18 vss 3.13114e-17
C2672 b_1_20 vss 3.13114e-17
C2673 b_1_19 vss 3.13114e-17
C2674 b_1_21 vss 3.13114e-17
C2675 b_1_20 vss 3.13114e-17
C2676 b_1_22 vss 3.13114e-17
C2677 b_1_21 vss 3.13114e-17
C2678 b_1_23 vss 2.42663e-16
C2679 b_1_22 vss 2.42663e-16
C2680 b_1_24 vss 3.13114e-17
C2681 b_1_23 vss 3.13114e-17
C2682 b_1_25 vss 3.13114e-17
C2683 b_1_24 vss 3.13114e-17
C2684 b_1_26 vss 3.13114e-17
C2685 b_1_25 vss 3.13114e-17
C2686 b_1_27 vss 3.13114e-17
C2687 b_1_26 vss 3.13114e-17
C2688 b_1_28 vss 3.13114e-17
C2689 b_1_27 vss 3.13114e-17
C2690 b_1_29 vss 3.13114e-17
C2691 b_1_28 vss 3.13114e-17
C2692 b_1_30 vss 3.13114e-17
C2693 b_1_29 vss 3.13114e-17
C2694 b_1_31 vss 3.13114e-17
C2695 b_1_30 vss 3.13114e-17
C2696 b_1_32 vss 3.13114e-17
C2697 b_1_31 vss 3.13114e-17
C2698 b_1_33 vss 3.13114e-17
C2699 b_1_32 vss 3.13114e-17
C2700 b_1_34 vss 3.13114e-17
C2701 b_1_33 vss 3.13114e-17
C2702 b_1_35 vss 3.13114e-17
C2703 b_1_34 vss 3.13114e-17
C2704 b_1_36 vss 3.13114e-17
C2705 b_1_35 vss 3.13114e-17
C2706 b_1_37 vss 3.13114e-17
C2707 b_1_36 vss 3.13114e-17
C2708 b_1_38 vss 3.13114e-17
C2709 b_1_37 vss 3.13114e-17
C2710 b_1_39 vss 3.13114e-17
C2711 b_1_38 vss 3.13114e-17
C2712 b_1_40 vss 3.13114e-17
C2713 b_1_39 vss 3.13114e-17
C2714 b_1_41 vss 3.13114e-17
C2715 b_1_40 vss 3.13114e-17
C2716 b_1_42 vss 3.13114e-17
C2717 b_1_41 vss 3.13114e-17
C2718 b_1_43 vss 1.40901e-17
C2719 b_1_42 vss 1.40901e-17
C2720 b_1_46 vss 6.34418e-17
C2721 b_1_44 vss 6.34418e-17
C2722 b_1_45 vss 1.42197e-16
C2723 b_1_46 vss 1.42197e-16
C2724 b_1_47 vss 1.40901e-16
C2725 b_1_46 vss 1.40901e-16
C2726 b_1_48 vss 3.13114e-17
C2727 b_1_47 vss 3.13114e-17
C2728 b_1_49 vss 3.13114e-17
C2729 b_1_48 vss 3.13114e-17
C2730 b_1_50 vss 3.13114e-17
C2731 b_1_49 vss 3.13114e-17
C2732 b_1_51 vss 3.13114e-17
C2733 b_1_50 vss 3.13114e-17
C2734 b_1_52 vss 3.13114e-17
C2735 b_1_51 vss 3.13114e-17
C2736 b_1_53 vss 3.13114e-17
C2737 b_1_52 vss 3.13114e-17
C2738 b_1_54 vss 3.13114e-17
C2739 b_1_53 vss 3.13114e-17
C2740 b_1_55 vss 2.42663e-16
C2741 b_1_54 vss 2.42663e-16
C2742 b_1_56 vss 3.13114e-17
C2743 b_1_55 vss 3.13114e-17
C2744 b_1_57 vss 3.13114e-17
C2745 b_1_56 vss 3.13114e-17
C2746 b_1_58 vss 3.13114e-17
C2747 b_1_57 vss 3.13114e-17
C2748 b_1_59 vss 3.13114e-17
C2749 b_1_58 vss 3.13114e-17
C2750 b_1_60 vss 3.13114e-17
C2751 b_1_59 vss 3.13114e-17
C2752 b_1_61 vss 3.13114e-17
C2753 b_1_60 vss 3.13114e-17
C2754 b_1_62 vss 3.13114e-17
C2755 b_1_61 vss 3.13114e-17
C2756 b_1_63 vss 3.13114e-17
C2757 b_1_62 vss 3.13114e-17
C2758 b_1_64 vss 3.13114e-17
C2759 b_1_63 vss 3.13114e-17
C2760 b_1_65 vss 3.13114e-17
C2761 b_1_64 vss 3.13114e-17
C2762 b_1_66 vss 3.13114e-17
C2763 b_1_65 vss 3.13114e-17
C2764 b_1_67 vss 3.13114e-17
C2765 b_1_66 vss 3.13114e-17
C2766 b_1_68 vss 3.13114e-17
C2767 b_1_67 vss 3.13114e-17
C2768 b_1_69 vss 3.13114e-17
C2769 b_1_68 vss 3.13114e-17
C2770 b_1_70 vss 3.13114e-17
C2771 b_1_69 vss 3.13114e-17
C2772 b_1_71 vss 3.13114e-17
C2773 b_1_70 vss 3.13114e-17
C2774 b_1_72 vss 3.13114e-17
C2775 b_1_71 vss 3.13114e-17
C2776 b_1_73 vss 3.13114e-17
C2777 b_1_72 vss 3.13114e-17
C2778 b_1_74 vss 3.13114e-17
C2779 b_1_73 vss 3.13114e-17
C2780 b_1_75 vss 1.40901e-17
C2781 b_1_74 vss 1.40901e-17
C2782 b_1_76 vss 8.14095e-17
C2783 b_1_75 vss 8.14095e-17
C2784 b_1_77 vss 1.25245e-17
C2785 b_1_76 vss 1.25245e-17
C2786 b_1_78 vss 2.50491e-17
C2787 b_1_77 vss 2.50491e-17
C2788 b_1_78 vss 2.97458e-16
C2789 b_1_79 vss 2.97458e-16
C2790 b_1_80 vss 6.18399e-16
C2791 b_1_79 vss 6.18399e-16
C2792 b_1_6 vss 9.46242e-17
C2793 b_1_5 vss 9.46242e-17
C2794 b_1_83 vss 9.39341e-17
C2795 b_1_80 vss 9.39341e-17
C2796 b_1_82 vss 1.40901e-17
C2797 b_1_81 vss 1.40901e-17
C2798 b_1_83 vss 7.04506e-17
C2799 b_1_82 vss 7.04506e-17
C2800 b_1_84 vss 7.82784e-17
C2801 b_1_83 vss 7.82784e-17
C2802 b_1_85 vss 1.40901e-17
C2803 b_1_84 vss 1.40901e-17
C2804 b_1_1 vss 3.15414e-17
C2805 b_1_2 vss 3.15414e-17
C2806 b_1_3 vss 3.15414e-17
C2807 b_1_2 vss 3.15414e-17
C2808 b_1_4 vss 6.30828e-17
C2809 b_1_3 vss 6.30828e-17

R52_1 n1625_7 n1625_39 0.001
R52_2 n1625_38 n1625_2 0.001
R52_3 n1625_1 n1625_18 0.001
R52_4 n1625_19 n1625_8 0.001
R52_5 n1625_7 n1625_36 0.001
R52_6 n1625_7 n1625_37 0.001
R52_7 n1625_16 n1625_8 0.001
R52_8 n1625_17 n1625_8 0.001
R52_9 n1625_30 n1625_4 0.001
R52_10 n1625_34 n1625_3 0.001
R52_11 n1625_7 n1625_35 0.001
R52_12 n1625_15 n1625_8 0.001
R52_13 n1625_20 n1625_10 0.001
R52_14 n1625_29 n1625_9 0.001
R52_15 n1625_28 n1625_13 0.001
R52_16 n1625_27 n1625_13 0.001
R52_17 n1625_26 n1625_13 0.001
R52_18 n1625_24 n1625_13 0.001
R52_19 n1625_25 n1625_13 0.001
R52_20 n1625_10 n1625_9 7.2
R52_21 n1625_11 n1625_10 21.6
R52_22 n1625_12 n1625_11 0.001
R52_23 n1625_15 n1625_14 0.001
R52_24 n1625_16 n1625_15 0.108
R52_25 n1625_17 n1625_16 0.108
R52_26 n1625_18 n1625_17 0.108
R52_27 n1625_19 n1625_18 0.108
R52_28 n1625_22 n1625_19 0.324
R52_29 n1625_2 n1625_1 0.216
R52_30 n1625_4 n1625_3 7.2
R52_31 n1625_5 n1625_4 21.6
R52_32 n1625 n1625_5 0.001
R52_33 n1625_20 n1625_29 0.108
R52_34 n1625_21 n1625_20 0.001
R52_35 n1625_40 n1625_22 0.324
R52_36 n1625_24 n1625_23 0.001
R52_37 n1625_25 n1625_24 0.108
R52_38 n1625_26 n1625_25 0.108
R52_39 n1625_27 n1625_26 0.108
R52_40 n1625_28 n1625_27 0.108
R52_41 n1625_29 n1625_28 0.108
R52_42 n1625_32 n1625_29 0.216
R52_43 n1625_30 n1625_34 0.108
R52_44 n1625_31 n1625_30 0.001
R52_45 n1625_33 n1625_32 0.108
R52_46 n1625_34 n1625_33 0.216
R52_47 n1625_35 n1625_34 0.108
R52_48 n1625_36 n1625_35 0.108
R52_49 n1625_37 n1625_36 0.108
R52_50 n1625_38 n1625_37 0.108
R52_51 n1625_39 n1625_38 0.108
R52_52 n1625_40 n1625_39 0.324

C2810 n1625_10 vss 4.20552e-17
C2811 n1625_9 vss 4.20552e-17
C2812 n1625_11 vss 9.46242e-17
C2813 n1625_10 vss 9.46242e-17
C2814 n1625_12 vss 5.47139e-16
C2815 n1625_11 vss 5.47139e-16
C2816 n1625_15 vss 1.40901e-17
C2817 n1625_14 vss 1.40901e-17
C2818 n1625_16 vss 3.91392e-17
C2819 n1625_15 vss 3.91392e-17
C2820 n1625_17 vss 3.91392e-17
C2821 n1625_16 vss 3.91392e-17
C2822 n1625_18 vss 3.91392e-17
C2823 n1625_17 vss 3.91392e-17
C2824 n1625_19 vss 3.91392e-17
C2825 n1625_18 vss 3.91392e-17
C2826 n1625_22 vss 1.0959e-16
C2827 n1625_19 vss 1.0959e-16
C2828 n1625_2 vss 7.81488e-17
C2829 n1625_1 vss 7.81488e-17
C2830 n1625_4 vss 4.20552e-17
C2831 n1625_3 vss 4.20552e-17
C2832 n1625_5 vss 9.46242e-17
C2833 n1625_4 vss 9.46242e-17
C2834 n1625 vss 3.05111e-16
C2835 n1625_5 vss 3.05111e-16
C2836 n1625_20 vss 3.71822e-17
C2837 n1625_29 vss 3.71822e-17
C2838 n1625_21 vss 1.40901e-17
C2839 n1625_20 vss 1.40901e-17
C2840 n1625_40 vss 9.39341e-17
C2841 n1625_22 vss 9.39341e-17
C2842 n1625_24 vss 1.40901e-17
C2843 n1625_23 vss 1.40901e-17
C2844 n1625_25 vss 3.91392e-17
C2845 n1625_24 vss 3.91392e-17
C2846 n1625_26 vss 3.91392e-17
C2847 n1625_25 vss 3.91392e-17
C2848 n1625_27 vss 4.6967e-17
C2849 n1625_26 vss 4.6967e-17
C2850 n1625_28 vss 3.91392e-17
C2851 n1625_27 vss 3.91392e-17
C2852 n1625_29 vss 4.6967e-17
C2853 n1625_28 vss 4.6967e-17
C2854 n1625_32 vss 6.41883e-17
C2855 n1625_29 vss 6.41883e-17
C2856 n1625_30 vss 3.71822e-17
C2857 n1625_34 vss 3.71822e-17
C2858 n1625_31 vss 1.40901e-17
C2859 n1625_30 vss 1.40901e-17
C2860 n1625_33 vss 2.81802e-17
C2861 n1625_32 vss 2.81802e-17
C2862 n1625_34 vss 5.63604e-17
C2863 n1625_33 vss 5.63604e-17
C2864 n1625_35 vss 4.6967e-17
C2865 n1625_34 vss 4.6967e-17
C2866 n1625_36 vss 3.91392e-17
C2867 n1625_35 vss 3.91392e-17
C2868 n1625_37 vss 3.91392e-17
C2869 n1625_36 vss 3.91392e-17
C2870 n1625_38 vss 3.91392e-17
C2871 n1625_37 vss 3.91392e-17
C2872 n1625_39 vss 3.91392e-17
C2873 n1625_38 vss 3.91392e-17
C2874 n1625_40 vss 1.0959e-16
C2875 n1625_39 vss 1.0959e-16

R53_1 n1644_2 n1644_33 0.001
R53_2 n1644_20 n1644_6 0.001
R53_3 n1644_1 n1644_32 0.001
R53_4 n1644_29 n1644_5 0.001
R53_5 n1644_39 n1644_9 0.001
R53_6 n1644_38 n1644_9 0.001
R53_7 n1644_36 n1644_9 0.001
R53_8 n1644_37 n1644_9 0.001
R53_9 n1644_35 n1644_9 0.001
R53_10 n1644_28 n1644_10 0.001
R53_11 n1644_26 n1644_10 0.001
R53_12 n1644_27 n1644_10 0.001
R53_13 n1644_24 n1644_10 0.001
R53_14 n1644_25 n1644_12 0.001
R53_15 n1644_17 n1644_13 0.001
R53_16 n1644_16 n1644_13 0.001
R53_17 n1644_18 n1644_13 0.001
R53_18 n1644_11 n1644_15 0.001
R53_19 n1644_14 n1644_13 0.001
R53_20 n1644_6 n1644_5 7.2
R53_21 n1644_7 n1644_6 21.6
R53_22 n1644 n1644_7 0.001
R53_23 n1644_14 n1644_22 0.324
R53_24 n1644_15 n1644_14 0.108
R53_25 n1644_16 n1644_15 0.108
R53_26 n1644_17 n1644_16 0.108
R53_27 n1644_18 n1644_17 0.108
R53_28 n1644_19 n1644_18 0.001
R53_29 n1644_12 n1644_11 0.216
R53_30 n1644_20 n1644_29 0.108
R53_31 n1644_21 n1644_20 0.001
R53_32 n1644_23 n1644_22 0.324
R53_33 n1644_24 n1644_23 0.324
R53_34 n1644_25 n1644_24 0.108
R53_35 n1644_26 n1644_25 0.108
R53_36 n1644_27 n1644_26 0.108
R53_37 n1644_28 n1644_27 0.108
R53_38 n1644_29 n1644_28 0.108
R53_39 n1644_30 n1644_29 0.216
R53_40 n1644_31 n1644_30 0.108
R53_41 n1644_32 n1644_31 0.216
R53_42 n1644_35 n1644_32 0.108
R53_43 n1644_36 n1644_35 0.108
R53_44 n1644_37 n1644_36 0.108
R53_45 n1644_38 n1644_37 0.108
R53_46 n1644_39 n1644_38 0.108
R53_47 n1644_40 n1644_39 0.001
R53_48 n1644_33 n1644_32 0.108
R53_49 n1644_34 n1644_33 0.001
R53_50 n1644_2 n1644_1 7.2
R53_51 n1644_3 n1644_2 21.6
R53_52 n1644_4 n1644_3 0.001

C2876 n1644_6 vss 4.20552e-17
C2877 n1644_5 vss 4.20552e-17
C2878 n1644_7 vss 9.46242e-17
C2879 n1644_6 vss 9.46242e-17
C2880 n1644 vss 3.05111e-16
C2881 n1644_7 vss 3.05111e-16
C2882 n1644_14 vss 1.0959e-16
C2883 n1644_22 vss 1.0959e-16
C2884 n1644_15 vss 3.91392e-17
C2885 n1644_14 vss 3.91392e-17
C2886 n1644_16 vss 3.91392e-17
C2887 n1644_15 vss 3.91392e-17
C2888 n1644_17 vss 3.91392e-17
C2889 n1644_16 vss 3.91392e-17
C2890 n1644_18 vss 3.91392e-17
C2891 n1644_17 vss 3.91392e-17
C2892 n1644_19 vss 1.40901e-17
C2893 n1644_18 vss 1.40901e-17
C2894 n1644_12 vss 7.81488e-17
C2895 n1644_11 vss 7.81488e-17
C2896 n1644_20 vss 3.71822e-17
C2897 n1644_29 vss 3.71822e-17
C2898 n1644_21 vss 1.40901e-17
C2899 n1644_20 vss 1.40901e-17
C2900 n1644_23 vss 9.39341e-17
C2901 n1644_22 vss 9.39341e-17
C2902 n1644_24 vss 1.0959e-16
C2903 n1644_23 vss 1.0959e-16
C2904 n1644_25 vss 3.91392e-17
C2905 n1644_24 vss 3.91392e-17
C2906 n1644_26 vss 3.91392e-17
C2907 n1644_25 vss 3.91392e-17
C2908 n1644_27 vss 3.91392e-17
C2909 n1644_26 vss 3.91392e-17
C2910 n1644_28 vss 3.91392e-17
C2911 n1644_27 vss 3.91392e-17
C2912 n1644_29 vss 4.6967e-17
C2913 n1644_28 vss 4.6967e-17
C2914 n1644_30 vss 5.63604e-17
C2915 n1644_29 vss 5.63604e-17
C2916 n1644_31 vss 2.81802e-17
C2917 n1644_30 vss 2.81802e-17
C2918 n1644_32 vss 6.41883e-17
C2919 n1644_31 vss 6.41883e-17
C2920 n1644_35 vss 4.6967e-17
C2921 n1644_32 vss 4.6967e-17
C2922 n1644_36 vss 3.91392e-17
C2923 n1644_35 vss 3.91392e-17
C2924 n1644_37 vss 4.6967e-17
C2925 n1644_36 vss 4.6967e-17
C2926 n1644_38 vss 3.91392e-17
C2927 n1644_37 vss 3.91392e-17
C2928 n1644_39 vss 3.91392e-17
C2929 n1644_38 vss 3.91392e-17
C2930 n1644_40 vss 1.40901e-17
C2931 n1644_39 vss 1.40901e-17
C2932 n1644_33 vss 3.71822e-17
C2933 n1644_32 vss 3.71822e-17
C2934 n1644_34 vss 1.40901e-17
C2935 n1644_33 vss 1.40901e-17
C2936 n1644_2 vss 4.20552e-17
C2937 n1644_1 vss 4.20552e-17
C2938 n1644_3 vss 9.46242e-17
C2939 n1644_2 vss 9.46242e-17
C2940 n1644_4 vss 5.47139e-16
C2941 n1644_3 vss 5.47139e-16

R1_1 b_0_50 b_0_1 0.001
R1_2 b_0_48 b_0_1 0.001
R1_3 b_0_49 b_0_1 0.001
R1_4 b_0_47 b_0_1 0.001
R1_5 b_0_46 b_0_1 0.001
R1_6 b_0_45 b_0_1 0.001
R1_7 b_0_44 b_0_1 0.001
R1_8 b_0_43 b_0_1 0.001
R1_9 b_0_42 b_0_2 0.001
R1_10 b_0_41 b_0_2 0.001
R1_11 b_0_39 b_0_2 0.001
R1_12 b_0_40 b_0_2 0.001
R1_13 b_0_38 b_0_2 0.001
R1_14 b_0_37 b_0_2 0.001
R1_15 b_0_36 b_0_2 0.001
R1_16 b_0_35 b_0_2 0.001
R1_17 b_0_34 b_0_2 0.001
R1_18 b_0_33 b_0_2 0.001
R1_19 b_0_32 b_0_2 0.001
R1_20 b_0_30 b_0_2 0.001
R1_21 b_0_31 b_0_2 0.001
R1_22 b_0_29 b_0_2 0.001
R1_23 b_0_28 b_0_2 0.001
R1_24 b_0_27 b_0_2 0.001
R1_25 b_0_26 b_0_2 0.001
R1_26 b_0_25 b_0_2 0.001
R1_27 b_0_24 b_0_2 0.001
R1_28 b_0_23 b_0_2 0.001
R1_29 b_0_79 b_0_3 0.001
R1_30 b_0_77 b_0_3 0.001
R1_31 b_0_78 b_0_3 0.001
R1_32 b_0_76 b_0_3 0.001
R1_33 b_0_75 b_0_3 0.001
R1_34 b_0_73 b_0_3 0.001
R1_35 b_0_74 b_0_3 0.001
R1_36 b_0_72 b_0_3 0.001
R1_37 b_0_70 b_0_4 0.001
R1_38 b_0_71 b_0_4 0.001
R1_39 b_0_68 b_0_4 0.001
R1_40 b_0_69 b_0_4 0.001
R1_41 b_0_65 b_0_4 0.001
R1_42 b_0_67 b_0_4 0.001
R1_43 b_0_66 b_0_4 0.001
R1_44 b_0_64 b_0_4 0.001
R1_45 b_0_63 b_0_4 0.001
R1_46 b_0_61 b_0_4 0.001
R1_47 b_0_62 b_0_4 0.001
R1_48 b_0_59 b_0_4 0.001
R1_49 b_0_60 b_0_4 0.001
R1_50 b_0_58 b_0_4 0.001
R1_51 b_0_57 b_0_4 0.001
R1_52 b_0_55 b_0_4 0.001
R1_53 b_0_56 b_0_4 0.001
R1_54 b_0_53 b_0_4 0.001
R1_55 b_0_54 b_0_4 0.001
R1_56 b_0_52 b_0_4 0.001
R1_57 b_0_14 b_0_5 0.001
R1_58 b_0_13 b_0_8 0.001
R1_59 b_0 b_0_11 0.001
R1_60 b_0_6 b_0_5 21.6
R1_61 b_0_8 b_0_7 7.2
R1_62 b_0_9 b_0_8 7.2
R1_63 b_0_10 b_0_9 14.4
R1_64 b_0_13 b_0_12 0.001
R1_65 b_0_16 b_0_13 0.216
R1_66 b_0_14 b_0_16 0.216
R1_67 b_0_15 b_0_14 0.001
R1_68 b_0_16 b_0_17 0.324
R1_69 b_0_18 b_0_17 2.268
R1_70 b_0_19 b_0_18 1.08
R1_71 b_0_20 b_0_19 0.001
R1_72 b_0_21 b_0_20 0.001
R1_73 b_0_51 b_0_21 0.216
R1_74 b_0_23 b_0_22 0.001
R1_75 b_0_24 b_0_23 0.108
R1_76 b_0_25 b_0_24 0.108
R1_77 b_0_26 b_0_25 0.108
R1_78 b_0_27 b_0_26 0.108
R1_79 b_0_28 b_0_27 0.108
R1_80 b_0_29 b_0_28 0.108
R1_81 b_0_30 b_0_29 0.108
R1_82 b_0_31 b_0_30 0.108
R1_83 b_0_32 b_0_31 0.108
R1_84 b_0_33 b_0_32 0.108
R1_85 b_0_34 b_0_33 0.108
R1_86 b_0_35 b_0_34 0.108
R1_87 b_0_36 b_0_35 0.108
R1_88 b_0_37 b_0_36 0.108
R1_89 b_0_38 b_0_37 0.108
R1_90 b_0_39 b_0_38 0.108
R1_91 b_0_40 b_0_39 0.108
R1_92 b_0_41 b_0_40 0.108
R1_93 b_0_42 b_0_41 0.108
R1_94 b_0_43 b_0_42 0.864
R1_95 b_0_44 b_0_43 0.108
R1_96 b_0_45 b_0_44 0.108
R1_97 b_0_46 b_0_45 0.108
R1_98 b_0_47 b_0_46 0.108
R1_99 b_0_48 b_0_47 0.108
R1_100 b_0_49 b_0_48 0.108
R1_101 b_0_50 b_0_49 0.108
R1_102 b_0_81 b_0_50 0.54
R1_103 b_0_52 b_0_51 0.001
R1_104 b_0_53 b_0_52 0.108
R1_105 b_0_54 b_0_53 0.108
R1_106 b_0_55 b_0_54 0.108
R1_107 b_0_56 b_0_55 0.108
R1_108 b_0_57 b_0_56 0.108
R1_109 b_0_58 b_0_57 0.108
R1_110 b_0_59 b_0_58 0.108
R1_111 b_0_60 b_0_59 0.108
R1_112 b_0_61 b_0_60 0.108
R1_113 b_0_62 b_0_61 0.108
R1_114 b_0_63 b_0_62 0.108
R1_115 b_0_64 b_0_63 0.108
R1_116 b_0_65 b_0_64 0.108
R1_117 b_0_66 b_0_65 0.108
R1_118 b_0_67 b_0_66 0.108
R1_119 b_0_68 b_0_67 0.108
R1_120 b_0_69 b_0_68 0.108
R1_121 b_0_70 b_0_69 0.108
R1_122 b_0_71 b_0_70 0.108
R1_123 b_0_72 b_0_71 0.864
R1_124 b_0_73 b_0_72 0.108
R1_125 b_0_74 b_0_73 0.108
R1_126 b_0_75 b_0_74 0.108
R1_127 b_0_76 b_0_75 0.108
R1_128 b_0_77 b_0_76 0.108
R1_129 b_0_78 b_0_77 0.108
R1_130 b_0_79 b_0_78 0.108
R1_131 b_0_82 b_0_79 0.54
R1_132 b_0_82 b_0_80 0.001
R1_133 b_0_81 b_0_82 0.108
R1_134 b_0_83 b_0_82 0.54
R1_135 b_0_84 b_0_83 0.001
R1_136 b_0 b_0_84 0.001

C2942 b_0_6 vss 9.46242e-17
C2943 b_0_5 vss 9.46242e-17
C2944 b_0_8 vss 3.15414e-17
C2945 b_0_7 vss 3.15414e-17
C2946 b_0_9 vss 3.15414e-17
C2947 b_0_8 vss 3.15414e-17
C2948 b_0_10 vss 6.30828e-17
C2949 b_0_9 vss 6.30828e-17
C2950 b_0_13 vss 1.40901e-17
C2951 b_0_12 vss 1.40901e-17
C2952 b_0_16 vss 7.82784e-17
C2953 b_0_13 vss 7.82784e-17
C2954 b_0_14 vss 7.04506e-17
C2955 b_0_16 vss 7.04506e-17
C2956 b_0_15 vss 1.40901e-17
C2957 b_0_14 vss 1.40901e-17
C2958 b_0_16 vss 9.39341e-17
C2959 b_0_17 vss 9.39341e-17
C2960 b_0_18 vss 6.18399e-16
C2961 b_0_17 vss 6.18399e-16
C2962 b_0_19 vss 2.97458e-16
C2963 b_0_18 vss 2.97458e-16
C2964 b_0_20 vss 2.50491e-17
C2965 b_0_19 vss 2.50491e-17
C2966 b_0_21 vss 1.25245e-17
C2967 b_0_20 vss 1.25245e-17
C2968 b_0_51 vss 8.14095e-17
C2969 b_0_21 vss 8.14095e-17
C2970 b_0_23 vss 1.40901e-17
C2971 b_0_22 vss 1.40901e-17
C2972 b_0_24 vss 3.13114e-17
C2973 b_0_23 vss 3.13114e-17
C2974 b_0_25 vss 3.13114e-17
C2975 b_0_24 vss 3.13114e-17
C2976 b_0_26 vss 3.13114e-17
C2977 b_0_25 vss 3.13114e-17
C2978 b_0_27 vss 3.13114e-17
C2979 b_0_26 vss 3.13114e-17
C2980 b_0_28 vss 3.13114e-17
C2981 b_0_27 vss 3.13114e-17
C2982 b_0_29 vss 3.13114e-17
C2983 b_0_28 vss 3.13114e-17
C2984 b_0_30 vss 3.13114e-17
C2985 b_0_29 vss 3.13114e-17
C2986 b_0_31 vss 3.13114e-17
C2987 b_0_30 vss 3.13114e-17
C2988 b_0_32 vss 3.13114e-17
C2989 b_0_31 vss 3.13114e-17
C2990 b_0_33 vss 3.13114e-17
C2991 b_0_32 vss 3.13114e-17
C2992 b_0_34 vss 3.13114e-17
C2993 b_0_33 vss 3.13114e-17
C2994 b_0_35 vss 3.13114e-17
C2995 b_0_34 vss 3.13114e-17
C2996 b_0_36 vss 3.13114e-17
C2997 b_0_35 vss 3.13114e-17
C2998 b_0_37 vss 3.13114e-17
C2999 b_0_36 vss 3.13114e-17
C3000 b_0_38 vss 3.13114e-17
C3001 b_0_37 vss 3.13114e-17
C3002 b_0_39 vss 3.13114e-17
C3003 b_0_38 vss 3.13114e-17
C3004 b_0_40 vss 3.13114e-17
C3005 b_0_39 vss 3.13114e-17
C3006 b_0_41 vss 3.13114e-17
C3007 b_0_40 vss 3.13114e-17
C3008 b_0_42 vss 3.13114e-17
C3009 b_0_41 vss 3.13114e-17
C3010 b_0_43 vss 2.42663e-16
C3011 b_0_42 vss 2.42663e-16
C3012 b_0_44 vss 3.13114e-17
C3013 b_0_43 vss 3.13114e-17
C3014 b_0_45 vss 3.13114e-17
C3015 b_0_44 vss 3.13114e-17
C3016 b_0_46 vss 3.13114e-17
C3017 b_0_45 vss 3.13114e-17
C3018 b_0_47 vss 3.13114e-17
C3019 b_0_46 vss 3.13114e-17
C3020 b_0_48 vss 3.13114e-17
C3021 b_0_47 vss 3.13114e-17
C3022 b_0_49 vss 3.13114e-17
C3023 b_0_48 vss 3.13114e-17
C3024 b_0_50 vss 3.13114e-17
C3025 b_0_49 vss 3.13114e-17
C3026 b_0_81 vss 1.40901e-16
C3027 b_0_50 vss 1.40901e-16
C3028 b_0_52 vss 1.40901e-17
C3029 b_0_51 vss 1.40901e-17
C3030 b_0_53 vss 3.13114e-17
C3031 b_0_52 vss 3.13114e-17
C3032 b_0_54 vss 3.13114e-17
C3033 b_0_53 vss 3.13114e-17
C3034 b_0_55 vss 3.13114e-17
C3035 b_0_54 vss 3.13114e-17
C3036 b_0_56 vss 3.13114e-17
C3037 b_0_55 vss 3.13114e-17
C3038 b_0_57 vss 3.13114e-17
C3039 b_0_56 vss 3.13114e-17
C3040 b_0_58 vss 3.13114e-17
C3041 b_0_57 vss 3.13114e-17
C3042 b_0_59 vss 3.13114e-17
C3043 b_0_58 vss 3.13114e-17
C3044 b_0_60 vss 3.13114e-17
C3045 b_0_59 vss 3.13114e-17
C3046 b_0_61 vss 3.13114e-17
C3047 b_0_60 vss 3.13114e-17
C3048 b_0_62 vss 3.13114e-17
C3049 b_0_61 vss 3.13114e-17
C3050 b_0_63 vss 3.13114e-17
C3051 b_0_62 vss 3.13114e-17
C3052 b_0_64 vss 3.13114e-17
C3053 b_0_63 vss 3.13114e-17
C3054 b_0_65 vss 3.13114e-17
C3055 b_0_64 vss 3.13114e-17
C3056 b_0_66 vss 3.13114e-17
C3057 b_0_65 vss 3.13114e-17
C3058 b_0_67 vss 3.13114e-17
C3059 b_0_66 vss 3.13114e-17
C3060 b_0_68 vss 3.13114e-17
C3061 b_0_67 vss 3.13114e-17
C3062 b_0_69 vss 3.13114e-17
C3063 b_0_68 vss 3.13114e-17
C3064 b_0_70 vss 3.13114e-17
C3065 b_0_69 vss 3.13114e-17
C3066 b_0_71 vss 3.13114e-17
C3067 b_0_70 vss 3.13114e-17
C3068 b_0_72 vss 2.42663e-16
C3069 b_0_71 vss 2.42663e-16
C3070 b_0_73 vss 3.13114e-17
C3071 b_0_72 vss 3.13114e-17
C3072 b_0_74 vss 3.13114e-17
C3073 b_0_73 vss 3.13114e-17
C3074 b_0_75 vss 3.13114e-17
C3075 b_0_74 vss 3.13114e-17
C3076 b_0_76 vss 3.13114e-17
C3077 b_0_75 vss 3.13114e-17
C3078 b_0_77 vss 3.13114e-17
C3079 b_0_76 vss 3.13114e-17
C3080 b_0_78 vss 3.13114e-17
C3081 b_0_77 vss 3.13114e-17
C3082 b_0_79 vss 3.13114e-17
C3083 b_0_78 vss 3.13114e-17
C3084 b_0_82 vss 1.40901e-16
C3085 b_0_79 vss 1.40901e-16
C3086 b_0_82 vss 6.34418e-17
C3087 b_0_80 vss 6.34418e-17
C3088 b_0_81 vss 1.42197e-16
C3089 b_0_82 vss 1.42197e-16
C3090 b_0_83 vss 6.8969e-16
C3091 b_0_82 vss 6.8969e-16
C3092 b_0_84 vss 3.48676e-17
C3093 b_0_83 vss 3.48676e-17
C3094 b_0 vss 4.3846e-15
C3095 b_0_84 vss 4.3846e-15

R54_1 ck_101 ck_1 0.001
R54_2 ck_100 ck_1 0.001
R54_3 ck_99 ck_1 0.001
R54_4 ck_98 ck_1 0.001
R54_5 ck_97 ck_1 0.001
R54_6 ck_96 ck_1 0.001
R54_7 ck_95 ck_1 0.001
R54_8 ck_93 ck_1 0.001
R54_9 ck_94 ck_1 0.001
R54_10 ck_92 ck_1 0.001
R54_11 ck_91 ck_1 0.001
R54_12 ck_90 ck_1 0.001
R54_13 ck_89 ck_1 0.001
R54_14 ck_88 ck_1 0.001
R54_15 ck_87 ck_1 0.001
R54_16 ck_85 ck_1 0.001
R54_17 ck_86 ck_1 0.001
R54_18 ck_83 ck_1 0.001
R54_19 ck_84 ck_1 0.001
R54_20 ck_82 ck_1 0.001
R54_21 ck_81 ck_2 0.001
R54_22 ck_79 ck_2 0.001
R54_23 ck_80 ck_2 0.001
R54_24 ck_78 ck_2 0.001
R54_25 ck_77 ck_2 0.001
R54_26 ck_75 ck_2 0.001
R54_27 ck_76 ck_2 0.001
R54_28 ck_74 ck_2 0.001
R54_29 ck_66 ck_3 0.001
R54_30 ck_65 ck_3 0.001
R54_31 ck_64 ck_3 0.001
R54_32 ck_63 ck_3 0.001
R54_33 ck_62 ck_3 0.001
R54_34 ck_61 ck_3 0.001
R54_35 ck_60 ck_3 0.001
R54_36 ck_58 ck_3 0.001
R54_37 ck_59 ck_3 0.001
R54_38 ck_56 ck_3 0.001
R54_39 ck_57 ck_3 0.001
R54_40 ck_55 ck_3 0.001
R54_41 ck_54 ck_3 0.001
R54_42 ck_53 ck_3 0.001
R54_43 ck_52 ck_3 0.001
R54_44 ck_50 ck_3 0.001
R54_45 ck_51 ck_3 0.001
R54_46 ck_48 ck_3 0.001
R54_47 ck_49 ck_3 0.001
R54_48 ck_47 ck_3 0.001
R54_49 ck_46 ck_4 0.001
R54_50 ck_44 ck_4 0.001
R54_51 ck_45 ck_4 0.001
R54_52 ck_43 ck_4 0.001
R54_53 ck_42 ck_4 0.001
R54_54 ck_41 ck_4 0.001
R54_55 ck_40 ck_4 0.001
R54_56 ck_39 ck_4 0.001
R54_57 ck_29 ck_6 0.001
R54_58 ck_33 ck_5 0.001
R54_59 ck_35 ck_19 0.001
R54_60 ck_16 ck_28 0.001
R54_61 ck_13 ck_27 0.001
R54_62 ck ck_26 0.001
R54_63 ck_27 ck_31 0.324
R54_64 ck_28 ck_32 0.324
R54_65 ck_12 ck_11 14.4
R54_66 ck_13 ck_12 7.2
R54_67 ck_14 ck_13 7.2
R54_68 ck_15 ck_14 14.4
R54_69 ck_16 ck_15 7.2
R54_70 ck_17 ck_16 7.2
R54_71 ck_18 ck_17 14.4
R54_72 ck_19 ck_18 7.2
R54_73 ck_20 ck_19 7.2
R54_74 ck_21 ck_20 14.4
R54_75 ck_22 ck_21 14.4
R54_76 ck_23 ck_22 14.4
R54_77 ck_24 ck_23 14.4
R54_78 ck_25 ck_24 14.4
R54_79 ck_6 ck_5 7.2
R54_80 ck_7 ck_6 21.6
R54_81 ck_8 ck_7 14.4
R54_82 ck_9 ck_8 14.4
R54_83 ck_10 ck_9 14.4
R54_84 ck_29 ck_33 0.108
R54_85 ck_30 ck_29 0.001
R54_86 ck_32 ck_31 0.432
R54_87 ck_34 ck_32 0.432
R54_88 ck_33 ck_37 2.052
R54_89 ck_34 ck_33 0.216
R54_90 ck_35 ck_34 0.216
R54_91 ck_36 ck_35 0.001
R54_92 ck_38 ck_37 0.864
R54_93 ck_38 ck_67 0.432
R54_94 ck_39 ck_70 0.54
R54_95 ck_40 ck_39 0.108
R54_96 ck_41 ck_40 0.108
R54_97 ck_42 ck_41 0.108
R54_98 ck_43 ck_42 0.108
R54_99 ck_44 ck_43 0.108
R54_100 ck_45 ck_44 0.108
R54_101 ck_46 ck_45 0.108
R54_102 ck_47 ck_46 0.864
R54_103 ck_48 ck_47 0.108
R54_104 ck_49 ck_48 0.108
R54_105 ck_50 ck_49 0.108
R54_106 ck_51 ck_50 0.108
R54_107 ck_52 ck_51 0.108
R54_108 ck_53 ck_52 0.108
R54_109 ck_54 ck_53 0.108
R54_110 ck_55 ck_54 0.108
R54_111 ck_56 ck_55 0.108
R54_112 ck_57 ck_56 0.108
R54_113 ck_58 ck_57 0.108
R54_114 ck_59 ck_58 0.108
R54_115 ck_60 ck_59 0.108
R54_116 ck_61 ck_60 0.108
R54_117 ck_62 ck_61 0.108
R54_118 ck_63 ck_62 0.108
R54_119 ck_64 ck_63 0.108
R54_120 ck_65 ck_64 0.108
R54_121 ck_66 ck_65 0.108
R54_122 ck_67 ck_66 0.001
R54_123 ck_74 ck_69 0.54
R54_124 ck_75 ck_74 0.108
R54_125 ck_76 ck_75 0.108
R54_126 ck_77 ck_76 0.108
R54_127 ck_78 ck_77 0.108
R54_128 ck_79 ck_78 0.108
R54_129 ck_80 ck_79 0.108
R54_130 ck_81 ck_80 0.108
R54_131 ck_82 ck_81 0.864
R54_132 ck_83 ck_82 0.108
R54_133 ck_84 ck_83 0.108
R54_134 ck_85 ck_84 0.108
R54_135 ck_86 ck_85 0.108
R54_136 ck_87 ck_86 0.108
R54_137 ck_88 ck_87 0.108
R54_138 ck_89 ck_88 0.108
R54_139 ck_90 ck_89 0.108
R54_140 ck_91 ck_90 0.108
R54_141 ck_92 ck_91 0.108
R54_142 ck_93 ck_92 0.108
R54_143 ck_94 ck_93 0.108
R54_144 ck_95 ck_94 0.108
R54_145 ck_96 ck_95 0.108
R54_146 ck_97 ck_96 0.108
R54_147 ck_98 ck_97 0.108
R54_148 ck_99 ck_98 0.108
R54_149 ck_100 ck_99 0.108
R54_150 ck_101 ck_100 0.108
R54_151 ck_102 ck_101 0.001
R54_152 ck_70 ck_68 0.001
R54_153 ck_69 ck_70 0.108
R54_154 ck_70 ck_73 0.54
R54_155 ck ck_72 0.001
R54_156 ck_73 ck_72 0.001

C3096 ck_27 vss 6.5785e-17
C3097 ck_31 vss 6.5785e-17
C3098 ck_28 vss 6.5785e-17
C3099 ck_32 vss 6.5785e-17
C3100 ck_12 vss 6.30828e-17
C3101 ck_11 vss 6.30828e-17
C3102 ck_13 vss 3.15414e-17
C3103 ck_12 vss 3.15414e-17
C3104 ck_14 vss 3.15414e-17
C3105 ck_13 vss 3.15414e-17
C3106 ck_15 vss 6.30828e-17
C3107 ck_14 vss 6.30828e-17
C3108 ck_16 vss 3.15414e-17
C3109 ck_15 vss 3.15414e-17
C3110 ck_17 vss 3.15414e-17
C3111 ck_16 vss 3.15414e-17
C3112 ck_18 vss 6.30828e-17
C3113 ck_17 vss 6.30828e-17
C3114 ck_19 vss 3.15414e-17
C3115 ck_18 vss 3.15414e-17
C3116 ck_20 vss 3.15414e-17
C3117 ck_19 vss 3.15414e-17
C3118 ck_21 vss 6.30828e-17
C3119 ck_20 vss 6.30828e-17
C3120 ck_22 vss 6.30828e-17
C3121 ck_21 vss 6.30828e-17
C3122 ck_23 vss 6.30828e-17
C3123 ck_22 vss 6.30828e-17
C3124 ck_24 vss 6.30828e-17
C3125 ck_23 vss 6.30828e-17
C3126 ck_25 vss 6.30828e-17
C3127 ck_24 vss 6.30828e-17
C3128 ck_6 vss 4.20552e-17
C3129 ck_5 vss 4.20552e-17
C3130 ck_7 vss 9.46242e-17
C3131 ck_6 vss 9.46242e-17
C3132 ck_8 vss 6.30828e-17
C3133 ck_7 vss 6.30828e-17
C3134 ck_9 vss 6.30828e-17
C3135 ck_8 vss 6.30828e-17
C3136 ck_10 vss 6.30828e-17
C3137 ck_9 vss 6.30828e-17
C3138 ck_29 vss 4.10962e-17
C3139 ck_33 vss 4.10962e-17
C3140 ck_30 vss 1.40901e-17
C3141 ck_29 vss 1.40901e-17
C3142 ck_32 vss 8.77133e-17
C3143 ck_31 vss 8.77133e-17
C3144 ck_34 vss 8.77133e-17
C3145 ck_32 vss 8.77133e-17
C3146 ck_33 vss 5.47949e-16
C3147 ck_37 vss 5.47949e-16
C3148 ck_34 vss 7.82784e-17
C3149 ck_33 vss 7.82784e-17
C3150 ck_35 vss 7.04506e-17
C3151 ck_34 vss 7.04506e-17
C3152 ck_36 vss 1.40901e-17
C3153 ck_35 vss 1.40901e-17
C3154 ck_38 vss 2.50491e-16
C3155 ck_37 vss 2.50491e-16
C3156 ck_38 vss 1.18983e-16
C3157 ck_67 vss 1.18983e-16
C3158 ck_39 vss 1.40901e-16
C3159 ck_70 vss 1.40901e-16
C3160 ck_40 vss 3.13114e-17
C3161 ck_39 vss 3.13114e-17
C3162 ck_41 vss 3.13114e-17
C3163 ck_40 vss 3.13114e-17
C3164 ck_42 vss 3.13114e-17
C3165 ck_41 vss 3.13114e-17
C3166 ck_43 vss 3.13114e-17
C3167 ck_42 vss 3.13114e-17
C3168 ck_44 vss 3.13114e-17
C3169 ck_43 vss 3.13114e-17
C3170 ck_45 vss 3.13114e-17
C3171 ck_44 vss 3.13114e-17
C3172 ck_46 vss 3.13114e-17
C3173 ck_45 vss 3.13114e-17
C3174 ck_47 vss 2.42663e-16
C3175 ck_46 vss 2.42663e-16
C3176 ck_48 vss 3.13114e-17
C3177 ck_47 vss 3.13114e-17
C3178 ck_49 vss 3.13114e-17
C3179 ck_48 vss 3.13114e-17
C3180 ck_50 vss 3.13114e-17
C3181 ck_49 vss 3.13114e-17
C3182 ck_51 vss 3.13114e-17
C3183 ck_50 vss 3.13114e-17
C3184 ck_52 vss 3.13114e-17
C3185 ck_51 vss 3.13114e-17
C3186 ck_53 vss 3.13114e-17
C3187 ck_52 vss 3.13114e-17
C3188 ck_54 vss 3.13114e-17
C3189 ck_53 vss 3.13114e-17
C3190 ck_55 vss 3.13114e-17
C3191 ck_54 vss 3.13114e-17
C3192 ck_56 vss 3.13114e-17
C3193 ck_55 vss 3.13114e-17
C3194 ck_57 vss 3.13114e-17
C3195 ck_56 vss 3.13114e-17
C3196 ck_58 vss 3.13114e-17
C3197 ck_57 vss 3.13114e-17
C3198 ck_59 vss 3.13114e-17
C3199 ck_58 vss 3.13114e-17
C3200 ck_60 vss 3.13114e-17
C3201 ck_59 vss 3.13114e-17
C3202 ck_61 vss 3.13114e-17
C3203 ck_60 vss 3.13114e-17
C3204 ck_62 vss 3.13114e-17
C3205 ck_61 vss 3.13114e-17
C3206 ck_63 vss 3.13114e-17
C3207 ck_62 vss 3.13114e-17
C3208 ck_64 vss 3.13114e-17
C3209 ck_63 vss 3.13114e-17
C3210 ck_65 vss 3.13114e-17
C3211 ck_64 vss 3.13114e-17
C3212 ck_66 vss 3.13114e-17
C3213 ck_65 vss 3.13114e-17
C3214 ck_67 vss 1.40901e-17
C3215 ck_66 vss 1.40901e-17
C3216 ck_74 vss 1.40901e-16
C3217 ck_69 vss 1.40901e-16
C3218 ck_75 vss 3.13114e-17
C3219 ck_74 vss 3.13114e-17
C3220 ck_76 vss 3.13114e-17
C3221 ck_75 vss 3.13114e-17
C3222 ck_77 vss 3.13114e-17
C3223 ck_76 vss 3.13114e-17
C3224 ck_78 vss 3.13114e-17
C3225 ck_77 vss 3.13114e-17
C3226 ck_79 vss 3.13114e-17
C3227 ck_78 vss 3.13114e-17
C3228 ck_80 vss 3.13114e-17
C3229 ck_79 vss 3.13114e-17
C3230 ck_81 vss 3.13114e-17
C3231 ck_80 vss 3.13114e-17
C3232 ck_82 vss 2.42663e-16
C3233 ck_81 vss 2.42663e-16
C3234 ck_83 vss 3.13114e-17
C3235 ck_82 vss 3.13114e-17
C3236 ck_84 vss 3.13114e-17
C3237 ck_83 vss 3.13114e-17
C3238 ck_85 vss 3.13114e-17
C3239 ck_84 vss 3.13114e-17
C3240 ck_86 vss 3.13114e-17
C3241 ck_85 vss 3.13114e-17
C3242 ck_87 vss 3.13114e-17
C3243 ck_86 vss 3.13114e-17
C3244 ck_88 vss 3.13114e-17
C3245 ck_87 vss 3.13114e-17
C3246 ck_89 vss 3.13114e-17
C3247 ck_88 vss 3.13114e-17
C3248 ck_90 vss 3.13114e-17
C3249 ck_89 vss 3.13114e-17
C3250 ck_91 vss 3.13114e-17
C3251 ck_90 vss 3.13114e-17
C3252 ck_92 vss 3.13114e-17
C3253 ck_91 vss 3.13114e-17
C3254 ck_93 vss 3.13114e-17
C3255 ck_92 vss 3.13114e-17
C3256 ck_94 vss 3.13114e-17
C3257 ck_93 vss 3.13114e-17
C3258 ck_95 vss 3.13114e-17
C3259 ck_94 vss 3.13114e-17
C3260 ck_96 vss 3.13114e-17
C3261 ck_95 vss 3.13114e-17
C3262 ck_97 vss 3.13114e-17
C3263 ck_96 vss 3.13114e-17
C3264 ck_98 vss 3.13114e-17
C3265 ck_97 vss 3.13114e-17
C3266 ck_99 vss 3.13114e-17
C3267 ck_98 vss 3.13114e-17
C3268 ck_100 vss 3.13114e-17
C3269 ck_99 vss 3.13114e-17
C3270 ck_101 vss 3.13114e-17
C3271 ck_100 vss 3.13114e-17
C3272 ck_102 vss 1.40901e-17
C3273 ck_101 vss 1.40901e-17
C3274 ck_70 vss 6.34418e-17
C3275 ck_68 vss 6.34418e-17
C3276 ck_69 vss 1.42197e-16
C3277 ck_70 vss 1.42197e-16
C3278 ck_70 vss 6.8969e-16
C3279 ck_73 vss 6.8969e-16
C3280 ck vss 4.3846e-15
C3281 ck_72 vss 4.3846e-15
C3282 ck_73 vss 3.48676e-17
C3283 ck_72 vss 3.48676e-17

R55_1 n1874_101 n1874_1 0.001
R55_2 n1874_100 n1874_1 0.001
R55_3 n1874_99 n1874_1 0.001
R55_4 n1874_98 n1874_1 0.001
R55_5 n1874_97 n1874_1 0.001
R55_6 n1874_3 n1874_95 0.001
R55_7 n1874_2 n1874_94 0.001
R55_8 n1874_91 n1874_12 0.001
R55_9 n1874_77 n1874_13 0.001
R55_10 n1874_90 n1874_22 0.001
R55_11 n1874_89 n1874_22 0.001
R55_12 n1874_87 n1874_22 0.001
R55_13 n1874_88 n1874_22 0.001
R55_14 n1874_86 n1874_22 0.001
R55_15 n1874_41 n1874_23 0.001
R55_16 n1874_40 n1874_23 0.001
R55_17 n1874_39 n1874_23 0.001
R55_18 n1874_38 n1874_23 0.001
R55_19 n1874_37 n1874_23 0.001
R55_20 n1874_36 n1874_24 0.001
R55_21 n1874_35 n1874_24 0.001
R55_22 n1874_34 n1874_24 0.001
R55_23 n1874_33 n1874_24 0.001
R55_24 n1874_32 n1874_24 0.001
R55_25 n1874_58 n1874_25 0.001
R55_26 n1874_57 n1874_25 0.001
R55_27 n1874_56 n1874_25 0.001
R55_28 n1874_55 n1874_25 0.001
R55_29 n1874_54 n1874_25 0.001
R55_30 n1874_53 n1874_26 0.001
R55_31 n1874_52 n1874_26 0.001
R55_32 n1874_51 n1874_26 0.001
R55_33 n1874_50 n1874_26 0.001
R55_34 n1874_49 n1874_26 0.001
R55_35 n1874_47 n1874_27 0.001
R55_36 n1874_45 n1874_27 0.001
R55_37 n1874_46 n1874_27 0.001
R55_38 n1874_44 n1874_27 0.001
R55_39 n1874_43 n1874_27 0.001
R55_40 n1874_76 n1874_28 0.001
R55_41 n1874_75 n1874_28 0.001
R55_42 n1874_74 n1874_28 0.001
R55_43 n1874_73 n1874_28 0.001
R55_44 n1874_72 n1874_28 0.001
R55_45 n1874_64 n1874 0.001
R55_46 n1874_62 n1874 0.001
R55_47 n1874_63 n1874 0.001
R55_48 n1874_61 n1874 0.001
R55_49 n1874_60 n1874 0.001
R55_50 n1874_70 n1874_30 0.001
R55_51 n1874_68 n1874_30 0.001
R55_52 n1874_69 n1874_30 0.001
R55_53 n1874_67 n1874_30 0.001
R55_54 n1874_66 n1874_30 0.001
R55_55 n1874_13 n1874_12 7.2
R55_56 n1874_14 n1874_13 21.6
R55_57 n1874_15 n1874_14 0.001
R55_58 n1874_16 n1874_15 0.001
R55_59 n1874_17 n1874_16 0.001
R55_60 n1874_18 n1874_17 0.001
R55_61 n1874_19 n1874_18 0.001
R55_62 n1874_20 n1874_19 0.001
R55_63 n1874_21 n1874_20 0.001
R55_64 n1874_32 n1874_31 0.001
R55_65 n1874_33 n1874_32 0.108
R55_66 n1874_34 n1874_33 0.108
R55_67 n1874_35 n1874_34 0.108
R55_68 n1874_36 n1874_35 0.108
R55_69 n1874_37 n1874_36 0.864
R55_70 n1874_38 n1874_37 0.108
R55_71 n1874_39 n1874_38 0.108
R55_72 n1874_40 n1874_39 0.108
R55_73 n1874_41 n1874_40 0.108
R55_74 n1874_84 n1874_41 0.324
R55_75 n1874_43 n1874_42 0.001
R55_76 n1874_44 n1874_43 0.108
R55_77 n1874_45 n1874_44 0.108
R55_78 n1874_46 n1874_45 0.108
R55_79 n1874_47 n1874_46 0.108
R55_80 n1874_82 n1874_47 0.324
R55_81 n1874_49 n1874_48 0.001
R55_82 n1874_50 n1874_49 0.108
R55_83 n1874_51 n1874_50 0.108
R55_84 n1874_52 n1874_51 0.108
R55_85 n1874_53 n1874_52 0.108
R55_86 n1874_54 n1874_53 0.864
R55_87 n1874_55 n1874_54 0.108
R55_88 n1874_56 n1874_55 0.108
R55_89 n1874_57 n1874_56 0.108
R55_90 n1874_58 n1874_57 0.108
R55_91 n1874_83 n1874_58 0.324
R55_92 n1874_60 n1874_59 0.001
R55_93 n1874_61 n1874_60 0.108
R55_94 n1874_62 n1874_61 0.108
R55_95 n1874_63 n1874_62 0.108
R55_96 n1874_64 n1874_63 0.108
R55_97 n1874_80 n1874_64 0.324
R55_98 n1874_66 n1874_65 0.001
R55_99 n1874_67 n1874_66 0.108
R55_100 n1874_68 n1874_67 0.108
R55_101 n1874_69 n1874_68 0.108
R55_102 n1874_70 n1874_69 0.108
R55_103 n1874_79 n1874_70 0.324
R55_104 n1874_72 n1874_71 0.001
R55_105 n1874_73 n1874_72 0.108
R55_106 n1874_74 n1874_73 0.108
R55_107 n1874_75 n1874_74 0.108
R55_108 n1874_76 n1874_75 0.108
R55_109 n1874_81 n1874_76 0.324
R55_110 n1874_77 n1874_91 0.108
R55_111 n1874_78 n1874_77 0.001
R55_112 n1874_80 n1874_79 0.324
R55_113 n1874_81 n1874_80 0.324
R55_114 n1874_82 n1874_81 0.324
R55_115 n1874_83 n1874_82 0.324
R55_116 n1874_84 n1874_83 0.324
R55_117 n1874_102 n1874_84 0.324
R55_118 n1874_86 n1874_85 0.001
R55_119 n1874_87 n1874_86 0.108
R55_120 n1874_88 n1874_87 0.108
R55_121 n1874_89 n1874_88 0.108
R55_122 n1874_90 n1874_89 0.108
R55_123 n1874_91 n1874_90 0.108
R55_124 n1874_92 n1874_91 0.216
R55_125 n1874_93 n1874_92 0.108
R55_126 n1874_94 n1874_93 0.216
R55_127 n1874_97 n1874_94 0.108
R55_128 n1874_98 n1874_97 0.108
R55_129 n1874_99 n1874_98 0.108
R55_130 n1874_100 n1874_99 0.108
R55_131 n1874_101 n1874_100 0.108
R55_132 n1874_102 n1874_101 0.324
R55_133 n1874_95 n1874_94 0.108
R55_134 n1874_96 n1874_95 0.001
R55_135 n1874_3 n1874_2 7.2
R55_136 n1874_4 n1874_3 21.6
R55_137 n1874_5 n1874_4 0.001
R55_138 n1874_6 n1874_5 0.001
R55_139 n1874_7 n1874_6 0.001
R55_140 n1874_8 n1874_7 0.001
R55_141 n1874_9 n1874_8 0.001
R55_142 n1874_10 n1874_9 0.001
R55_143 n1874_11 n1874_10 0.001

C3284 n1874_13 vss 4.20552e-17
C3285 n1874_12 vss 4.20552e-17
C3286 n1874_14 vss 9.46242e-17
C3287 n1874_13 vss 9.46242e-17
C3288 n1874_15 vss 5.47139e-16
C3289 n1874_14 vss 5.47139e-16
C3290 n1874_16 vss 5.47139e-16
C3291 n1874_15 vss 5.47139e-16
C3292 n1874_17 vss 5.47139e-16
C3293 n1874_16 vss 5.47139e-16
C3294 n1874_18 vss 5.47139e-16
C3295 n1874_17 vss 5.47139e-16
C3296 n1874_19 vss 5.47139e-16
C3297 n1874_18 vss 5.47139e-16
C3298 n1874_20 vss 5.47139e-16
C3299 n1874_19 vss 5.47139e-16
C3300 n1874_21 vss 5.47139e-16
C3301 n1874_20 vss 5.47139e-16
C3302 n1874_32 vss 1.40901e-17
C3303 n1874_31 vss 1.40901e-17
C3304 n1874_33 vss 3.91392e-17
C3305 n1874_32 vss 3.91392e-17
C3306 n1874_34 vss 3.91392e-17
C3307 n1874_33 vss 3.91392e-17
C3308 n1874_35 vss 4.6967e-17
C3309 n1874_34 vss 4.6967e-17
C3310 n1874_36 vss 3.91392e-17
C3311 n1874_35 vss 3.91392e-17
C3312 n1874_37 vss 2.42663e-16
C3313 n1874_36 vss 2.42663e-16
C3314 n1874_38 vss 3.91392e-17
C3315 n1874_37 vss 3.91392e-17
C3316 n1874_39 vss 3.91392e-17
C3317 n1874_38 vss 3.91392e-17
C3318 n1874_40 vss 3.91392e-17
C3319 n1874_39 vss 3.91392e-17
C3320 n1874_41 vss 3.91392e-17
C3321 n1874_40 vss 3.91392e-17
C3322 n1874_84 vss 1.0959e-16
C3323 n1874_41 vss 1.0959e-16
C3324 n1874_43 vss 1.40901e-17
C3325 n1874_42 vss 1.40901e-17
C3326 n1874_44 vss 3.91392e-17
C3327 n1874_43 vss 3.91392e-17
C3328 n1874_45 vss 3.91392e-17
C3329 n1874_44 vss 3.91392e-17
C3330 n1874_46 vss 3.91392e-17
C3331 n1874_45 vss 3.91392e-17
C3332 n1874_47 vss 3.91392e-17
C3333 n1874_46 vss 3.91392e-17
C3334 n1874_82 vss 1.0959e-16
C3335 n1874_47 vss 1.0959e-16
C3336 n1874_49 vss 1.40901e-17
C3337 n1874_48 vss 1.40901e-17
C3338 n1874_50 vss 3.91392e-17
C3339 n1874_49 vss 3.91392e-17
C3340 n1874_51 vss 3.91392e-17
C3341 n1874_50 vss 3.91392e-17
C3342 n1874_52 vss 4.6967e-17
C3343 n1874_51 vss 4.6967e-17
C3344 n1874_53 vss 3.91392e-17
C3345 n1874_52 vss 3.91392e-17
C3346 n1874_54 vss 2.42663e-16
C3347 n1874_53 vss 2.42663e-16
C3348 n1874_55 vss 3.91392e-17
C3349 n1874_54 vss 3.91392e-17
C3350 n1874_56 vss 3.91392e-17
C3351 n1874_55 vss 3.91392e-17
C3352 n1874_57 vss 3.91392e-17
C3353 n1874_56 vss 3.91392e-17
C3354 n1874_58 vss 3.91392e-17
C3355 n1874_57 vss 3.91392e-17
C3356 n1874_83 vss 1.0959e-16
C3357 n1874_58 vss 1.0959e-16
C3358 n1874_60 vss 1.40901e-17
C3359 n1874_59 vss 1.40901e-17
C3360 n1874_61 vss 3.91392e-17
C3361 n1874_60 vss 3.91392e-17
C3362 n1874_62 vss 3.91392e-17
C3363 n1874_61 vss 3.91392e-17
C3364 n1874_63 vss 3.91392e-17
C3365 n1874_62 vss 3.91392e-17
C3366 n1874_64 vss 3.91392e-17
C3367 n1874_63 vss 3.91392e-17
C3368 n1874_80 vss 1.0959e-16
C3369 n1874_64 vss 1.0959e-16
C3370 n1874_66 vss 1.40901e-17
C3371 n1874_65 vss 1.40901e-17
C3372 n1874_67 vss 3.91392e-17
C3373 n1874_66 vss 3.91392e-17
C3374 n1874_68 vss 3.91392e-17
C3375 n1874_67 vss 3.91392e-17
C3376 n1874_69 vss 3.91392e-17
C3377 n1874_68 vss 3.91392e-17
C3378 n1874_70 vss 3.91392e-17
C3379 n1874_69 vss 3.91392e-17
C3380 n1874_79 vss 1.0959e-16
C3381 n1874_70 vss 1.0959e-16
C3382 n1874_72 vss 1.40901e-17
C3383 n1874_71 vss 1.40901e-17
C3384 n1874_73 vss 3.91392e-17
C3385 n1874_72 vss 3.91392e-17
C3386 n1874_74 vss 3.91392e-17
C3387 n1874_73 vss 3.91392e-17
C3388 n1874_75 vss 3.91392e-17
C3389 n1874_74 vss 3.91392e-17
C3390 n1874_76 vss 3.91392e-17
C3391 n1874_75 vss 3.91392e-17
C3392 n1874_81 vss 1.0959e-16
C3393 n1874_76 vss 1.0959e-16
C3394 n1874_77 vss 3.71822e-17
C3395 n1874_91 vss 3.71822e-17
C3396 n1874_78 vss 1.40901e-17
C3397 n1874_77 vss 1.40901e-17
C3398 n1874_80 vss 9.39341e-17
C3399 n1874_79 vss 9.39341e-17
C3400 n1874_81 vss 9.39341e-17
C3401 n1874_80 vss 9.39341e-17
C3402 n1874_82 vss 9.39341e-17
C3403 n1874_81 vss 9.39341e-17
C3404 n1874_83 vss 9.39341e-17
C3405 n1874_82 vss 9.39341e-17
C3406 n1874_84 vss 9.39341e-17
C3407 n1874_83 vss 9.39341e-17
C3408 n1874_102 vss 9.39341e-17
C3409 n1874_84 vss 9.39341e-17
C3410 n1874_86 vss 1.40901e-17
C3411 n1874_85 vss 1.40901e-17
C3412 n1874_87 vss 3.91392e-17
C3413 n1874_86 vss 3.91392e-17
C3414 n1874_88 vss 3.91392e-17
C3415 n1874_87 vss 3.91392e-17
C3416 n1874_89 vss 4.6967e-17
C3417 n1874_88 vss 4.6967e-17
C3418 n1874_90 vss 3.91392e-17
C3419 n1874_89 vss 3.91392e-17
C3420 n1874_91 vss 4.6967e-17
C3421 n1874_90 vss 4.6967e-17
C3422 n1874_92 vss 6.41883e-17
C3423 n1874_91 vss 6.41883e-17
C3424 n1874_93 vss 2.81802e-17
C3425 n1874_92 vss 2.81802e-17
C3426 n1874_94 vss 5.63604e-17
C3427 n1874_93 vss 5.63604e-17
C3428 n1874_97 vss 4.6967e-17
C3429 n1874_94 vss 4.6967e-17
C3430 n1874_98 vss 3.91392e-17
C3431 n1874_97 vss 3.91392e-17
C3432 n1874_99 vss 3.91392e-17
C3433 n1874_98 vss 3.91392e-17
C3434 n1874_100 vss 3.91392e-17
C3435 n1874_99 vss 3.91392e-17
C3436 n1874_101 vss 3.91392e-17
C3437 n1874_100 vss 3.91392e-17
C3438 n1874_102 vss 1.0959e-16
C3439 n1874_101 vss 1.0959e-16
C3440 n1874_95 vss 3.71822e-17
C3441 n1874_94 vss 3.71822e-17
C3442 n1874_96 vss 1.40901e-17
C3443 n1874_95 vss 1.40901e-17
C3444 n1874_3 vss 4.20552e-17
C3445 n1874_2 vss 4.20552e-17
C3446 n1874_4 vss 9.46242e-17
C3447 n1874_3 vss 9.46242e-17
C3448 n1874_5 vss 3.05111e-16
C3449 n1874_4 vss 3.05111e-16
C3450 n1874_6 vss 3.05111e-16
C3451 n1874_5 vss 3.05111e-16
C3452 n1874_7 vss 3.05111e-16
C3453 n1874_6 vss 3.05111e-16
C3454 n1874_8 vss 3.05111e-16
C3455 n1874_7 vss 3.05111e-16
C3456 n1874_9 vss 3.05111e-16
C3457 n1874_8 vss 3.05111e-16
C3458 n1874_10 vss 3.05111e-16
C3459 n1874_9 vss 3.05111e-16
C3460 n1874_11 vss 3.05111e-16
C3461 n1874_10 vss 3.05111e-16

R56_1 n1981_2 n1981_33 0.001
R56_2 n1981_20 n1981_6 0.001
R56_3 n1981_1 n1981_32 0.001
R56_4 n1981_29 n1981_5 0.001
R56_5 n1981_38 n1981_9 0.001
R56_6 n1981_39 n1981_9 0.001
R56_7 n1981_36 n1981_9 0.001
R56_8 n1981_37 n1981_9 0.001
R56_9 n1981_35 n1981_9 0.001
R56_10 n1981_27 n1981_10 0.001
R56_11 n1981_28 n1981_10 0.001
R56_12 n1981_26 n1981_10 0.001
R56_13 n1981_24 n1981_10 0.001
R56_14 n1981_25 n1981_12 0.001
R56_15 n1981_16 n1981_13 0.001
R56_16 n1981_18 n1981_13 0.001
R56_17 n1981_17 n1981_13 0.001
R56_18 n1981_11 n1981_15 0.001
R56_19 n1981_14 n1981_13 0.001
R56_20 n1981_6 n1981_5 7.2
R56_21 n1981_7 n1981_6 21.6
R56_22 n1981 n1981_7 0.001
R56_23 n1981_14 n1981_22 0.324
R56_24 n1981_15 n1981_14 0.108
R56_25 n1981_16 n1981_15 0.108
R56_26 n1981_17 n1981_16 0.108
R56_27 n1981_18 n1981_17 0.108
R56_28 n1981_19 n1981_18 0.001
R56_29 n1981_12 n1981_11 0.216
R56_30 n1981_20 n1981_29 0.108
R56_31 n1981_21 n1981_20 0.001
R56_32 n1981_23 n1981_22 0.324
R56_33 n1981_24 n1981_23 0.324
R56_34 n1981_25 n1981_24 0.108
R56_35 n1981_26 n1981_25 0.108
R56_36 n1981_27 n1981_26 0.108
R56_37 n1981_28 n1981_27 0.108
R56_38 n1981_29 n1981_28 0.108
R56_39 n1981_30 n1981_29 0.216
R56_40 n1981_31 n1981_30 0.108
R56_41 n1981_32 n1981_31 0.216
R56_42 n1981_35 n1981_32 0.108
R56_43 n1981_36 n1981_35 0.108
R56_44 n1981_37 n1981_36 0.108
R56_45 n1981_38 n1981_37 0.108
R56_46 n1981_39 n1981_38 0.108
R56_47 n1981_40 n1981_39 0.001
R56_48 n1981_33 n1981_32 0.108
R56_49 n1981_34 n1981_33 0.001
R56_50 n1981_2 n1981_1 7.2
R56_51 n1981_3 n1981_2 21.6
R56_52 n1981_4 n1981_3 0.001

C3462 n1981_6 vss 4.20552e-17
C3463 n1981_5 vss 4.20552e-17
C3464 n1981_7 vss 9.46242e-17
C3465 n1981_6 vss 9.46242e-17
C3466 n1981 vss 3.05111e-16
C3467 n1981_7 vss 3.05111e-16
C3468 n1981_14 vss 1.0959e-16
C3469 n1981_22 vss 1.0959e-16
C3470 n1981_15 vss 3.91392e-17
C3471 n1981_14 vss 3.91392e-17
C3472 n1981_16 vss 3.91392e-17
C3473 n1981_15 vss 3.91392e-17
C3474 n1981_17 vss 3.91392e-17
C3475 n1981_16 vss 3.91392e-17
C3476 n1981_18 vss 3.91392e-17
C3477 n1981_17 vss 3.91392e-17
C3478 n1981_19 vss 1.40901e-17
C3479 n1981_18 vss 1.40901e-17
C3480 n1981_12 vss 7.81488e-17
C3481 n1981_11 vss 7.81488e-17
C3482 n1981_20 vss 3.71822e-17
C3483 n1981_29 vss 3.71822e-17
C3484 n1981_21 vss 1.40901e-17
C3485 n1981_20 vss 1.40901e-17
C3486 n1981_23 vss 9.39341e-17
C3487 n1981_22 vss 9.39341e-17
C3488 n1981_24 vss 1.0959e-16
C3489 n1981_23 vss 1.0959e-16
C3490 n1981_25 vss 3.91392e-17
C3491 n1981_24 vss 3.91392e-17
C3492 n1981_26 vss 3.91392e-17
C3493 n1981_25 vss 3.91392e-17
C3494 n1981_27 vss 3.91392e-17
C3495 n1981_26 vss 3.91392e-17
C3496 n1981_28 vss 3.91392e-17
C3497 n1981_27 vss 3.91392e-17
C3498 n1981_29 vss 4.6967e-17
C3499 n1981_28 vss 4.6967e-17
C3500 n1981_30 vss 5.63604e-17
C3501 n1981_29 vss 5.63604e-17
C3502 n1981_31 vss 2.81802e-17
C3503 n1981_30 vss 2.81802e-17
C3504 n1981_32 vss 6.41883e-17
C3505 n1981_31 vss 6.41883e-17
C3506 n1981_35 vss 4.6967e-17
C3507 n1981_32 vss 4.6967e-17
C3508 n1981_36 vss 3.91392e-17
C3509 n1981_35 vss 3.91392e-17
C3510 n1981_37 vss 4.6967e-17
C3511 n1981_36 vss 4.6967e-17
C3512 n1981_38 vss 3.91392e-17
C3513 n1981_37 vss 3.91392e-17
C3514 n1981_39 vss 3.91392e-17
C3515 n1981_38 vss 3.91392e-17
C3516 n1981_40 vss 1.40901e-17
C3517 n1981_39 vss 1.40901e-17
C3518 n1981_33 vss 3.71822e-17
C3519 n1981_32 vss 3.71822e-17
C3520 n1981_34 vss 1.40901e-17
C3521 n1981_33 vss 1.40901e-17
C3522 n1981_2 vss 4.20552e-17
C3523 n1981_1 vss 4.20552e-17
C3524 n1981_3 vss 9.46242e-17
C3525 n1981_2 vss 9.46242e-17
C3526 n1981_4 vss 5.47139e-16
C3527 n1981_3 vss 5.47139e-16

R2_1 a_3_50 a_3_1 0.001
R2_2 a_3_48 a_3_1 0.001
R2_3 a_3_49 a_3_1 0.001
R2_4 a_3_47 a_3_1 0.001
R2_5 a_3_46 a_3_1 0.001
R2_6 a_3_45 a_3_1 0.001
R2_7 a_3_44 a_3_1 0.001
R2_8 a_3_43 a_3_1 0.001
R2_9 a_3_42 a_3_2 0.001
R2_10 a_3_41 a_3_2 0.001
R2_11 a_3_39 a_3_2 0.001
R2_12 a_3_40 a_3_2 0.001
R2_13 a_3_36 a_3_2 0.001
R2_14 a_3_38 a_3_2 0.001
R2_15 a_3_37 a_3_2 0.001
R2_16 a_3_34 a_3_2 0.001
R2_17 a_3_35 a_3_2 0.001
R2_18 a_3_33 a_3_2 0.001
R2_19 a_3_32 a_3_2 0.001
R2_20 a_3_30 a_3_2 0.001
R2_21 a_3_31 a_3_2 0.001
R2_22 a_3_29 a_3_2 0.001
R2_23 a_3_28 a_3_2 0.001
R2_24 a_3_27 a_3_2 0.001
R2_25 a_3_26 a_3_2 0.001
R2_26 a_3_25 a_3_2 0.001
R2_27 a_3_24 a_3_2 0.001
R2_28 a_3_23 a_3_2 0.001
R2_29 a_3_79 a_3_3 0.001
R2_30 a_3_77 a_3_3 0.001
R2_31 a_3_78 a_3_3 0.001
R2_32 a_3_76 a_3_3 0.001
R2_33 a_3_75 a_3_3 0.001
R2_34 a_3_73 a_3_3 0.001
R2_35 a_3_74 a_3_3 0.001
R2_36 a_3_72 a_3_3 0.001
R2_37 a_3_71 a_3_4 0.001
R2_38 a_3_70 a_3_4 0.001
R2_39 a_3_68 a_3_4 0.001
R2_40 a_3_69 a_3_4 0.001
R2_41 a_3_65 a_3_4 0.001
R2_42 a_3_67 a_3_4 0.001
R2_43 a_3_66 a_3_4 0.001
R2_44 a_3_64 a_3_4 0.001
R2_45 a_3_63 a_3_4 0.001
R2_46 a_3_61 a_3_4 0.001
R2_47 a_3_62 a_3_4 0.001
R2_48 a_3_59 a_3_4 0.001
R2_49 a_3_60 a_3_4 0.001
R2_50 a_3_58 a_3_4 0.001
R2_51 a_3_57 a_3_4 0.001
R2_52 a_3_56 a_3_4 0.001
R2_53 a_3_55 a_3_4 0.001
R2_54 a_3_54 a_3_4 0.001
R2_55 a_3_53 a_3_4 0.001
R2_56 a_3_52 a_3_4 0.001
R2_57 a_3_14 a_3_5 0.001
R2_58 a_3_13 a_3_8 0.001
R2_59 a_3 a_3_11 0.001
R2_60 a_3_6 a_3_5 21.6
R2_61 a_3_8 a_3_7 7.2
R2_62 a_3_9 a_3_8 7.2
R2_63 a_3_10 a_3_9 14.4
R2_64 a_3_13 a_3_12 0.001
R2_65 a_3_16 a_3_13 0.216
R2_66 a_3_14 a_3_16 0.216
R2_67 a_3_15 a_3_14 0.001
R2_68 a_3_16 a_3_17 0.324
R2_69 a_3_18 a_3_17 2.268
R2_70 a_3_19 a_3_18 1.08
R2_71 a_3_20 a_3_19 0.001
R2_72 a_3_21 a_3_20 0.001
R2_73 a_3_51 a_3_21 0.216
R2_74 a_3_23 a_3_22 0.001
R2_75 a_3_24 a_3_23 0.108
R2_76 a_3_25 a_3_24 0.108
R2_77 a_3_26 a_3_25 0.108
R2_78 a_3_27 a_3_26 0.108
R2_79 a_3_28 a_3_27 0.108
R2_80 a_3_29 a_3_28 0.108
R2_81 a_3_30 a_3_29 0.108
R2_82 a_3_31 a_3_30 0.108
R2_83 a_3_32 a_3_31 0.108
R2_84 a_3_33 a_3_32 0.108
R2_85 a_3_34 a_3_33 0.108
R2_86 a_3_35 a_3_34 0.108
R2_87 a_3_36 a_3_35 0.108
R2_88 a_3_37 a_3_36 0.108
R2_89 a_3_38 a_3_37 0.108
R2_90 a_3_39 a_3_38 0.108
R2_91 a_3_40 a_3_39 0.108
R2_92 a_3_41 a_3_40 0.108
R2_93 a_3_42 a_3_41 0.108
R2_94 a_3_43 a_3_42 0.864
R2_95 a_3_44 a_3_43 0.108
R2_96 a_3_45 a_3_44 0.108
R2_97 a_3_46 a_3_45 0.108
R2_98 a_3_47 a_3_46 0.108
R2_99 a_3_48 a_3_47 0.108
R2_100 a_3_49 a_3_48 0.108
R2_101 a_3_50 a_3_49 0.108
R2_102 a_3_81 a_3_50 0.54
R2_103 a_3_52 a_3_51 0.001
R2_104 a_3_53 a_3_52 0.108
R2_105 a_3_54 a_3_53 0.108
R2_106 a_3_55 a_3_54 0.108
R2_107 a_3_56 a_3_55 0.108
R2_108 a_3_57 a_3_56 0.108
R2_109 a_3_58 a_3_57 0.108
R2_110 a_3_59 a_3_58 0.108
R2_111 a_3_60 a_3_59 0.108
R2_112 a_3_61 a_3_60 0.108
R2_113 a_3_62 a_3_61 0.108
R2_114 a_3_63 a_3_62 0.108
R2_115 a_3_64 a_3_63 0.108
R2_116 a_3_65 a_3_64 0.108
R2_117 a_3_66 a_3_65 0.108
R2_118 a_3_67 a_3_66 0.108
R2_119 a_3_68 a_3_67 0.108
R2_120 a_3_69 a_3_68 0.108
R2_121 a_3_70 a_3_69 0.108
R2_122 a_3_71 a_3_70 0.108
R2_123 a_3_72 a_3_71 0.864
R2_124 a_3_73 a_3_72 0.108
R2_125 a_3_74 a_3_73 0.108
R2_126 a_3_75 a_3_74 0.108
R2_127 a_3_76 a_3_75 0.108
R2_128 a_3_77 a_3_76 0.108
R2_129 a_3_78 a_3_77 0.108
R2_130 a_3_79 a_3_78 0.108
R2_131 a_3_82 a_3_79 0.54
R2_132 a_3_82 a_3_80 0.001
R2_133 a_3_81 a_3_82 0.108
R2_134 a_3_83 a_3_82 0.54
R2_135 a_3_84 a_3_83 0.001
R2_136 a_3 a_3_84 0.001

C3528 a_3_6 vss 9.46242e-17
C3529 a_3_5 vss 9.46242e-17
C3530 a_3_8 vss 3.15414e-17
C3531 a_3_7 vss 3.15414e-17
C3532 a_3_9 vss 3.15414e-17
C3533 a_3_8 vss 3.15414e-17
C3534 a_3_10 vss 6.30828e-17
C3535 a_3_9 vss 6.30828e-17
C3536 a_3_13 vss 1.40901e-17
C3537 a_3_12 vss 1.40901e-17
C3538 a_3_16 vss 7.82784e-17
C3539 a_3_13 vss 7.82784e-17
C3540 a_3_14 vss 7.04506e-17
C3541 a_3_16 vss 7.04506e-17
C3542 a_3_15 vss 1.40901e-17
C3543 a_3_14 vss 1.40901e-17
C3544 a_3_16 vss 9.39341e-17
C3545 a_3_17 vss 9.39341e-17
C3546 a_3_18 vss 6.18399e-16
C3547 a_3_17 vss 6.18399e-16
C3548 a_3_19 vss 2.97458e-16
C3549 a_3_18 vss 2.97458e-16
C3550 a_3_20 vss 2.50491e-17
C3551 a_3_19 vss 2.50491e-17
C3552 a_3_21 vss 1.25245e-17
C3553 a_3_20 vss 1.25245e-17
C3554 a_3_51 vss 8.14095e-17
C3555 a_3_21 vss 8.14095e-17
C3556 a_3_23 vss 1.40901e-17
C3557 a_3_22 vss 1.40901e-17
C3558 a_3_24 vss 3.13114e-17
C3559 a_3_23 vss 3.13114e-17
C3560 a_3_25 vss 3.13114e-17
C3561 a_3_24 vss 3.13114e-17
C3562 a_3_26 vss 3.13114e-17
C3563 a_3_25 vss 3.13114e-17
C3564 a_3_27 vss 3.13114e-17
C3565 a_3_26 vss 3.13114e-17
C3566 a_3_28 vss 3.13114e-17
C3567 a_3_27 vss 3.13114e-17
C3568 a_3_29 vss 3.13114e-17
C3569 a_3_28 vss 3.13114e-17
C3570 a_3_30 vss 3.13114e-17
C3571 a_3_29 vss 3.13114e-17
C3572 a_3_31 vss 3.13114e-17
C3573 a_3_30 vss 3.13114e-17
C3574 a_3_32 vss 3.13114e-17
C3575 a_3_31 vss 3.13114e-17
C3576 a_3_33 vss 3.13114e-17
C3577 a_3_32 vss 3.13114e-17
C3578 a_3_34 vss 3.13114e-17
C3579 a_3_33 vss 3.13114e-17
C3580 a_3_35 vss 3.13114e-17
C3581 a_3_34 vss 3.13114e-17
C3582 a_3_36 vss 3.13114e-17
C3583 a_3_35 vss 3.13114e-17
C3584 a_3_37 vss 3.13114e-17
C3585 a_3_36 vss 3.13114e-17
C3586 a_3_38 vss 3.13114e-17
C3587 a_3_37 vss 3.13114e-17
C3588 a_3_39 vss 3.13114e-17
C3589 a_3_38 vss 3.13114e-17
C3590 a_3_40 vss 3.13114e-17
C3591 a_3_39 vss 3.13114e-17
C3592 a_3_41 vss 3.13114e-17
C3593 a_3_40 vss 3.13114e-17
C3594 a_3_42 vss 3.13114e-17
C3595 a_3_41 vss 3.13114e-17
C3596 a_3_43 vss 2.42663e-16
C3597 a_3_42 vss 2.42663e-16
C3598 a_3_44 vss 3.13114e-17
C3599 a_3_43 vss 3.13114e-17
C3600 a_3_45 vss 3.13114e-17
C3601 a_3_44 vss 3.13114e-17
C3602 a_3_46 vss 3.13114e-17
C3603 a_3_45 vss 3.13114e-17
C3604 a_3_47 vss 3.13114e-17
C3605 a_3_46 vss 3.13114e-17
C3606 a_3_48 vss 3.13114e-17
C3607 a_3_47 vss 3.13114e-17
C3608 a_3_49 vss 3.13114e-17
C3609 a_3_48 vss 3.13114e-17
C3610 a_3_50 vss 3.13114e-17
C3611 a_3_49 vss 3.13114e-17
C3612 a_3_81 vss 1.40901e-16
C3613 a_3_50 vss 1.40901e-16
C3614 a_3_52 vss 1.40901e-17
C3615 a_3_51 vss 1.40901e-17
C3616 a_3_53 vss 3.13114e-17
C3617 a_3_52 vss 3.13114e-17
C3618 a_3_54 vss 3.13114e-17
C3619 a_3_53 vss 3.13114e-17
C3620 a_3_55 vss 3.13114e-17
C3621 a_3_54 vss 3.13114e-17
C3622 a_3_56 vss 3.13114e-17
C3623 a_3_55 vss 3.13114e-17
C3624 a_3_57 vss 3.13114e-17
C3625 a_3_56 vss 3.13114e-17
C3626 a_3_58 vss 3.13114e-17
C3627 a_3_57 vss 3.13114e-17
C3628 a_3_59 vss 3.13114e-17
C3629 a_3_58 vss 3.13114e-17
C3630 a_3_60 vss 3.13114e-17
C3631 a_3_59 vss 3.13114e-17
C3632 a_3_61 vss 3.13114e-17
C3633 a_3_60 vss 3.13114e-17
C3634 a_3_62 vss 3.13114e-17
C3635 a_3_61 vss 3.13114e-17
C3636 a_3_63 vss 3.13114e-17
C3637 a_3_62 vss 3.13114e-17
C3638 a_3_64 vss 3.13114e-17
C3639 a_3_63 vss 3.13114e-17
C3640 a_3_65 vss 3.13114e-17
C3641 a_3_64 vss 3.13114e-17
C3642 a_3_66 vss 3.13114e-17
C3643 a_3_65 vss 3.13114e-17
C3644 a_3_67 vss 3.13114e-17
C3645 a_3_66 vss 3.13114e-17
C3646 a_3_68 vss 3.13114e-17
C3647 a_3_67 vss 3.13114e-17
C3648 a_3_69 vss 3.13114e-17
C3649 a_3_68 vss 3.13114e-17
C3650 a_3_70 vss 3.13114e-17
C3651 a_3_69 vss 3.13114e-17
C3652 a_3_71 vss 3.13114e-17
C3653 a_3_70 vss 3.13114e-17
C3654 a_3_72 vss 2.42663e-16
C3655 a_3_71 vss 2.42663e-16
C3656 a_3_73 vss 3.13114e-17
C3657 a_3_72 vss 3.13114e-17
C3658 a_3_74 vss 3.13114e-17
C3659 a_3_73 vss 3.13114e-17
C3660 a_3_75 vss 3.13114e-17
C3661 a_3_74 vss 3.13114e-17
C3662 a_3_76 vss 3.13114e-17
C3663 a_3_75 vss 3.13114e-17
C3664 a_3_77 vss 3.13114e-17
C3665 a_3_76 vss 3.13114e-17
C3666 a_3_78 vss 3.13114e-17
C3667 a_3_77 vss 3.13114e-17
C3668 a_3_79 vss 3.13114e-17
C3669 a_3_78 vss 3.13114e-17
C3670 a_3_82 vss 1.40901e-16
C3671 a_3_79 vss 1.40901e-16
C3672 a_3_82 vss 6.34418e-17
C3673 a_3_80 vss 6.34418e-17
C3674 a_3_81 vss 1.42197e-16
C3675 a_3_82 vss 1.42197e-16
C3676 a_3_83 vss 6.8969e-16
C3677 a_3_82 vss 6.8969e-16
C3678 a_3_84 vss 3.48676e-17
C3679 a_3_83 vss 3.48676e-17
C3680 a_3 vss 4.3846e-15
C3681 a_3_84 vss 4.3846e-15

R57_1 n2124_2 n2124_30 0.001
R57_2 n2124_20 n2124_6 0.001
R57_3 n2124_1 n2124_34 0.001
R57_4 n2124_29 n2124_5 0.001
R57_5 n2124_39 n2124_9 0.001
R57_6 n2124_38 n2124_12 0.001
R57_7 n2124_36 n2124_9 0.001
R57_8 n2124_37 n2124_9 0.001
R57_9 n2124_35 n2124_9 0.001
R57_10 n2124_28 n2124_10 0.001
R57_11 n2124_26 n2124_10 0.001
R57_12 n2124_27 n2124_10 0.001
R57_13 n2124_25 n2124_10 0.001
R57_14 n2124_24 n2124_10 0.001
R57_15 n2124_11 n2124_18 0.001
R57_16 n2124_19 n2124_13 0.001
R57_17 n2124_17 n2124_13 0.001
R57_18 n2124_16 n2124_13 0.001
R57_19 n2124_15 n2124_13 0.001
R57_20 n2124_6 n2124_5 7.2
R57_21 n2124_7 n2124_6 21.6
R57_22 n2124_8 n2124_7 0.001
R57_23 n2124_15 n2124_14 0.001
R57_24 n2124_16 n2124_15 0.108
R57_25 n2124_17 n2124_16 0.108
R57_26 n2124_18 n2124_17 0.108
R57_27 n2124_19 n2124_18 0.108
R57_28 n2124_22 n2124_19 0.324
R57_29 n2124_12 n2124_11 0.216
R57_30 n2124_20 n2124_29 0.108
R57_31 n2124_21 n2124_20 0.001
R57_32 n2124_40 n2124_22 0.324
R57_33 n2124_24 n2124_23 0.001
R57_34 n2124_25 n2124_24 0.108
R57_35 n2124_26 n2124_25 0.108
R57_36 n2124_27 n2124_26 0.108
R57_37 n2124_28 n2124_27 0.108
R57_38 n2124_29 n2124_28 0.108
R57_39 n2124_32 n2124_29 0.216
R57_40 n2124_30 n2124_34 0.108
R57_41 n2124_31 n2124_30 0.001
R57_42 n2124_33 n2124_32 0.108
R57_43 n2124_34 n2124_33 0.216
R57_44 n2124_35 n2124_34 0.108
R57_45 n2124_36 n2124_35 0.108
R57_46 n2124_37 n2124_36 0.108
R57_47 n2124_38 n2124_37 0.108
R57_48 n2124_39 n2124_38 0.108
R57_49 n2124_40 n2124_39 0.324
R57_50 n2124_2 n2124_1 7.2
R57_51 n2124_3 n2124_2 21.6
R57_52 n2124 n2124_3 0.001

C3682 n2124_6 vss 4.20552e-17
C3683 n2124_5 vss 4.20552e-17
C3684 n2124_7 vss 9.46242e-17
C3685 n2124_6 vss 9.46242e-17
C3686 n2124_8 vss 5.47139e-16
C3687 n2124_7 vss 5.47139e-16
C3688 n2124_15 vss 1.40901e-17
C3689 n2124_14 vss 1.40901e-17
C3690 n2124_16 vss 3.91392e-17
C3691 n2124_15 vss 3.91392e-17
C3692 n2124_17 vss 3.91392e-17
C3693 n2124_16 vss 3.91392e-17
C3694 n2124_18 vss 3.91392e-17
C3695 n2124_17 vss 3.91392e-17
C3696 n2124_19 vss 3.91392e-17
C3697 n2124_18 vss 3.91392e-17
C3698 n2124_22 vss 1.0959e-16
C3699 n2124_19 vss 1.0959e-16
C3700 n2124_12 vss 7.81488e-17
C3701 n2124_11 vss 7.81488e-17
C3702 n2124_20 vss 3.71822e-17
C3703 n2124_29 vss 3.71822e-17
C3704 n2124_21 vss 1.40901e-17
C3705 n2124_20 vss 1.40901e-17
C3706 n2124_40 vss 9.39341e-17
C3707 n2124_22 vss 9.39341e-17
C3708 n2124_24 vss 1.40901e-17
C3709 n2124_23 vss 1.40901e-17
C3710 n2124_25 vss 3.91392e-17
C3711 n2124_24 vss 3.91392e-17
C3712 n2124_26 vss 3.91392e-17
C3713 n2124_25 vss 3.91392e-17
C3714 n2124_27 vss 4.6967e-17
C3715 n2124_26 vss 4.6967e-17
C3716 n2124_28 vss 3.91392e-17
C3717 n2124_27 vss 3.91392e-17
C3718 n2124_29 vss 4.6967e-17
C3719 n2124_28 vss 4.6967e-17
C3720 n2124_32 vss 6.41883e-17
C3721 n2124_29 vss 6.41883e-17
C3722 n2124_30 vss 3.71822e-17
C3723 n2124_34 vss 3.71822e-17
C3724 n2124_31 vss 1.40901e-17
C3725 n2124_30 vss 1.40901e-17
C3726 n2124_33 vss 2.81802e-17
C3727 n2124_32 vss 2.81802e-17
C3728 n2124_34 vss 5.63604e-17
C3729 n2124_33 vss 5.63604e-17
C3730 n2124_35 vss 4.6967e-17
C3731 n2124_34 vss 4.6967e-17
C3732 n2124_36 vss 3.91392e-17
C3733 n2124_35 vss 3.91392e-17
C3734 n2124_37 vss 3.91392e-17
C3735 n2124_36 vss 3.91392e-17
C3736 n2124_38 vss 3.91392e-17
C3737 n2124_37 vss 3.91392e-17
C3738 n2124_39 vss 3.91392e-17
C3739 n2124_38 vss 3.91392e-17
C3740 n2124_40 vss 1.0959e-16
C3741 n2124_39 vss 1.0959e-16
C3742 n2124_2 vss 4.20552e-17
C3743 n2124_1 vss 4.20552e-17
C3744 n2124_3 vss 9.46242e-17
C3745 n2124_2 vss 9.46242e-17
C3746 n2124 vss 3.05111e-16
C3747 n2124_3 vss 3.05111e-16

R58_1 n2145_1 n2145_4 0.001
R58_2 n2145_3 n2145 0.001
R58_3 n2145_4 n2145_3 0.756

C3748 n2145_4 vss 8.14925e-17
C3749 n2145_3 vss 8.14925e-17

R59_1 n2151_1 n2151_4 0.001
R59_2 n2151_3 n2151 0.001
R59_3 n2151_4 n2151_3 0.756

C3750 n2151_4 vss 8.14925e-17
C3751 n2151_3 vss 8.14925e-17

R60_1 n2169_1 n2169_4 0.001
R60_2 n2169_3 n2169 0.001
R60_3 n2169_4 n2169_3 0.756

C3752 n2169_4 vss 8.14925e-17
C3753 n2169_3 vss 8.14925e-17

R61_1 n2181_1 n2181_4 0.001
R61_2 n2181_3 n2181 0.001
R61_3 n2181_4 n2181_3 0.756

C3754 n2181_4 vss 8.14925e-17
C3755 n2181_3 vss 8.14925e-17

R62_1 sel_49 sel_1 0.001
R62_2 sel_48 sel_1 0.001
R62_3 sel_47 sel_1 0.001
R62_4 sel_45 sel_1 0.001
R62_5 sel_46 sel_1 0.001
R62_6 sel_43 sel_1 0.001
R62_7 sel_44 sel_1 0.001
R62_8 sel_42 sel_1 0.001
R62_9 sel_41 sel_1 0.001
R62_10 sel_39 sel_1 0.001
R62_11 sel_40 sel_1 0.001
R62_12 sel_37 sel_1 0.001
R62_13 sel_38 sel_1 0.001
R62_14 sel_35 sel_1 0.001
R62_15 sel_36 sel_1 0.001
R62_16 sel_34 sel_1 0.001
R62_17 sel_33 sel_1 0.001
R62_18 sel_31 sel_1 0.001
R62_19 sel_32 sel_1 0.001
R62_20 sel_30 sel_1 0.001
R62_21 sel_29 sel_2 0.001
R62_22 sel_27 sel_2 0.001
R62_23 sel_28 sel_2 0.001
R62_24 sel_25 sel_2 0.001
R62_25 sel_26 sel_2 0.001
R62_26 sel_23 sel_2 0.001
R62_27 sel_24 sel_2 0.001
R62_28 sel_22 sel_2 0.001
R62_29 sel_84 sel_3 0.001
R62_30 sel_83 sel_3 0.001
R62_31 sel_82 sel_3 0.001
R62_32 sel_80 sel_3 0.001
R62_33 sel_81 sel_3 0.001
R62_34 sel_78 sel_3 0.001
R62_35 sel_79 sel_3 0.001
R62_36 sel_76 sel_3 0.001
R62_37 sel_77 sel_3 0.001
R62_38 sel_74 sel_3 0.001
R62_39 sel_75 sel_3 0.001
R62_40 sel_72 sel_3 0.001
R62_41 sel_73 sel_3 0.001
R62_42 sel_70 sel_3 0.001
R62_43 sel_71 sel_3 0.001
R62_44 sel_69 sel_3 0.001
R62_45 sel_68 sel_3 0.001
R62_46 sel_66 sel_3 0.001
R62_47 sel_67 sel_3 0.001
R62_48 sel_65 sel_3 0.001
R62_49 sel_64 sel_4 0.001
R62_50 sel_62 sel_4 0.001
R62_51 sel_63 sel_4 0.001
R62_52 sel_61 sel_4 0.001
R62_53 sel_60 sel_4 0.001
R62_54 sel_58 sel_4 0.001
R62_55 sel_59 sel_4 0.001
R62_56 sel_57 sel_4 0.001
R62_57 sel_14 sel_6 0.001
R62_58 sel_13 sel_9 0.001
R62_59 sel sel_11 0.001
R62_60 sel_6 sel_5 7.2
R62_61 sel_7 sel_6 7.2
R62_62 sel_8 sel_7 14.4
R62_63 sel_10 sel_9 21.6
R62_64 sel_13 sel_12 0.001
R62_65 sel_16 sel_13 0.216
R62_66 sel_14 sel_16 0.216
R62_67 sel_15 sel_14 0.001
R62_68 sel_16 sel_17 0.324
R62_69 sel_17 sel_18 2.268
R62_70 sel_19 sel_18 1.08
R62_71 sel_19 sel_21 0.001
R62_72 sel_20 sel_85 0.216
R62_73 sel_21 sel_20 0.001
R62_74 sel_22 sel_52 0.54
R62_75 sel_23 sel_22 0.108
R62_76 sel_24 sel_23 0.108
R62_77 sel_25 sel_24 0.108
R62_78 sel_26 sel_25 0.108
R62_79 sel_27 sel_26 0.108
R62_80 sel_28 sel_27 0.108
R62_81 sel_29 sel_28 0.108
R62_82 sel_30 sel_29 0.864
R62_83 sel_31 sel_30 0.108
R62_84 sel_32 sel_31 0.108
R62_85 sel_33 sel_32 0.108
R62_86 sel_34 sel_33 0.108
R62_87 sel_35 sel_34 0.108
R62_88 sel_36 sel_35 0.108
R62_89 sel_37 sel_36 0.108
R62_90 sel_38 sel_37 0.108
R62_91 sel_39 sel_38 0.108
R62_92 sel_40 sel_39 0.108
R62_93 sel_41 sel_40 0.108
R62_94 sel_42 sel_41 0.108
R62_95 sel_43 sel_42 0.108
R62_96 sel_44 sel_43 0.108
R62_97 sel_45 sel_44 0.108
R62_98 sel_46 sel_45 0.108
R62_99 sel_47 sel_46 0.108
R62_100 sel_48 sel_47 0.108
R62_101 sel_49 sel_48 0.108
R62_102 sel_50 sel_49 0.001
R62_103 sel_57 sel_53 0.54
R62_104 sel_58 sel_57 0.108
R62_105 sel_59 sel_58 0.108
R62_106 sel_60 sel_59 0.108
R62_107 sel_61 sel_60 0.108
R62_108 sel_62 sel_61 0.108
R62_109 sel_63 sel_62 0.108
R62_110 sel_64 sel_63 0.108
R62_111 sel_65 sel_64 0.864
R62_112 sel_66 sel_65 0.108
R62_113 sel_67 sel_66 0.108
R62_114 sel_68 sel_67 0.108
R62_115 sel_69 sel_68 0.108
R62_116 sel_70 sel_69 0.108
R62_117 sel_71 sel_70 0.108
R62_118 sel_72 sel_71 0.108
R62_119 sel_73 sel_72 0.108
R62_120 sel_74 sel_73 0.108
R62_121 sel_75 sel_74 0.108
R62_122 sel_76 sel_75 0.108
R62_123 sel_77 sel_76 0.108
R62_124 sel_78 sel_77 0.108
R62_125 sel_79 sel_78 0.108
R62_126 sel_80 sel_79 0.108
R62_127 sel_81 sel_80 0.108
R62_128 sel_82 sel_81 0.108
R62_129 sel_83 sel_82 0.108
R62_130 sel_84 sel_83 0.108
R62_131 sel_85 sel_84 0.001
R62_132 sel_53 sel_51 0.001
R62_133 sel_52 sel_53 0.108
R62_134 sel_53 sel_56 0.54
R62_135 sel sel_55 0.001
R62_136 sel_56 sel_55 0.001

C3756 sel_6 vss 3.15414e-17
C3757 sel_5 vss 3.15414e-17
C3758 sel_7 vss 3.15414e-17
C3759 sel_6 vss 3.15414e-17
C3760 sel_8 vss 6.30828e-17
C3761 sel_7 vss 6.30828e-17
C3762 sel_10 vss 9.46242e-17
C3763 sel_9 vss 9.46242e-17
C3764 sel_13 vss 1.40901e-17
C3765 sel_12 vss 1.40901e-17
C3766 sel_16 vss 7.04506e-17
C3767 sel_13 vss 7.04506e-17
C3768 sel_14 vss 7.82784e-17
C3769 sel_16 vss 7.82784e-17
C3770 sel_15 vss 1.40901e-17
C3771 sel_14 vss 1.40901e-17
C3772 sel_16 vss 9.39341e-17
C3773 sel_17 vss 9.39341e-17
C3774 sel_17 vss 6.18399e-16
C3775 sel_18 vss 6.18399e-16
C3776 sel_19 vss 2.97458e-16
C3777 sel_18 vss 2.97458e-16
C3778 sel_19 vss 2.50491e-17
C3779 sel_21 vss 2.50491e-17
C3780 sel_20 vss 8.14095e-17
C3781 sel_85 vss 8.14095e-17
C3782 sel_21 vss 1.25245e-17
C3783 sel_20 vss 1.25245e-17
C3784 sel_22 vss 1.40901e-16
C3785 sel_52 vss 1.40901e-16
C3786 sel_23 vss 3.13114e-17
C3787 sel_22 vss 3.13114e-17
C3788 sel_24 vss 3.13114e-17
C3789 sel_23 vss 3.13114e-17
C3790 sel_25 vss 3.13114e-17
C3791 sel_24 vss 3.13114e-17
C3792 sel_26 vss 3.13114e-17
C3793 sel_25 vss 3.13114e-17
C3794 sel_27 vss 3.13114e-17
C3795 sel_26 vss 3.13114e-17
C3796 sel_28 vss 3.13114e-17
C3797 sel_27 vss 3.13114e-17
C3798 sel_29 vss 3.13114e-17
C3799 sel_28 vss 3.13114e-17
C3800 sel_30 vss 2.42663e-16
C3801 sel_29 vss 2.42663e-16
C3802 sel_31 vss 3.13114e-17
C3803 sel_30 vss 3.13114e-17
C3804 sel_32 vss 3.13114e-17
C3805 sel_31 vss 3.13114e-17
C3806 sel_33 vss 3.13114e-17
C3807 sel_32 vss 3.13114e-17
C3808 sel_34 vss 3.13114e-17
C3809 sel_33 vss 3.13114e-17
C3810 sel_35 vss 3.13114e-17
C3811 sel_34 vss 3.13114e-17
C3812 sel_36 vss 3.13114e-17
C3813 sel_35 vss 3.13114e-17
C3814 sel_37 vss 3.13114e-17
C3815 sel_36 vss 3.13114e-17
C3816 sel_38 vss 3.13114e-17
C3817 sel_37 vss 3.13114e-17
C3818 sel_39 vss 3.13114e-17
C3819 sel_38 vss 3.13114e-17
C3820 sel_40 vss 3.13114e-17
C3821 sel_39 vss 3.13114e-17
C3822 sel_41 vss 3.13114e-17
C3823 sel_40 vss 3.13114e-17
C3824 sel_42 vss 3.13114e-17
C3825 sel_41 vss 3.13114e-17
C3826 sel_43 vss 3.13114e-17
C3827 sel_42 vss 3.13114e-17
C3828 sel_44 vss 3.13114e-17
C3829 sel_43 vss 3.13114e-17
C3830 sel_45 vss 3.13114e-17
C3831 sel_44 vss 3.13114e-17
C3832 sel_46 vss 3.13114e-17
C3833 sel_45 vss 3.13114e-17
C3834 sel_47 vss 3.13114e-17
C3835 sel_46 vss 3.13114e-17
C3836 sel_48 vss 3.13114e-17
C3837 sel_47 vss 3.13114e-17
C3838 sel_49 vss 3.13114e-17
C3839 sel_48 vss 3.13114e-17
C3840 sel_50 vss 1.40901e-17
C3841 sel_49 vss 1.40901e-17
C3842 sel_57 vss 1.40901e-16
C3843 sel_53 vss 1.40901e-16
C3844 sel_58 vss 3.13114e-17
C3845 sel_57 vss 3.13114e-17
C3846 sel_59 vss 3.13114e-17
C3847 sel_58 vss 3.13114e-17
C3848 sel_60 vss 3.13114e-17
C3849 sel_59 vss 3.13114e-17
C3850 sel_61 vss 3.13114e-17
C3851 sel_60 vss 3.13114e-17
C3852 sel_62 vss 3.13114e-17
C3853 sel_61 vss 3.13114e-17
C3854 sel_63 vss 3.13114e-17
C3855 sel_62 vss 3.13114e-17
C3856 sel_64 vss 3.13114e-17
C3857 sel_63 vss 3.13114e-17
C3858 sel_65 vss 2.42663e-16
C3859 sel_64 vss 2.42663e-16
C3860 sel_66 vss 3.13114e-17
C3861 sel_65 vss 3.13114e-17
C3862 sel_67 vss 3.13114e-17
C3863 sel_66 vss 3.13114e-17
C3864 sel_68 vss 3.13114e-17
C3865 sel_67 vss 3.13114e-17
C3866 sel_69 vss 3.13114e-17
C3867 sel_68 vss 3.13114e-17
C3868 sel_70 vss 3.13114e-17
C3869 sel_69 vss 3.13114e-17
C3870 sel_71 vss 3.13114e-17
C3871 sel_70 vss 3.13114e-17
C3872 sel_72 vss 3.13114e-17
C3873 sel_71 vss 3.13114e-17
C3874 sel_73 vss 3.13114e-17
C3875 sel_72 vss 3.13114e-17
C3876 sel_74 vss 3.13114e-17
C3877 sel_73 vss 3.13114e-17
C3878 sel_75 vss 3.13114e-17
C3879 sel_74 vss 3.13114e-17
C3880 sel_76 vss 3.13114e-17
C3881 sel_75 vss 3.13114e-17
C3882 sel_77 vss 3.13114e-17
C3883 sel_76 vss 3.13114e-17
C3884 sel_78 vss 3.13114e-17
C3885 sel_77 vss 3.13114e-17
C3886 sel_79 vss 3.13114e-17
C3887 sel_78 vss 3.13114e-17
C3888 sel_80 vss 3.13114e-17
C3889 sel_79 vss 3.13114e-17
C3890 sel_81 vss 3.13114e-17
C3891 sel_80 vss 3.13114e-17
C3892 sel_82 vss 3.13114e-17
C3893 sel_81 vss 3.13114e-17
C3894 sel_83 vss 3.13114e-17
C3895 sel_82 vss 3.13114e-17
C3896 sel_84 vss 3.13114e-17
C3897 sel_83 vss 3.13114e-17
C3898 sel_85 vss 1.40901e-17
C3899 sel_84 vss 1.40901e-17
C3900 sel_53 vss 6.34418e-17
C3901 sel_51 vss 6.34418e-17
C3902 sel_52 vss 1.42197e-16
C3903 sel_53 vss 1.42197e-16
C3904 sel_53 vss 6.8969e-16
C3905 sel_56 vss 6.8969e-16
C3906 sel vss 4.3846e-15
C3907 sel_55 vss 4.3846e-15
C3908 sel_56 vss 3.48676e-17
C3909 sel_55 vss 3.48676e-17

R63_1 bb_3_3 bb_3_6 0.001
R63_2 bb_3_7 bb_3_19 0.001
R63_3 bb_3_5 bb_3_11 0.001
R63_4 bb_3_13 bb_3_24 0.001
R63_5 bb_3_14 bb_3_12 0.001
R63_6 bb_3_22 bb_3_46 0.001
R63_7 bb_3_43 bb_3_25 0.001
R63_8 bb_3_42 bb_3_25 0.001
R63_9 bb_3_45 bb_3_25 0.001
R63_10 bb_3_44 bb_3_25 0.001
R63_11 bb_3_35 bb_3_26 0.001
R63_12 bb_3_34 bb_3_26 0.001
R63_13 bb_3_33 bb_3_26 0.001
R63_14 bb_3_28 bb_3_26 0.001
R63_15 bb_3_29 bb_3_26 0.001
R63_16 bb_3_30 bb_3_26 0.001
R63_17 bb_3_31 bb_3_26 0.001
R63_18 bb_3_32 bb_3_26 0.001
R63_19 bb_3_37 bb_3_26 0.001
R63_20 bb_3_39 bb_3_26 0.001
R63_21 bb_3_38 bb_3_26 0.001
R63_22 bb_3_40 bb_3_26 0.001
R63_23 bb_3_41 bb_3_26 0.001
R63_24 bb_3_36 bb_3_26 0.001
R63_25 bb_3_28 bb_3_27 0.001
R63_26 bb_3_29 bb_3_28 0.108
R63_27 bb_3_30 bb_3_29 0.108
R63_28 bb_3_31 bb_3_30 0.108
R63_29 bb_3_32 bb_3_31 0.108
R63_30 bb_3_33 bb_3_32 0.108
R63_31 bb_3_34 bb_3_33 0.108
R63_32 bb_3_35 bb_3_34 0.108
R63_33 bb_3_36 bb_3_35 0.108
R63_34 bb_3_37 bb_3_36 0.108
R63_35 bb_3_38 bb_3_37 0.108
R63_36 bb_3_39 bb_3_38 0.108
R63_37 bb_3_40 bb_3_39 0.108
R63_38 bb_3_41 bb_3_40 0.108
R63_39 bb_3_42 bb_3_41 0.864
R63_40 bb_3_43 bb_3_42 0.108
R63_41 bb_3_44 bb_3_43 0.108
R63_42 bb_3_45 bb_3_44 0.108
R63_43 bb_3_46 bb_3_45 0.54
R63_44 bb_3_47 bb_3_46 0.001
R63_45 bb_3_22 bb_3_21 0.001
R63_46 bb_3_23 bb_3_22 0.054
R63_47 bb_3_24 bb_3_23 5.724
R63_48 bb_3_13 bb_3_12 17.712
R63_49 bb_3_15 bb_3_14 0.648
R63_50 bb_3_10 bb_3_8 115.2
R63_51 bb_3 bb_3_10 64.8
R63_52 bb_3_16 bb_3_15 0.054
R63_53 bb_3_17 bb_3_16 0.378
R63_54 bb_3_11 bb_3_10 7.2
R63_55 bb_3_18 bb_3_17 0.054
R63_56 bb_3_19 bb_3_18 0.702
R63_57 bb_3_20 bb_3_19 0.378
R63_58 bb_3_6 bb_3_5 0.756
R63_59 bb_3_7 bb_3_6 0.108
R63_60 bb_3_4 bb_3_1 115.2
R63_61 bb_3_2 bb_3_4 43.2
R63_62 bb_3_4 bb_3_3 7.2

C3910 bb_3_28 vss 1.40901e-17
C3911 bb_3_27 vss 1.40901e-17
C3912 bb_3_29 vss 3.13114e-17
C3913 bb_3_28 vss 3.13114e-17
C3914 bb_3_30 vss 3.13114e-17
C3915 bb_3_29 vss 3.13114e-17
C3916 bb_3_31 vss 3.13114e-17
C3917 bb_3_30 vss 3.13114e-17
C3918 bb_3_32 vss 3.13114e-17
C3919 bb_3_31 vss 3.13114e-17
C3920 bb_3_33 vss 3.13114e-17
C3921 bb_3_32 vss 3.13114e-17
C3922 bb_3_34 vss 3.13114e-17
C3923 bb_3_33 vss 3.13114e-17
C3924 bb_3_35 vss 3.13114e-17
C3925 bb_3_34 vss 3.13114e-17
C3926 bb_3_36 vss 3.13114e-17
C3927 bb_3_35 vss 3.13114e-17
C3928 bb_3_37 vss 3.13114e-17
C3929 bb_3_36 vss 3.13114e-17
C3930 bb_3_38 vss 3.13114e-17
C3931 bb_3_37 vss 3.13114e-17
C3932 bb_3_39 vss 3.13114e-17
C3933 bb_3_38 vss 3.13114e-17
C3934 bb_3_40 vss 3.13114e-17
C3935 bb_3_39 vss 3.13114e-17
C3936 bb_3_41 vss 3.13114e-17
C3937 bb_3_40 vss 3.13114e-17
C3938 bb_3_42 vss 2.42663e-16
C3939 bb_3_41 vss 2.42663e-16
C3940 bb_3_43 vss 3.91392e-17
C3941 bb_3_42 vss 3.91392e-17
C3942 bb_3_44 vss 3.91392e-17
C3943 bb_3_43 vss 3.91392e-17
C3944 bb_3_45 vss 3.91392e-17
C3945 bb_3_44 vss 3.91392e-17
C3946 bb_3_46 vss 1.64385e-16
C3947 bb_3_45 vss 1.64385e-16
C3948 bb_3_47 vss 2.1918e-17
C3949 bb_3_46 vss 2.1918e-17
C3950 bb_3_22 vss 1.30248e-17
C3951 bb_3_21 vss 1.30248e-17
C3952 bb_3_23 vss 1.95372e-17
C3953 bb_3_22 vss 1.95372e-17
C3954 bb_3_24 vss 2.07745e-15
C3955 bb_3_23 vss 2.07745e-15
C3956 bb_3_13 vss 1.78604e-15
C3957 bb_3_12 vss 1.78604e-15
C3958 bb_3_15 vss 1.47744e-16
C3959 bb_3_14 vss 1.47744e-16
C3960 bb_3_10 vss 1.25194e-16
C3961 bb_3_8 vss 1.25194e-16
C3962 bb_3 vss 7.43336e-17
C3963 bb_3_10 vss 7.43336e-17
C3964 bb_3_16 vss 1.2312e-17
C3965 bb_3_15 vss 1.2312e-17
C3966 bb_3_17 vss 9.234e-17
C3967 bb_3_16 vss 9.234e-17
C3968 bb_3_11 vss 3.15414e-17
C3969 bb_3_10 vss 3.15414e-17
C3970 bb_3_18 vss 1.2312e-17
C3971 bb_3_17 vss 1.2312e-17
C3972 bb_3_19 vss 1.66212e-16
C3973 bb_3_18 vss 1.66212e-16
C3974 bb_3_20 vss 9.234e-17
C3975 bb_3_19 vss 9.234e-17
C3976 bb_3_6 vss 8.14925e-17
C3977 bb_3_5 vss 8.14925e-17
C3978 bb_3_7 vss 3.65472e-17
C3979 bb_3_6 vss 3.65472e-17
C3980 bb_3_4 vss 1.25194e-16
C3981 bb_3_1 vss 1.25194e-16
C3982 bb_3_2 vss 5.086e-17
C3983 bb_3_4 vss 5.086e-17
C3984 bb_3_4 vss 3.15414e-17
C3985 bb_3_3 vss 3.15414e-17

R64_1 n2333_1 n2333_10 0.001
R64_2 n2333_9 n2333_5 0.001
R64_3 n2333_6 n2333_3 0.001
R64_4 n2333_8 n2333_5 0.001
R64_5 n2333_3 n2333_2 115.2
R64_6 n2333 n2333_3 43.2
R64_7 n2333_6 n2333_7 0.54
R64_8 n2333_9 n2333_7 2.376
R64_9 n2333_9 n2333_8 0.216
R64_10 n2333_11 n2333_9 0.756
R64_11 n2333_11 n2333_10 0.324

C3986 n2333_3 vss 1.25194e-16
C3987 n2333_2 vss 1.25194e-16
C3988 n2333 vss 5.086e-17
C3989 n2333_3 vss 5.086e-17
C3990 n2333_6 vss 5.43283e-17
C3991 n2333_7 vss 5.43283e-17
C3992 n2333_9 vss 2.44477e-16
C3993 n2333_7 vss 2.44477e-16
C3994 n2333_9 vss 3.83746e-17
C3995 n2333_8 vss 3.83746e-17
C3996 n2333_11 vss 8.65858e-17
C3997 n2333_9 vss 8.65858e-17
C3998 n2333_11 vss 4.07462e-17
C3999 n2333_10 vss 4.07462e-17

R65_1 core_int_9_15 core_int_9_2 0.001
R65_2 core_int_9_1 core_int_9_8 0.001
R65_3 core_int_9_26 core_int_9_17 0.001
R65_4 core_int_9_10 core_int_9_3 0.001
R65_5 core_int_9_21 core_int_9_30 0.001
R65_6 core_int_9_27 core_int_9_24 0.001
R65_7 core_int_9_5 core_int_9_13 0.001
R65_8 core_int_9_11 core_int_9_9 0.001
R65_9 core_int_9_12 core_int_9_9 0.001
R65_10 core_int_9_10 core_int_9_14 0.324
R65_11 core_int_9_12 core_int_9_11 0.216
R65_12 core_int_9_13 core_int_9_12 0.216
R65_13 core_int_9_14 core_int_9_13 0.108
R65_14 core_int_9_5 core_int_9_4 0.648
R65_15 core_int_9_6 core_int_9_5 0.486
R65_16 core_int_9_7 core_int_9_6 0.054
R65_17 core_int_9_8 core_int_9_7 0.108
R65_18 core_int_9_2 core_int_9_1 3.996
R65_19 core_int_9_15 core_int_9_19 0.108
R65_20 core_int_9_17 core_int_9_16 0.81
R65_21 core_int_9_18 core_int_9_17 0.324
R65_22 core_int_9_19 core_int_9_18 0.054
R65_23 core_int_9_24 core_int_9_23 115.2
R65_24 core_int_9 core_int_9_24 64.8
R65_25 core_int_9_26 core_int_9_27 0.216
R65_26 core_int_9_27 core_int_9_28 0.216
R65_27 core_int_9_29 core_int_9_28 1.62
R65_28 core_int_9_30 core_int_9_29 0.108
R65_29 core_int_9_21 core_int_9_20 115.2
R65_30 core_int_9_22 core_int_9_21 43.2

C4000 core_int_9_10 vss 4.07462e-17
C4001 core_int_9_14 vss 4.07462e-17
C4002 core_int_9_12 vss 4.38566e-17
C4003 core_int_9_11 vss 4.38566e-17
C4004 core_int_9_13 vss 4.38566e-17
C4005 core_int_9_12 vss 4.38566e-17
C4006 core_int_9_14 vss 3.65472e-17
C4007 core_int_9_13 vss 3.65472e-17
C4008 core_int_9_5 vss 1.47744e-16
C4009 core_int_9_4 vss 1.47744e-16
C4010 core_int_9_6 vss 1.10808e-16
C4011 core_int_9_5 vss 1.10808e-16
C4012 core_int_9_7 vss 1.2312e-17
C4013 core_int_9_6 vss 1.2312e-17
C4014 core_int_9_8 vss 3.078e-17
C4015 core_int_9_7 vss 3.078e-17
C4016 core_int_9_2 vss 4.07462e-16
C4017 core_int_9_1 vss 4.07462e-16
C4018 core_int_9_15 vss 3.078e-17
C4019 core_int_9_19 vss 3.078e-17
C4020 core_int_9_17 vss 1.8468e-16
C4021 core_int_9_16 vss 1.8468e-16
C4022 core_int_9_18 vss 7.3872e-17
C4023 core_int_9_17 vss 7.3872e-17
C4024 core_int_9_19 vss 1.2312e-17
C4025 core_int_9_18 vss 1.2312e-17
C4026 core_int_9_24 vss 1.25194e-16
C4027 core_int_9_23 vss 1.25194e-16
C4028 core_int_9 vss 7.43336e-17
C4029 core_int_9_24 vss 7.43336e-17
C4030 core_int_9_26 vss 4.38566e-17
C4031 core_int_9_27 vss 4.38566e-17
C4032 core_int_9_27 vss 2.71642e-17
C4033 core_int_9_28 vss 2.71642e-17
C4034 core_int_9_29 vss 1.69776e-16
C4035 core_int_9_28 vss 1.69776e-16
C4036 core_int_9_30 vss 2.92378e-17
C4037 core_int_9_29 vss 2.92378e-17
C4038 core_int_9_21 vss 1.25194e-16
C4039 core_int_9_20 vss 1.25194e-16
C4040 core_int_9_22 vss 5.086e-17
C4041 core_int_9_21 vss 5.086e-17

R66_1 n2381_1 n2381_10 0.001
R66_2 n2381_9 n2381_5 0.001
R66_3 n2381_6 n2381_3 0.001
R66_4 n2381_8 n2381_5 0.001
R66_5 n2381_3 n2381_2 115.2
R66_6 n2381 n2381_3 43.2
R66_7 n2381_6 n2381_7 0.54
R66_8 n2381_9 n2381_7 2.376
R66_9 n2381_9 n2381_8 0.216
R66_10 n2381_11 n2381_9 0.756
R66_11 n2381_11 n2381_10 0.324

C4042 n2381_3 vss 1.25194e-16
C4043 n2381_2 vss 1.25194e-16
C4044 n2381 vss 5.086e-17
C4045 n2381_3 vss 5.086e-17
C4046 n2381_6 vss 5.43283e-17
C4047 n2381_7 vss 5.43283e-17
C4048 n2381_9 vss 2.44477e-16
C4049 n2381_7 vss 2.44477e-16
C4050 n2381_9 vss 3.83746e-17
C4051 n2381_8 vss 3.83746e-17
C4052 n2381_11 vss 8.65858e-17
C4053 n2381_9 vss 8.65858e-17
C4054 n2381_11 vss 4.07462e-17
C4055 n2381_10 vss 4.07462e-17

R67_1 n2400_8 n2400 0.001
R67_2 n2400_10 n2400_2 0.001
R67_3 n2400_4 n2400_13 0.001
R67_4 n2400_9 n2400_6 0.001
R67_5 n2400_7 n2400_6 0.001
R67_6 n2400_9 n2400_7 0.108
R67_7 n2400_8 n2400_12 0.432
R67_8 n2400_11 n2400_9 0.648
R67_9 n2400_10 n2400_11 0.432
R67_10 n2400_12 n2400_11 0.864
R67_11 n2400_13 n2400_12 0.324
R67_12 n2400_4 n2400_3 79.2
R67_13 n2400_5 n2400_4 43.2

C4056 n2400_9 vss 2.92378e-17
C4057 n2400_7 vss 2.92378e-17
C4058 n2400_8 vss 4.75373e-17
C4059 n2400_12 vss 4.75373e-17
C4060 n2400_11 vss 7.47014e-17
C4061 n2400_9 vss 7.47014e-17
C4062 n2400_10 vss 4.75373e-17
C4063 n2400_11 vss 4.75373e-17
C4064 n2400_12 vss 9.50746e-17
C4065 n2400_11 vss 9.50746e-17
C4066 n2400_13 vss 4.07462e-17
C4067 n2400_12 vss 4.07462e-17
C4068 n2400_4 vss 8.9983e-17
C4069 n2400_3 vss 8.9983e-17
C4070 n2400_5 vss 5.086e-17
C4071 n2400_4 vss 5.086e-17

R68_1 n2412_1 n2412_10 0.001
R68_2 n2412_9 n2412_5 0.001
R68_3 n2412_6 n2412_3 0.001
R68_4 n2412_8 n2412_5 0.001
R68_5 n2412_3 n2412_2 115.2
R68_6 n2412 n2412_3 43.2
R68_7 n2412_6 n2412_7 0.54
R68_8 n2412_9 n2412_7 2.376
R68_9 n2412_9 n2412_8 0.216
R68_10 n2412_11 n2412_9 0.756
R68_11 n2412_11 n2412_10 0.324

C4072 n2412_3 vss 1.25194e-16
C4073 n2412_2 vss 1.25194e-16
C4074 n2412 vss 5.086e-17
C4075 n2412_3 vss 5.086e-17
C4076 n2412_6 vss 5.43283e-17
C4077 n2412_7 vss 5.43283e-17
C4078 n2412_9 vss 2.44477e-16
C4079 n2412_7 vss 2.44477e-16
C4080 n2412_9 vss 3.83746e-17
C4081 n2412_8 vss 3.83746e-17
C4082 n2412_11 vss 8.65858e-17
C4083 n2412_9 vss 8.65858e-17
C4084 n2412_11 vss 4.07462e-17
C4085 n2412_10 vss 4.07462e-17

R69_1 n2427_6 n2427 0.001
R69_2 n2427_3 n2427_11 0.001
R69_3 n2427_7 n2427_5 0.001
R69_4 n2427_9 n2427_6 0.108
R69_5 n2427_8 n2427_7 0.108
R69_6 n2427_10 n2427_8 0.756
R69_7 n2427_9 n2427_10 0.216
R69_8 n2427_12 n2427_10 0.54
R69_9 n2427_12 n2427_11 0.108
R69_10 n2427_3 n2427_2 79.2
R69_11 n2427_4 n2427_3 43.2

C4086 n2427_9 vss 2.92378e-17
C4087 n2427_6 vss 2.92378e-17
C4088 n2427_8 vss 2.19283e-17
C4089 n2427_7 vss 2.19283e-17
C4090 n2427_10 vss 8.14925e-17
C4091 n2427_8 vss 8.14925e-17
C4092 n2427_9 vss 2.71642e-17
C4093 n2427_10 vss 2.71642e-17
C4094 n2427_12 vss 6.11194e-17
C4095 n2427_10 vss 6.11194e-17
C4096 n2427_12 vss 2.19283e-17
C4097 n2427_11 vss 2.19283e-17
C4098 n2427_3 vss 8.9983e-17
C4099 n2427_2 vss 8.9983e-17
C4100 n2427_4 vss 5.086e-17
C4101 n2427_3 vss 5.086e-17

R70_1 n2447_6 n2447 0.001
R70_2 n2447_3 n2447_11 0.001
R70_3 n2447_7 n2447_5 0.001
R70_4 n2447_9 n2447_6 0.108
R70_5 n2447_8 n2447_7 0.108
R70_6 n2447_10 n2447_8 0.756
R70_7 n2447_9 n2447_10 0.216
R70_8 n2447_12 n2447_10 0.54
R70_9 n2447_12 n2447_11 0.108
R70_10 n2447_3 n2447_2 79.2
R70_11 n2447_4 n2447_3 43.2

C4102 n2447_9 vss 2.92378e-17
C4103 n2447_6 vss 2.92378e-17
C4104 n2447_8 vss 2.19283e-17
C4105 n2447_7 vss 2.19283e-17
C4106 n2447_10 vss 8.14925e-17
C4107 n2447_8 vss 8.14925e-17
C4108 n2447_9 vss 2.71642e-17
C4109 n2447_10 vss 2.71642e-17
C4110 n2447_12 vss 6.11194e-17
C4111 n2447_10 vss 6.11194e-17
C4112 n2447_12 vss 2.19283e-17
C4113 n2447_11 vss 2.19283e-17
C4114 n2447_3 vss 8.9983e-17
C4115 n2447_2 vss 8.9983e-17
C4116 n2447_4 vss 5.086e-17
C4117 n2447_3 vss 5.086e-17

R71_1 core_int_7_13 core_int_7_2 0.001
R71_2 core_int_7_1 core_int_7_11 0.001
R71_3 core_int_7 core_int_7_22 0.001
R71_4 core_int_7_21 core_int_7_15 0.001
R71_5 core_int_7_6 core_int_7_3 0.001
R71_6 core_int_7_20 core_int_7_18 0.001
R71_7 core_int_7_19 core_int_7_18 0.001
R71_8 core_int_7_8 core_int_7_5 0.001
R71_9 core_int_7_4 core_int_7_3 136.8
R71_10 core_int_7_6 core_int_7_5 0.648
R71_11 core_int_7_8 core_int_7_7 0.324
R71_12 core_int_7_9 core_int_7_8 0.81
R71_13 core_int_7_10 core_int_7_9 0.054
R71_14 core_int_7_11 core_int_7_10 0.108
R71_15 core_int_7_2 core_int_7_1 7.236
R71_16 core_int_7_13 core_int_7_17 0.108
R71_17 core_int_7_15 core_int_7_14 0.648
R71_18 core_int_7_16 core_int_7_15 0.432
R71_19 core_int_7_17 core_int_7_16 0.054
R71_20 core_int_7_20 core_int_7_19 0.216
R71_21 core_int_7_21 core_int_7_20 0.216
R71_22 core_int_7_22 core_int_7_21 0.216

C4118 core_int_7_4 vss 1.54536e-16
C4119 core_int_7_3 vss 1.54536e-16
C4120 core_int_7_6 vss 6.62126e-17
C4121 core_int_7_5 vss 6.62126e-17
C4122 core_int_7_8 vss 7.3872e-17
C4123 core_int_7_7 vss 7.3872e-17
C4124 core_int_7_9 vss 1.8468e-16
C4125 core_int_7_8 vss 1.8468e-16
C4126 core_int_7_10 vss 1.2312e-17
C4127 core_int_7_9 vss 1.2312e-17
C4128 core_int_7_11 vss 3.078e-17
C4129 core_int_7_10 vss 3.078e-17
C4130 core_int_7_2 vss 7.33432e-16
C4131 core_int_7_1 vss 7.33432e-16
C4132 core_int_7_13 vss 3.078e-17
C4133 core_int_7_17 vss 3.078e-17
C4134 core_int_7_15 vss 1.539e-16
C4135 core_int_7_14 vss 1.539e-16
C4136 core_int_7_16 vss 1.04652e-16
C4137 core_int_7_15 vss 1.04652e-16
C4138 core_int_7_17 vss 1.2312e-17
C4139 core_int_7_16 vss 1.2312e-17
C4140 core_int_7_20 vss 4.38566e-17
C4141 core_int_7_19 vss 4.38566e-17
C4142 core_int_7_21 vss 5.11661e-17
C4143 core_int_7_20 vss 5.11661e-17
C4144 core_int_7_22 vss 5.11661e-17
C4145 core_int_7_21 vss 5.11661e-17

R72_1 n2489_8 n2489 0.001
R72_2 n2489_10 n2489_2 0.001
R72_3 n2489_4 n2489_13 0.001
R72_4 n2489_9 n2489_6 0.001
R72_5 n2489_7 n2489_6 0.001
R72_6 n2489_9 n2489_7 0.108
R72_7 n2489_8 n2489_12 0.432
R72_8 n2489_11 n2489_9 0.648
R72_9 n2489_10 n2489_11 0.432
R72_10 n2489_12 n2489_11 0.864
R72_11 n2489_13 n2489_12 0.324
R72_12 n2489_4 n2489_3 79.2
R72_13 n2489_5 n2489_4 43.2

C4146 n2489_9 vss 2.92378e-17
C4147 n2489_7 vss 2.92378e-17
C4148 n2489_8 vss 4.75373e-17
C4149 n2489_12 vss 4.75373e-17
C4150 n2489_11 vss 7.47014e-17
C4151 n2489_9 vss 7.47014e-17
C4152 n2489_10 vss 4.75373e-17
C4153 n2489_11 vss 4.75373e-17
C4154 n2489_12 vss 9.50746e-17
C4155 n2489_11 vss 9.50746e-17
C4156 n2489_13 vss 4.07462e-17
C4157 n2489_12 vss 4.07462e-17
C4158 n2489_4 vss 8.9983e-17
C4159 n2489_3 vss 8.9983e-17
C4160 n2489_5 vss 5.086e-17
C4161 n2489_4 vss 5.086e-17

R73_1 n2503_6 n2503 0.001
R73_2 n2503_3 n2503_11 0.001
R73_3 n2503_7 n2503_5 0.001
R73_4 n2503_9 n2503_6 0.108
R73_5 n2503_8 n2503_7 0.108
R73_6 n2503_10 n2503_8 0.756
R73_7 n2503_9 n2503_10 0.216
R73_8 n2503_12 n2503_10 0.54
R73_9 n2503_12 n2503_11 0.108
R73_10 n2503_3 n2503_2 79.2
R73_11 n2503_4 n2503_3 43.2

C4162 n2503_9 vss 2.92378e-17
C4163 n2503_6 vss 2.92378e-17
C4164 n2503_8 vss 2.19283e-17
C4165 n2503_7 vss 2.19283e-17
C4166 n2503_10 vss 8.14925e-17
C4167 n2503_8 vss 8.14925e-17
C4168 n2503_9 vss 2.71642e-17
C4169 n2503_10 vss 2.71642e-17
C4170 n2503_12 vss 6.11194e-17
C4171 n2503_10 vss 6.11194e-17
C4172 n2503_12 vss 2.19283e-17
C4173 n2503_11 vss 2.19283e-17
C4174 n2503_3 vss 8.9983e-17
C4175 n2503_2 vss 8.9983e-17
C4176 n2503_4 vss 5.086e-17
C4177 n2503_3 vss 5.086e-17

R74_1 n2517 n2517_11 0.001
R74_2 n2517_6 n2517_3 0.001
R74_3 n2517_8 n2517_5 0.001
R74_4 n2517_3 n2517_2 79.2
R74_5 n2517_4 n2517_3 43.2
R74_6 n2517_7 n2517_6 0.108
R74_7 n2517_7 n2517_10 0.54
R74_8 n2517_9 n2517_8 0.108
R74_9 n2517_10 n2517_9 0.756
R74_10 n2517_12 n2517_10 0.216
R74_11 n2517_12 n2517_11 0.108

C4178 n2517_3 vss 8.9983e-17
C4179 n2517_2 vss 8.9983e-17
C4180 n2517_4 vss 5.086e-17
C4181 n2517_3 vss 5.086e-17
C4182 n2517_7 vss 2.19283e-17
C4183 n2517_6 vss 2.19283e-17
C4184 n2517_7 vss 6.11194e-17
C4185 n2517_10 vss 6.11194e-17
C4186 n2517_9 vss 2.19283e-17
C4187 n2517_8 vss 2.19283e-17
C4188 n2517_10 vss 8.14925e-17
C4189 n2517_9 vss 8.14925e-17
C4190 n2517_12 vss 2.71642e-17
C4191 n2517_10 vss 2.71642e-17
C4192 n2517_12 vss 2.92378e-17
C4193 n2517_11 vss 2.92378e-17

R75_1 core_int_3_13 core_int_3_2 0.001
R75_2 core_int_3_1 core_int_3_11 0.001
R75_3 core_int_3 core_int_3_22 0.001
R75_4 core_int_3_21 core_int_3_15 0.001
R75_5 core_int_3_6 core_int_3_3 0.001
R75_6 core_int_3_19 core_int_3_18 0.001
R75_7 core_int_3_20 core_int_3_18 0.001
R75_8 core_int_3_8 core_int_3_5 0.001
R75_9 core_int_3_4 core_int_3_3 136.8
R75_10 core_int_3_6 core_int_3_5 0.648
R75_11 core_int_3_8 core_int_3_7 0.324
R75_12 core_int_3_9 core_int_3_8 0.81
R75_13 core_int_3_10 core_int_3_9 0.054
R75_14 core_int_3_11 core_int_3_10 0.108
R75_15 core_int_3_2 core_int_3_1 6.48
R75_16 core_int_3_13 core_int_3_17 0.108
R75_17 core_int_3_15 core_int_3_14 0.648
R75_18 core_int_3_16 core_int_3_15 0.432
R75_19 core_int_3_17 core_int_3_16 0.054
R75_20 core_int_3_20 core_int_3_19 0.216
R75_21 core_int_3_21 core_int_3_20 0.216
R75_22 core_int_3_22 core_int_3_21 0.216

C4194 core_int_3_4 vss 1.54536e-16
C4195 core_int_3_3 vss 1.54536e-16
C4196 core_int_3_6 vss 6.62126e-17
C4197 core_int_3_5 vss 6.62126e-17
C4198 core_int_3_8 vss 7.3872e-17
C4199 core_int_3_7 vss 7.3872e-17
C4200 core_int_3_9 vss 1.8468e-16
C4201 core_int_3_8 vss 1.8468e-16
C4202 core_int_3_10 vss 1.2312e-17
C4203 core_int_3_9 vss 1.2312e-17
C4204 core_int_3_11 vss 3.078e-17
C4205 core_int_3_10 vss 3.078e-17
C4206 core_int_3_2 vss 6.5194e-16
C4207 core_int_3_1 vss 6.5194e-16
C4208 core_int_3_13 vss 3.078e-17
C4209 core_int_3_17 vss 3.078e-17
C4210 core_int_3_15 vss 1.539e-16
C4211 core_int_3_14 vss 1.539e-16
C4212 core_int_3_16 vss 1.04652e-16
C4213 core_int_3_15 vss 1.04652e-16
C4214 core_int_3_17 vss 1.2312e-17
C4215 core_int_3_16 vss 1.2312e-17
C4216 core_int_3_20 vss 4.38566e-17
C4217 core_int_3_19 vss 4.38566e-17
C4218 core_int_3_21 vss 5.11661e-17
C4219 core_int_3_20 vss 5.11661e-17
C4220 core_int_3_22 vss 5.11661e-17
C4221 core_int_3_21 vss 5.11661e-17

R76_1 n2561 n2561_10 0.001
R76_2 n2561_7 n2561_4 0.001
R76_3 n2561_6 n2561_5 0.001
R76_4 n2561_2 n2561_4 144
R76_5 n2561_4 n2561_3 72
R76_6 n2561_7 n2561_6 0.216
R76_7 n2561_7 n2561_8 0.54
R76_8 n2561_9 n2561_8 0.648
R76_9 n2561_10 n2561_9 0.432

C4222 n2561_2 vss 1.6236e-16
C4223 n2561_4 vss 1.6236e-16
C4224 n2561_4 vss 7.8246e-17
C4225 n2561_3 vss 7.8246e-17
C4226 n2561_7 vss 3.22574e-17
C4227 n2561_6 vss 3.22574e-17
C4228 n2561_7 vss 5.60261e-17
C4229 n2561_8 vss 5.60261e-17
C4230 n2561_9 vss 7.47014e-17
C4231 n2561_8 vss 7.47014e-17
C4232 n2561_10 vss 4.75373e-17
C4233 n2561_9 vss 4.75373e-17

R77_1 n2566 n2566_5 0.001
R77_2 n2566_3 n2566_2 0.001
R77_3 n2566_4 n2566_2 0.001
R77_4 n2566_4 n2566_3 0.108
R77_5 n2566_5 n2566_4 1.08

C4234 n2566_4 vss 3.10651e-17
C4235 n2566_3 vss 3.10651e-17
C4236 n2566_5 vss 1.18843e-16
C4237 n2566_4 vss 1.18843e-16

R78_1 core_l2_dff_s_1 core_l2_dff_s_6 0.001
R78_2 core_l2_dff_s_3 core_l2_dff_s_12 0.001
R78_3 core_l2_dff_s_4 core_l2_dff_s_2 0.001
R78_4 core_l2_dff_s core_l2_dff_s_9 180
R78_5 core_l2_dff_s_11 core_l2_dff_s_8 50.4
R78_6 core_l2_dff_s_11 core_l2_dff_s_9 43.2
R78_7 core_l2_dff_s_10 core_l2_dff_s_12 43.2
R78_8 core_l2_dff_s_12 core_l2_dff_s_11 28.8
R78_9 core_l2_dff_s_5 core_l2_dff_s_3 0.54
R78_10 core_l2_dff_s_5 core_l2_dff_s_4 0.648
R78_11 core_l2_dff_s_6 core_l2_dff_s_5 0.54

C4238 core_l2_dff_s vss 1.97571e-16
C4239 core_l2_dff_s_9 vss 1.97571e-16
C4240 core_l2_dff_s_11 vss 5.47722e-17
C4241 core_l2_dff_s_8 vss 5.47722e-17
C4242 core_l2_dff_s_11 vss 4.69476e-17
C4243 core_l2_dff_s_9 vss 4.69476e-17
C4244 core_l2_dff_s_10 vss 4.69476e-17
C4245 core_l2_dff_s_12 vss 4.69476e-17
C4246 core_l2_dff_s_12 vss 3.12984e-17
C4247 core_l2_dff_s_11 vss 3.12984e-17
C4248 core_l2_dff_s_5 vss 5.43283e-17
C4249 core_l2_dff_s_3 vss 5.43283e-17
C4250 core_l2_dff_s_5 vss 7.47014e-17
C4251 core_l2_dff_s_4 vss 7.47014e-17
C4252 core_l2_dff_s_6 vss 5.43283e-17
C4253 core_l2_dff_s_5 vss 5.43283e-17

R79_1 n2593 n2593_12 0.001
R79_2 n2593_10 n2593_5 0.001
R79_3 n2593_8 n2593_6 0.001
R79_4 n2593_7 n2593_6 0.001
R79_5 n2593_2 n2593_3 72
R79_6 n2593_8 n2593_7 0.108
R79_7 n2593_4 n2593_3 64.8
R79_8 n2593_8 n2593_9 0.324
R79_9 n2593_5 n2593_4 21.6
R79_10 n2593_10 n2593_9 0.648
R79_11 n2593_11 n2593_10 0.324
R79_12 n2593_12 n2593_11 0.324

C4254 n2593_2 vss 8.21582e-17
C4255 n2593_3 vss 8.21582e-17
C4256 n2593_8 vss 3.10651e-17
C4257 n2593_7 vss 3.10651e-17
C4258 n2593_4 vss 7.04214e-17
C4259 n2593_3 vss 7.04214e-17
C4260 n2593_8 vss 4.07462e-17
C4261 n2593_9 vss 4.07462e-17
C4262 n2593_5 vss 2.34738e-17
C4263 n2593_4 vss 2.34738e-17
C4264 n2593_10 vss 7.47014e-17
C4265 n2593_9 vss 7.47014e-17
C4266 n2593_11 vss 3.39552e-17
C4267 n2593_10 vss 3.39552e-17
C4268 n2593_12 vss 4.07462e-17
C4269 n2593_11 vss 4.07462e-17

R80_1 core_l2_dff_m core_l2_dff_m_12 0.001
R80_2 core_l2_dff_m_7 core_l2_dff_m_2 0.001
R80_3 core_l2_dff_m_6 core_l2_dff_m_4 0.001
R80_4 core_l2_dff_m_4 core_l2_dff_m_3 64.8
R80_5 core_l2_dff_m_5 core_l2_dff_m_4 93.6
R80_6 core_l2_dff_m_8 core_l2_dff_m_6 0.648
R80_7 core_l2_dff_m_8 core_l2_dff_m_7 0.216
R80_8 core_l2_dff_m_9 core_l2_dff_m_8 0.108
R80_9 core_l2_dff_m_10 core_l2_dff_m_9 0.648
R80_10 core_l2_dff_m_10 core_l2_dff_m_11 0.108
R80_11 core_l2_dff_m_12 core_l2_dff_m_11 0.216

C4270 core_l2_dff_m_4 vss 7.04214e-17
C4271 core_l2_dff_m_3 vss 7.04214e-17
C4272 core_l2_dff_m_5 vss 1.0172e-16
C4273 core_l2_dff_m_4 vss 1.0172e-16
C4274 core_l2_dff_m_8 vss 6.79104e-17
C4275 core_l2_dff_m_6 vss 6.79104e-17
C4276 core_l2_dff_m_8 vss 2.71642e-17
C4277 core_l2_dff_m_7 vss 2.71642e-17
C4278 core_l2_dff_m_9 vss 1.35821e-17
C4279 core_l2_dff_m_8 vss 1.35821e-17
C4280 core_l2_dff_m_10 vss 6.79104e-17
C4281 core_l2_dff_m_9 vss 6.79104e-17
C4282 core_l2_dff_m_10 vss 1.35821e-17
C4283 core_l2_dff_m_11 vss 1.35821e-17
C4284 core_l2_dff_m_12 vss 2.71642e-17
C4285 core_l2_dff_m_11 vss 2.71642e-17

R81_1 n2624 n2624_18 0.001
R81_2 n2624_17 n2624_7 0.001
R81_3 n2624_12 n2624_9 0.001
R81_4 n2624_15 n2624_14 0.001
R81_5 n2624_13 n2624_11 0.001
R81_6 n2624_6 n2624_4 0.001
R81_7 n2624_3 n2624_2 0.001
R81_8 n2624_10 n2624_9 43.2
R81_9 n2624_12 n2624_11 0.54
R81_10 n2624_6 n2624_5 36
R81_11 n2624_4 n2624_3 0.108
R81_12 n2624_14 n2624_13 57.6
R81_13 n2624_7 n2624_6 93.6
R81_14 n2624_16 n2624_15 0.54
R81_15 n2624_8 n2624_7 86.4
R81_16 n2624_17 n2624_16 0.972
R81_17 n2624_18 n2624_17 0.216

C4286 n2624_10 vss 5.086e-17
C4287 n2624_9 vss 5.086e-17
C4288 n2624_12 vss 5.43283e-17
C4289 n2624_11 vss 5.43283e-17
C4290 n2624_6 vss 3.9123e-17
C4291 n2624_5 vss 3.9123e-17
C4292 n2624_4 vss 2.92378e-17
C4293 n2624_3 vss 2.92378e-17
C4294 n2624_14 vss 6.25968e-17
C4295 n2624_13 vss 6.25968e-17
C4296 n2624_7 vss 1.0172e-16
C4297 n2624_6 vss 1.0172e-16
C4298 n2624_16 vss 5.43283e-17
C4299 n2624_15 vss 5.43283e-17
C4300 n2624_8 vss 9.97636e-17
C4301 n2624_7 vss 9.97636e-17
C4302 n2624_17 vss 1.00168e-16
C4303 n2624_16 vss 1.00168e-16
C4304 n2624_18 vss 2.71642e-17
C4305 n2624_17 vss 2.71642e-17

R82_1 n2635 n2635_5 0.001
R82_2 n2635_4 n2635_2 0.001
R82_3 n2635_3 n2635_2 0.001
R82_4 n2635_4 n2635_3 0.108
R82_5 n2635_5 n2635_4 1.188

C4306 n2635_4 vss 2.92378e-17
C4307 n2635_3 vss 2.92378e-17
C4308 n2635_5 vss 1.22239e-16
C4309 n2635_4 vss 1.22239e-16

R83_1 n2646 n2646_11 0.001
R83_2 n2646_6 n2646_3 0.001
R83_3 n2646_8 n2646_5 0.001
R83_4 n2646_3 n2646_2 79.2
R83_5 n2646_4 n2646_3 43.2
R83_6 n2646_7 n2646_6 0.108
R83_7 n2646_7 n2646_10 0.54
R83_8 n2646_9 n2646_8 0.108
R83_9 n2646_10 n2646_9 0.756
R83_10 n2646_12 n2646_10 0.216
R83_11 n2646_12 n2646_11 0.108

C4310 n2646_3 vss 8.9983e-17
C4311 n2646_2 vss 8.9983e-17
C4312 n2646_4 vss 5.086e-17
C4313 n2646_3 vss 5.086e-17
C4314 n2646_7 vss 2.19283e-17
C4315 n2646_6 vss 2.19283e-17
C4316 n2646_7 vss 6.11194e-17
C4317 n2646_10 vss 6.11194e-17
C4318 n2646_9 vss 2.19283e-17
C4319 n2646_8 vss 2.19283e-17
C4320 n2646_10 vss 8.14925e-17
C4321 n2646_9 vss 8.14925e-17
C4322 n2646_12 vss 2.71642e-17
C4323 n2646_10 vss 2.71642e-17
C4324 n2646_12 vss 2.92378e-17
C4325 n2646_11 vss 2.92378e-17

R84_1 bb_0_3 bb_0_6 0.001
R84_2 bb_0_7 bb_0_25 0.001
R84_3 bb_0_5 bb_0_11 0.001
R84_4 bb_0_31 bb_0_17 0.001
R84_5 bb_0_15 bb_0_13 0.001
R84_6 bb_0_19 bb_0_41 0.001
R84_7 bb_0_30 bb_0_20 0.001
R84_8 bb_0_21 bb_0_18 0.001
R84_9 bb_0_22 bb_0_28 0.001
R84_10 bb_0_27 bb_0_36 0.001
R84_11 bb_0_33 bb_0_29 0.001
R84_12 bb_0_58 bb_0_39 0.001
R84_13 bb_0_57 bb_0_39 0.001
R84_14 bb_0_55 bb_0_39 0.001
R84_15 bb_0_56 bb_0_39 0.001
R84_16 bb_0_62 bb_0_39 0.001
R84_17 bb_0_59 bb_0_39 0.001
R84_18 bb_0_60 bb_0_39 0.001
R84_19 bb_0_61 bb_0_39 0.001
R84_20 bb_0_66 bb_0_39 0.001
R84_21 bb_0_65 bb_0_39 0.001
R84_22 bb_0_64 bb_0_39 0.001
R84_23 bb_0_63 bb_0_39 0.001
R84_24 bb_0_51 bb_0_42 0.001
R84_25 bb_0_50 bb_0_42 0.001
R84_26 bb_0_52 bb_0_42 0.001
R84_27 bb_0_54 bb_0_39 0.001
R84_28 bb_0_53 bb_0_39 0.001
R84_29 bb_0_40 bb_0_46 0.001
R84_30 bb_0_49 bb_0_42 0.001
R84_31 bb_0_48 bb_0_44 0.001
R84_32 bb_0_44 bb_0_43 0.054
R84_33 bb_0_45 bb_0_44 0.001
R84_34 bb_0_49 bb_0_48 0.54
R84_35 bb_0_50 bb_0_49 0.108
R84_36 bb_0_51 bb_0_50 0.108
R84_37 bb_0_52 bb_0_51 0.108
R84_38 bb_0_53 bb_0_52 0.864
R84_39 bb_0_54 bb_0_53 0.108
R84_40 bb_0_55 bb_0_54 0.108
R84_41 bb_0_56 bb_0_55 0.108
R84_42 bb_0_57 bb_0_56 0.108
R84_43 bb_0_58 bb_0_57 0.108
R84_44 bb_0_59 bb_0_58 0.108
R84_45 bb_0_60 bb_0_59 0.108
R84_46 bb_0_61 bb_0_60 0.108
R84_47 bb_0_62 bb_0_61 0.108
R84_48 bb_0_63 bb_0_62 0.108
R84_49 bb_0_64 bb_0_63 0.108
R84_50 bb_0_65 bb_0_64 0.108
R84_51 bb_0_66 bb_0_65 0.108
R84_52 bb_0_67 bb_0_66 0.001
R84_53 bb_0_47 bb_0_46 0.54
R84_54 bb_0_48 bb_0_47 0.001
R84_55 bb_0_41 bb_0_40 7.02
R84_56 bb_0_13 bb_0_12 72
R84_57 bb_0_14 bb_0_13 50.4
R84_58 bb_0_19 bb_0_18 10.044
R84_59 bb_0_15 bb_0_16 0.216
R84_60 bb_0_21 bb_0_20 0.378
R84_61 bb_0_17 bb_0_16 0.216
R84_62 bb_0_30 bb_0_29 9.288
R84_63 bb_0_31 bb_0_38 0.432
R84_64 bb_0_32 bb_0_31 0.702
R84_65 bb_0_34 bb_0_33 0.216
R84_66 bb_0_35 bb_0_34 0.054
R84_67 bb_0_36 bb_0_35 0.108
R84_68 bb_0_37 bb_0_36 0.27
R84_69 bb_0_38 bb_0_37 0.054
R84_70 bb_0_28 bb_0_27 2.808
R84_71 bb_0_10 bb_0_8 115.2
R84_72 bb_0 bb_0_10 64.8
R84_73 bb_0_23 bb_0_22 0.27
R84_74 bb_0_11 bb_0_10 7.2
R84_75 bb_0_24 bb_0_23 0.054
R84_76 bb_0_25 bb_0_24 0.702
R84_77 bb_0_26 bb_0_25 0.378
R84_78 bb_0_6 bb_0_5 0.756
R84_79 bb_0_7 bb_0_6 0.108
R84_80 bb_0_4 bb_0_1 115.2
R84_81 bb_0_2 bb_0_4 43.2
R84_82 bb_0_4 bb_0_3 7.2

C4326 bb_0_44 vss 1.95372e-17
C4327 bb_0_43 vss 1.95372e-17
C4328 bb_0_45 vss 1.30248e-17
C4329 bb_0_44 vss 1.30248e-17
C4330 bb_0_49 vss 1.64385e-16
C4331 bb_0_48 vss 1.64385e-16
C4332 bb_0_50 vss 3.91392e-17
C4333 bb_0_49 vss 3.91392e-17
C4334 bb_0_51 vss 3.91392e-17
C4335 bb_0_50 vss 3.91392e-17
C4336 bb_0_52 vss 3.91392e-17
C4337 bb_0_51 vss 3.91392e-17
C4338 bb_0_53 vss 2.42663e-16
C4339 bb_0_52 vss 2.42663e-16
C4340 bb_0_54 vss 3.13114e-17
C4341 bb_0_53 vss 3.13114e-17
C4342 bb_0_55 vss 3.13114e-17
C4343 bb_0_54 vss 3.13114e-17
C4344 bb_0_56 vss 3.13114e-17
C4345 bb_0_55 vss 3.13114e-17
C4346 bb_0_57 vss 3.13114e-17
C4347 bb_0_56 vss 3.13114e-17
C4348 bb_0_58 vss 3.13114e-17
C4349 bb_0_57 vss 3.13114e-17
C4350 bb_0_59 vss 3.13114e-17
C4351 bb_0_58 vss 3.13114e-17
C4352 bb_0_60 vss 3.13114e-17
C4353 bb_0_59 vss 3.13114e-17
C4354 bb_0_61 vss 3.13114e-17
C4355 bb_0_60 vss 3.13114e-17
C4356 bb_0_62 vss 3.13114e-17
C4357 bb_0_61 vss 3.13114e-17
C4358 bb_0_63 vss 3.13114e-17
C4359 bb_0_62 vss 3.13114e-17
C4360 bb_0_64 vss 3.13114e-17
C4361 bb_0_63 vss 3.13114e-17
C4362 bb_0_65 vss 3.13114e-17
C4363 bb_0_64 vss 3.13114e-17
C4364 bb_0_66 vss 3.13114e-17
C4365 bb_0_65 vss 3.13114e-17
C4366 bb_0_67 vss 1.40901e-17
C4367 bb_0_66 vss 1.40901e-17
C4368 bb_0_47 vss 6.24776e-17
C4369 bb_0_46 vss 6.24776e-17
C4370 bb_0_48 vss 2.1918e-17
C4371 bb_0_47 vss 2.1918e-17
C4372 bb_0_41 vss 1.60056e-15
C4373 bb_0_40 vss 1.60056e-15
C4374 bb_0_13 vss 8.21582e-17
C4375 bb_0_12 vss 8.21582e-17
C4376 bb_0_14 vss 5.86844e-17
C4377 bb_0_13 vss 5.86844e-17
C4378 bb_0_19 vss 1.01866e-15
C4379 bb_0_18 vss 1.01866e-15
C4380 bb_0_15 vss 2.71642e-17
C4381 bb_0_16 vss 2.71642e-17
C4382 bb_0_21 vss 9.234e-17
C4383 bb_0_20 vss 9.234e-17
C4384 bb_0_17 vss 2.54664e-17
C4385 bb_0_16 vss 2.54664e-17
C4386 bb_0_30 vss 9.43955e-16
C4387 bb_0_29 vss 9.43955e-16
C4388 bb_0_31 vss 9.8496e-17
C4389 bb_0_38 vss 9.8496e-17
C4390 bb_0_32 vss 1.60056e-16
C4391 bb_0_31 vss 1.60056e-16
C4392 bb_0_34 vss 5.5404e-17
C4393 bb_0_33 vss 5.5404e-17
C4394 bb_0_35 vss 1.2312e-17
C4395 bb_0_34 vss 1.2312e-17
C4396 bb_0_36 vss 3.078e-17
C4397 bb_0_35 vss 3.078e-17
C4398 bb_0_37 vss 6.156e-17
C4399 bb_0_36 vss 6.156e-17
C4400 bb_0_38 vss 1.2312e-17
C4401 bb_0_37 vss 1.2312e-17
C4402 bb_0_28 vss 2.85224e-16
C4403 bb_0_27 vss 2.85224e-16
C4404 bb_0_10 vss 1.25194e-16
C4405 bb_0_8 vss 1.25194e-16
C4406 bb_0 vss 7.43336e-17
C4407 bb_0_10 vss 7.43336e-17
C4408 bb_0_23 vss 6.156e-17
C4409 bb_0_22 vss 6.156e-17
C4410 bb_0_11 vss 3.15414e-17
C4411 bb_0_10 vss 3.15414e-17
C4412 bb_0_24 vss 1.2312e-17
C4413 bb_0_23 vss 1.2312e-17
C4414 bb_0_25 vss 1.66212e-16
C4415 bb_0_24 vss 1.66212e-16
C4416 bb_0_26 vss 9.234e-17
C4417 bb_0_25 vss 9.234e-17
C4418 bb_0_6 vss 8.14925e-17
C4419 bb_0_5 vss 8.14925e-17
C4420 bb_0_7 vss 3.65472e-17
C4421 bb_0_6 vss 3.65472e-17
C4422 bb_0_4 vss 1.25194e-16
C4423 bb_0_1 vss 1.25194e-16
C4424 bb_0_2 vss 5.086e-17
C4425 bb_0_4 vss 5.086e-17
C4426 bb_0_4 vss 3.15414e-17
C4427 bb_0_3 vss 3.15414e-17

R85_1 n2733_1 n2733_10 0.001
R85_2 n2733_9 n2733_5 0.001
R85_3 n2733_6 n2733_3 0.001
R85_4 n2733_8 n2733_5 0.001
R85_5 n2733_3 n2733_2 115.2
R85_6 n2733 n2733_3 43.2
R85_7 n2733_6 n2733_7 0.54
R85_8 n2733_9 n2733_7 2.376
R85_9 n2733_9 n2733_8 0.216
R85_10 n2733_11 n2733_9 0.756
R85_11 n2733_11 n2733_10 0.324

C4428 n2733_3 vss 1.25194e-16
C4429 n2733_2 vss 1.25194e-16
C4430 n2733 vss 5.086e-17
C4431 n2733_3 vss 5.086e-17
C4432 n2733_6 vss 5.43283e-17
C4433 n2733_7 vss 5.43283e-17
C4434 n2733_9 vss 2.44477e-16
C4435 n2733_7 vss 2.44477e-16
C4436 n2733_9 vss 3.83746e-17
C4437 n2733_8 vss 3.83746e-17
C4438 n2733_11 vss 8.65858e-17
C4439 n2733_9 vss 8.65858e-17
C4440 n2733_11 vss 4.07462e-17
C4441 n2733_10 vss 4.07462e-17

R86_1 n2750 n2750_12 0.001
R86_2 n2750_10 n2750_5 0.001
R86_3 n2750_8 n2750_6 0.001
R86_4 n2750_7 n2750_6 0.001
R86_5 n2750_2 n2750_3 72
R86_6 n2750_8 n2750_7 0.108
R86_7 n2750_4 n2750_3 64.8
R86_8 n2750_8 n2750_9 0.324
R86_9 n2750_5 n2750_4 21.6
R86_10 n2750_10 n2750_9 0.648
R86_11 n2750_11 n2750_10 0.324
R86_12 n2750_12 n2750_11 0.324

C4442 n2750_2 vss 8.21582e-17
C4443 n2750_3 vss 8.21582e-17
C4444 n2750_8 vss 3.10651e-17
C4445 n2750_7 vss 3.10651e-17
C4446 n2750_4 vss 7.04214e-17
C4447 n2750_3 vss 7.04214e-17
C4448 n2750_8 vss 4.07462e-17
C4449 n2750_9 vss 4.07462e-17
C4450 n2750_5 vss 2.34738e-17
C4451 n2750_4 vss 2.34738e-17
C4452 n2750_10 vss 7.47014e-17
C4453 n2750_9 vss 7.47014e-17
C4454 n2750_11 vss 3.39552e-17
C4455 n2750_10 vss 3.39552e-17
C4456 n2750_12 vss 4.07462e-17
C4457 n2750_11 vss 4.07462e-17

R87_1 n2765 n2765_10 0.001
R87_2 n2765_7 n2765_3 0.001
R87_3 n2765_6 n2765_5 0.001
R87_4 n2765_3 n2765_2 72
R87_5 n2765_4 n2765_3 144
R87_6 n2765_7 n2765_6 0.216
R87_7 n2765_7 n2765_8 0.54
R87_8 n2765_9 n2765_8 0.648
R87_9 n2765_10 n2765_9 0.432

C4458 n2765_3 vss 7.8246e-17
C4459 n2765_2 vss 7.8246e-17
C4460 n2765_4 vss 1.6236e-16
C4461 n2765_3 vss 1.6236e-16
C4462 n2765_7 vss 3.22574e-17
C4463 n2765_6 vss 3.22574e-17
C4464 n2765_7 vss 5.60261e-17
C4465 n2765_8 vss 5.60261e-17
C4466 n2765_9 vss 7.47014e-17
C4467 n2765_8 vss 7.47014e-17
C4468 n2765_10 vss 4.75373e-17
C4469 n2765_9 vss 4.75373e-17

R88_1 n2770 n2770_5 0.001
R88_2 n2770_4 n2770_2 0.001
R88_3 n2770_3 n2770_2 0.001
R88_4 n2770_4 n2770_3 0.108
R88_5 n2770_5 n2770_4 1.08

C4470 n2770_4 vss 3.10651e-17
C4471 n2770_3 vss 3.10651e-17
C4472 n2770_5 vss 1.18843e-16
C4473 n2770_4 vss 1.18843e-16

R89_1 core_l0_dff_s_1 core_l0_dff_s_6 0.001
R89_2 core_l0_dff_s_3 core_l0_dff_s_12 0.001
R89_3 core_l0_dff_s_4 core_l0_dff_s_2 0.001
R89_4 core_l0_dff_s core_l0_dff_s_9 180
R89_5 core_l0_dff_s_11 core_l0_dff_s_8 50.4
R89_6 core_l0_dff_s_11 core_l0_dff_s_9 43.2
R89_7 core_l0_dff_s_10 core_l0_dff_s_12 43.2
R89_8 core_l0_dff_s_12 core_l0_dff_s_11 28.8
R89_9 core_l0_dff_s_5 core_l0_dff_s_3 0.54
R89_10 core_l0_dff_s_5 core_l0_dff_s_4 0.648
R89_11 core_l0_dff_s_6 core_l0_dff_s_5 0.54

C4474 core_l0_dff_s vss 1.97571e-16
C4475 core_l0_dff_s_9 vss 1.97571e-16
C4476 core_l0_dff_s_11 vss 5.47722e-17
C4477 core_l0_dff_s_8 vss 5.47722e-17
C4478 core_l0_dff_s_11 vss 4.69476e-17
C4479 core_l0_dff_s_9 vss 4.69476e-17
C4480 core_l0_dff_s_10 vss 4.69476e-17
C4481 core_l0_dff_s_12 vss 4.69476e-17
C4482 core_l0_dff_s_12 vss 3.12984e-17
C4483 core_l0_dff_s_11 vss 3.12984e-17
C4484 core_l0_dff_s_5 vss 5.43283e-17
C4485 core_l0_dff_s_3 vss 5.43283e-17
C4486 core_l0_dff_s_5 vss 7.47014e-17
C4487 core_l0_dff_s_4 vss 7.47014e-17
C4488 core_l0_dff_s_6 vss 5.43283e-17
C4489 core_l0_dff_s_5 vss 5.43283e-17

R90_1 ss_0_2 ss_0_5 0.001
R90_2 ss_0_4 ss_0_34 0.001
R90_3 ss_0_31 ss_0_7 0.001
R90_4 ss_0_28 ss_0_21 0.001
R90_5 ss_0_6 ss_0_10 0.001
R90_6 ss_0_8 ss_0_18 0.001
R90_7 ss_0_16 ss_0_13 0.001
R90_8 ss_0_17 ss_0_13 0.001
R90_9 ss_0_15 ss_0_14 0.001
R90_10 ss_0_20 ss_0_23 0.001
R90_11 ss_0_22 ss_0_27 0.001
R90_12 ss_0_26 ss_0_25 0.001
R90_13 ss_0_25 ss_0_24 475.2
R90_14 ss_0_15 ss_0_19 0.324
R90_15 ss_0_17 ss_0_16 0.216
R90_16 ss_0_18 ss_0_17 0.216
R90_17 ss_0_19 ss_0_18 0.108
R90_18 ss_0_27 ss_0_26 0.324
R90_19 ss_0_8 ss_0_12 0.594
R90_20 ss_0_9 ss_0_8 0.54
R90_21 ss_0_23 ss_0_22 5.94
R90_22 ss_0_11 ss_0_10 0.108
R90_23 ss_0_12 ss_0_11 0.054
R90_24 ss_0_21 ss_0_20 26.244
R90_25 ss_0_7 ss_0_6 7.668
R90_26 ss_0_29 ss_0_28 0.378
R90_27 ss_0_30 ss_0_29 0.054
R90_28 ss_0_31 ss_0_30 0.27
R90_29 ss_0_32 ss_0_31 0.108
R90_30 ss_0_33 ss_0_32 0.054
R90_31 ss_0_34 ss_0_33 0.54
R90_32 ss_0_35 ss_0_34 0.54
R90_33 ss_0_5 ss_0_4 0.216
R90_34 ss_0_2 ss_0_1 108
R90_35 ss_0 ss_0_2 50.4

C4490 ss_0_25 vss 5.18379e-16
C4491 ss_0_24 vss 5.18379e-16
C4492 ss_0_15 vss 4.07462e-17
C4493 ss_0_19 vss 4.07462e-17
C4494 ss_0_17 vss 4.38566e-17
C4495 ss_0_16 vss 4.38566e-17
C4496 ss_0_18 vss 4.38566e-17
C4497 ss_0_17 vss 4.38566e-17
C4498 ss_0_19 vss 3.65472e-17
C4499 ss_0_18 vss 3.65472e-17
C4500 ss_0_27 vss 7.30944e-17
C4501 ss_0_26 vss 7.30944e-17
C4502 ss_0_8 vss 1.35432e-16
C4503 ss_0_12 vss 1.35432e-16
C4504 ss_0_9 vss 1.2312e-16
C4505 ss_0_8 vss 1.2312e-16
C4506 ss_0_23 vss 2.14909e-15
C4507 ss_0_22 vss 2.14909e-15
C4508 ss_0_11 vss 3.078e-17
C4509 ss_0_10 vss 3.078e-17
C4510 ss_0_12 vss 1.2312e-17
C4511 ss_0_11 vss 1.2312e-17
C4512 ss_0_21 vss 2.64851e-15
C4513 ss_0_20 vss 2.64851e-15
C4514 ss_0_7 vss 7.74179e-16
C4515 ss_0_6 vss 7.74179e-16
C4516 ss_0_29 vss 8.6184e-17
C4517 ss_0_28 vss 8.6184e-17
C4518 ss_0_30 vss 1.2312e-17
C4519 ss_0_29 vss 1.2312e-17
C4520 ss_0_31 vss 6.156e-17
C4521 ss_0_30 vss 6.156e-17
C4522 ss_0_32 vss 3.078e-17
C4523 ss_0_31 vss 3.078e-17
C4524 ss_0_33 vss 1.2312e-17
C4525 ss_0_32 vss 1.2312e-17
C4526 ss_0_34 vss 1.29276e-16
C4527 ss_0_33 vss 1.29276e-16
C4528 ss_0_35 vss 1.29276e-16
C4529 ss_0_34 vss 1.29276e-16
C4530 ss_0_5 vss 2.71642e-17
C4531 ss_0_4 vss 2.71642e-17
C4532 ss_0_2 vss 1.21281e-16
C4533 ss_0_1 vss 1.21281e-16
C4534 ss_0 vss 5.86844e-17
C4535 ss_0_2 vss 5.86844e-17

R91_1 n2837 n2837_18 0.001
R91_2 n2837_17 n2837_7 0.001
R91_3 n2837_12 n2837_9 0.001
R91_4 n2837_15 n2837_14 0.001
R91_5 n2837_13 n2837_11 0.001
R91_6 n2837_6 n2837_4 0.001
R91_7 n2837_3 n2837_2 0.001
R91_8 n2837_10 n2837_9 43.2
R91_9 n2837_12 n2837_11 0.54
R91_10 n2837_6 n2837_5 36
R91_11 n2837_4 n2837_3 0.108
R91_12 n2837_14 n2837_13 57.6
R91_13 n2837_7 n2837_6 93.6
R91_14 n2837_16 n2837_15 0.54
R91_15 n2837_8 n2837_7 86.4
R91_16 n2837_17 n2837_16 0.972
R91_17 n2837_18 n2837_17 0.216

C4536 n2837_10 vss 5.086e-17
C4537 n2837_9 vss 5.086e-17
C4538 n2837_12 vss 5.43283e-17
C4539 n2837_11 vss 5.43283e-17
C4540 n2837_6 vss 3.9123e-17
C4541 n2837_5 vss 3.9123e-17
C4542 n2837_4 vss 2.92378e-17
C4543 n2837_3 vss 2.92378e-17
C4544 n2837_14 vss 6.25968e-17
C4545 n2837_13 vss 6.25968e-17
C4546 n2837_7 vss 1.0172e-16
C4547 n2837_6 vss 1.0172e-16
C4548 n2837_16 vss 5.43283e-17
C4549 n2837_15 vss 5.43283e-17
C4550 n2837_8 vss 9.97636e-17
C4551 n2837_7 vss 9.97636e-17
C4552 n2837_17 vss 1.00168e-16
C4553 n2837_16 vss 1.00168e-16
C4554 n2837_18 vss 2.71642e-17
C4555 n2837_17 vss 2.71642e-17

R92_1 n2848 n2848_5 0.001
R92_2 n2848_4 n2848_2 0.001
R92_3 n2848_3 n2848_2 0.001
R92_4 n2848_4 n2848_3 0.108
R92_5 n2848_5 n2848_4 1.188

C4556 n2848_4 vss 2.92378e-17
C4557 n2848_3 vss 2.92378e-17
C4558 n2848_5 vss 1.22239e-16
C4559 n2848_4 vss 1.22239e-16

R93_1 core_l0_dff_m core_l0_dff_m_12 0.001
R93_2 core_l0_dff_m_7 core_l0_dff_m_2 0.001
R93_3 core_l0_dff_m_6 core_l0_dff_m_4 0.001
R93_4 core_l0_dff_m_4 core_l0_dff_m_3 64.8
R93_5 core_l0_dff_m_5 core_l0_dff_m_4 93.6
R93_6 core_l0_dff_m_8 core_l0_dff_m_6 0.648
R93_7 core_l0_dff_m_8 core_l0_dff_m_7 0.216
R93_8 core_l0_dff_m_9 core_l0_dff_m_8 0.108
R93_9 core_l0_dff_m_10 core_l0_dff_m_9 0.648
R93_10 core_l0_dff_m_10 core_l0_dff_m_11 0.108
R93_11 core_l0_dff_m_12 core_l0_dff_m_11 0.216

C4560 core_l0_dff_m_4 vss 7.04214e-17
C4561 core_l0_dff_m_3 vss 7.04214e-17
C4562 core_l0_dff_m_5 vss 1.0172e-16
C4563 core_l0_dff_m_4 vss 1.0172e-16
C4564 core_l0_dff_m_8 vss 6.79104e-17
C4565 core_l0_dff_m_6 vss 6.79104e-17
C4566 core_l0_dff_m_8 vss 2.71642e-17
C4567 core_l0_dff_m_7 vss 2.71642e-17
C4568 core_l0_dff_m_9 vss 1.35821e-17
C4569 core_l0_dff_m_8 vss 1.35821e-17
C4570 core_l0_dff_m_10 vss 6.79104e-17
C4571 core_l0_dff_m_9 vss 6.79104e-17
C4572 core_l0_dff_m_10 vss 1.35821e-17
C4573 core_l0_dff_m_11 vss 1.35821e-17
C4574 core_l0_dff_m_12 vss 2.71642e-17
C4575 core_l0_dff_m_11 vss 2.71642e-17

R94_1 core_carry_2_13 core_carry_2_11 0.001
R94_2 core_carry_2_12 core_carry_2_15 0.001
R94_3 core_carry_2_14 core_carry_2_17 0.001
R94_4 core_carry_2_16 core_carry_2_22 0.001
R94_5 core_carry_2_6 core_carry_2 0.001
R94_6 core_carry_2_8 core_carry_2_5 0.001
R94_7 core_carry_2_19 core_carry_2_29 0.001
R94_8 core_carry_2_28 core_carry_2_25 0.001
R94_9 core_carry_2_27 core_carry_2_33 0.001
R94_10 core_carry_2_4 core_carry_2_2 0.001
R94_11 core_carry_2_3 core_carry_2_2 0.001
R94_12 core_carry_2_32 core_carry_2_30 115.2
R94_13 core_carry_2_31 core_carry_2_32 64.8
R94_14 core_carry_2_33 core_carry_2_32 7.2
R94_15 core_carry_2_26 core_carry_2_23 115.2
R94_16 core_carry_2_24 core_carry_2_26 43.2
R94_17 core_carry_2_26 core_carry_2_25 7.2
R94_18 core_carry_2_28 core_carry_2_27 0.756
R94_19 core_carry_2_29 core_carry_2_28 0.108
R94_20 core_carry_2_19 core_carry_2_18 0.756
R94_21 core_carry_2_20 core_carry_2_19 0.324
R94_22 core_carry_2_21 core_carry_2_20 0.054
R94_23 core_carry_2_22 core_carry_2_21 0.108
R94_24 core_carry_2_17 core_carry_2_16 1.188
R94_25 core_carry_2_4 core_carry_2_3 0.216
R94_26 core_carry_2_5 core_carry_2_4 0.324
R94_27 core_carry_2_6 core_carry_2_5 0.108
R94_28 core_carry_2_15 core_carry_2_14 0.27
R94_29 core_carry_2_8 core_carry_2_7 0.702
R94_30 core_carry_2_9 core_carry_2_8 0.378
R94_31 core_carry_2_10 core_carry_2_9 0.054
R94_32 core_carry_2_11 core_carry_2_10 0.378
R94_33 core_carry_2_13 core_carry_2_12 1.62

C4576 core_carry_2_32 vss 1.25194e-16
C4577 core_carry_2_30 vss 1.25194e-16
C4578 core_carry_2_31 vss 7.43336e-17
C4579 core_carry_2_32 vss 7.43336e-17
C4580 core_carry_2_33 vss 3.15414e-17
C4581 core_carry_2_32 vss 3.15414e-17
C4582 core_carry_2_26 vss 1.25194e-16
C4583 core_carry_2_23 vss 1.25194e-16
C4584 core_carry_2_24 vss 5.086e-17
C4585 core_carry_2_26 vss 5.086e-17
C4586 core_carry_2_26 vss 3.15414e-17
C4587 core_carry_2_25 vss 3.15414e-17
C4588 core_carry_2_28 vss 8.14925e-17
C4589 core_carry_2_27 vss 8.14925e-17
C4590 core_carry_2_29 vss 3.65472e-17
C4591 core_carry_2_28 vss 3.65472e-17
C4592 core_carry_2_19 vss 1.78524e-16
C4593 core_carry_2_18 vss 1.78524e-16
C4594 core_carry_2_20 vss 8.0028e-17
C4595 core_carry_2_19 vss 8.0028e-17
C4596 core_carry_2_21 vss 1.2312e-17
C4597 core_carry_2_20 vss 1.2312e-17
C4598 core_carry_2_22 vss 3.078e-17
C4599 core_carry_2_21 vss 3.078e-17
C4600 core_carry_2_17 vss 1.22239e-16
C4601 core_carry_2_16 vss 1.22239e-16
C4602 core_carry_2_4 vss 4.38566e-17
C4603 core_carry_2_3 vss 4.38566e-17
C4604 core_carry_2_5 vss 6.5785e-17
C4605 core_carry_2_4 vss 6.5785e-17
C4606 core_carry_2_6 vss 3.65472e-17
C4607 core_carry_2_5 vss 3.65472e-17
C4608 core_carry_2_15 vss 6.156e-17
C4609 core_carry_2_14 vss 6.156e-17
C4610 core_carry_2_8 vss 1.66212e-16
C4611 core_carry_2_7 vss 1.66212e-16
C4612 core_carry_2_9 vss 9.234e-17
C4613 core_carry_2_8 vss 9.234e-17
C4614 core_carry_2_10 vss 1.2312e-17
C4615 core_carry_2_9 vss 1.2312e-17
C4616 core_carry_2_11 vss 9.234e-17
C4617 core_carry_2_10 vss 9.234e-17
C4618 core_carry_2_13 vss 1.62985e-16
C4619 core_carry_2_12 vss 1.62985e-16

R95_1 core_int_8_13 core_int_8_5 0.001
R95_2 core_int_8_12 core_int_8_22 0.001
R95_3 core_int_8_2 core_int_8_10 0.001
R95_4 core_int_8_11 core_int_8 0.001
R95_5 core_int_8_9 core_int_8_7 0.001
R95_6 core_int_8_8 core_int_8_7 0.001
R95_7 core_int_8_19 core_int_8_16 0.001
R95_8 core_int_8_17 core_int_8_14 0.001
R95_9 core_int_8_15 core_int_8_14 136.8
R95_10 core_int_8_17 core_int_8_16 0.324
R95_11 core_int_8_9 core_int_8_8 0.216
R95_12 core_int_8_10 core_int_8_9 0.216
R95_13 core_int_8_11 core_int_8_10 0.216
R95_14 core_int_8_2 core_int_8_1 0.648
R95_15 core_int_8_3 core_int_8_2 0.432
R95_16 core_int_8_19 core_int_8_18 0.432
R95_17 core_int_8_20 core_int_8_19 0.702
R95_18 core_int_8_4 core_int_8_3 0.054
R95_19 core_int_8_5 core_int_8_4 0.54
R95_20 core_int_8_21 core_int_8_20 0.054
R95_21 core_int_8_22 core_int_8_21 0.54
R95_22 core_int_8_13 core_int_8_12 6.048

C4620 core_int_8_15 vss 1.54536e-16
C4621 core_int_8_14 vss 1.54536e-16
C4622 core_int_8_17 vss 3.90485e-17
C4623 core_int_8_16 vss 3.90485e-17
C4624 core_int_8_9 vss 4.38566e-17
C4625 core_int_8_8 vss 4.38566e-17
C4626 core_int_8_10 vss 5.11661e-17
C4627 core_int_8_9 vss 5.11661e-17
C4628 core_int_8_11 vss 5.11661e-17
C4629 core_int_8_10 vss 5.11661e-17
C4630 core_int_8_2 vss 1.539e-16
C4631 core_int_8_1 vss 1.539e-16
C4632 core_int_8_3 vss 1.04652e-16
C4633 core_int_8_2 vss 1.04652e-16
C4634 core_int_8_19 vss 9.8496e-17
C4635 core_int_8_18 vss 9.8496e-17
C4636 core_int_8_20 vss 1.60056e-16
C4637 core_int_8_19 vss 1.60056e-16
C4638 core_int_8_4 vss 1.2312e-17
C4639 core_int_8_3 vss 1.2312e-17
C4640 core_int_8_5 vss 1.2312e-16
C4641 core_int_8_4 vss 1.2312e-16
C4642 core_int_8_21 vss 1.2312e-17
C4643 core_int_8_20 vss 1.2312e-17
C4644 core_int_8_22 vss 1.2312e-16
C4645 core_int_8_21 vss 1.2312e-16
C4646 core_int_8_13 vss 6.11194e-16
C4647 core_int_8_12 vss 6.11194e-16

R96_1 core_carry_1_13 core_carry_1_5 0.001
R96_2 core_carry_1_12 core_carry_1_15 0.001
R96_3 core_carry_1_14 core_carry_1_41 0.001
R96_4 core_carry_1_40 core_carry_1_26 0.001
R96_5 core_carry_1_39 core_carry_1_37 0.001
R96_6 core_carry_1_38 core_carry_1_46 0.001
R96_7 core_carry_1_2 core_carry_1_10 0.001
R96_8 core_carry_1_11 core_carry_1 0.001
R96_9 core_carry_1_43 core_carry_1_53 0.001
R96_10 core_carry_1_19 core_carry_1_17 0.001
R96_11 core_carry_1_30 core_carry_1_28 0.001
R96_12 core_carry_1_52 core_carry_1_49 0.001
R96_13 core_carry_1_51 core_carry_1_57 0.001
R96_14 core_carry_1_9 core_carry_1_7 0.001
R96_15 core_carry_1_8 core_carry_1_7 0.001
R96_16 core_carry_1_23 core_carry_1_21 0.001
R96_17 core_carry_1_34 core_carry_1_32 0.001
R96_18 core_carry_1_17 core_carry_1_16 72
R96_19 core_carry_1_18 core_carry_1_17 50.4
R96_20 core_carry_1_28 core_carry_1_27 72
R96_21 core_carry_1_29 core_carry_1_28 50.4
R96_22 core_carry_1_56 core_carry_1_54 115.2
R96_23 core_carry_1_55 core_carry_1_56 64.8
R96_24 core_carry_1_57 core_carry_1_56 7.2
R96_25 core_carry_1_50 core_carry_1_47 115.2
R96_26 core_carry_1_48 core_carry_1_50 43.2
R96_27 core_carry_1_19 core_carry_1_20 0.216
R96_28 core_carry_1_30 core_carry_1_31 0.216
R96_29 core_carry_1_50 core_carry_1_49 7.2
R96_30 core_carry_1_21 core_carry_1_20 0.216
R96_31 core_carry_1_32 core_carry_1_31 0.216
R96_32 core_carry_1_52 core_carry_1_51 0.756
R96_33 core_carry_1_53 core_carry_1_52 0.108
R96_34 core_carry_1_23 core_carry_1_22 0.486
R96_35 core_carry_1_24 core_carry_1_23 0.648
R96_36 core_carry_1_34 core_carry_1_33 0.486
R96_37 core_carry_1_35 core_carry_1_34 0.648
R96_38 core_carry_1_43 core_carry_1_42 0.756
R96_39 core_carry_1_44 core_carry_1_43 0.324
R96_40 core_carry_1_25 core_carry_1_24 0.054
R96_41 core_carry_1_26 core_carry_1_25 0.27
R96_42 core_carry_1_36 core_carry_1_35 0.054
R96_43 core_carry_1_37 core_carry_1_36 0.27
R96_44 core_carry_1_45 core_carry_1_44 0.054
R96_45 core_carry_1_46 core_carry_1_45 0.27
R96_46 core_carry_1_39 core_carry_1_38 1.944
R96_47 core_carry_1_40 core_carry_1_39 1.62
R96_48 core_carry_1_41 core_carry_1_40 1.62
R96_49 core_carry_1_9 core_carry_1_8 0.216
R96_50 core_carry_1_10 core_carry_1_9 0.324
R96_51 core_carry_1_11 core_carry_1_10 0.108
R96_52 core_carry_1_15 core_carry_1_14 0.27
R96_53 core_carry_1_2 core_carry_1_1 0.702
R96_54 core_carry_1_3 core_carry_1_2 0.378
R96_55 core_carry_1_4 core_carry_1_3 0.054
R96_56 core_carry_1_5 core_carry_1_4 0.54
R96_57 core_carry_1_13 core_carry_1_12 0.756

C4648 core_carry_1_17 vss 8.21582e-17
C4649 core_carry_1_16 vss 8.21582e-17
C4650 core_carry_1_18 vss 5.86844e-17
C4651 core_carry_1_17 vss 5.86844e-17
C4652 core_carry_1_28 vss 8.21582e-17
C4653 core_carry_1_27 vss 8.21582e-17
C4654 core_carry_1_29 vss 5.86844e-17
C4655 core_carry_1_28 vss 5.86844e-17
C4656 core_carry_1_56 vss 1.25194e-16
C4657 core_carry_1_54 vss 1.25194e-16
C4658 core_carry_1_55 vss 7.43336e-17
C4659 core_carry_1_56 vss 7.43336e-17
C4660 core_carry_1_57 vss 3.15414e-17
C4661 core_carry_1_56 vss 3.15414e-17
C4662 core_carry_1_50 vss 1.25194e-16
C4663 core_carry_1_47 vss 1.25194e-16
C4664 core_carry_1_48 vss 5.086e-17
C4665 core_carry_1_50 vss 5.086e-17
C4666 core_carry_1_19 vss 2.71642e-17
C4667 core_carry_1_20 vss 2.71642e-17
C4668 core_carry_1_30 vss 2.71642e-17
C4669 core_carry_1_31 vss 2.71642e-17
C4670 core_carry_1_50 vss 3.15414e-17
C4671 core_carry_1_49 vss 3.15414e-17
C4672 core_carry_1_21 vss 2.54664e-17
C4673 core_carry_1_20 vss 2.54664e-17
C4674 core_carry_1_32 vss 2.54664e-17
C4675 core_carry_1_31 vss 2.54664e-17
C4676 core_carry_1_52 vss 8.14925e-17
C4677 core_carry_1_51 vss 8.14925e-17
C4678 core_carry_1_53 vss 3.65472e-17
C4679 core_carry_1_52 vss 3.65472e-17
C4680 core_carry_1_23 vss 1.10808e-16
C4681 core_carry_1_22 vss 1.10808e-16
C4682 core_carry_1_24 vss 1.47744e-16
C4683 core_carry_1_23 vss 1.47744e-16
C4684 core_carry_1_34 vss 1.10808e-16
C4685 core_carry_1_33 vss 1.10808e-16
C4686 core_carry_1_35 vss 1.47744e-16
C4687 core_carry_1_34 vss 1.47744e-16
C4688 core_carry_1_43 vss 1.78524e-16
C4689 core_carry_1_42 vss 1.78524e-16
C4690 core_carry_1_44 vss 8.0028e-17
C4691 core_carry_1_43 vss 8.0028e-17
C4692 core_carry_1_25 vss 1.2312e-17
C4693 core_carry_1_24 vss 1.2312e-17
C4694 core_carry_1_26 vss 6.156e-17
C4695 core_carry_1_25 vss 6.156e-17
C4696 core_carry_1_36 vss 1.2312e-17
C4697 core_carry_1_35 vss 1.2312e-17
C4698 core_carry_1_37 vss 6.156e-17
C4699 core_carry_1_36 vss 6.156e-17
C4700 core_carry_1_45 vss 1.2312e-17
C4701 core_carry_1_44 vss 1.2312e-17
C4702 core_carry_1_46 vss 6.156e-17
C4703 core_carry_1_45 vss 6.156e-17
C4704 core_carry_1_39 vss 2.03731e-16
C4705 core_carry_1_38 vss 2.03731e-16
C4706 core_carry_1_40 vss 1.62985e-16
C4707 core_carry_1_39 vss 1.62985e-16
C4708 core_carry_1_41 vss 1.62985e-16
C4709 core_carry_1_40 vss 1.62985e-16
C4710 core_carry_1_9 vss 4.38566e-17
C4711 core_carry_1_8 vss 4.38566e-17
C4712 core_carry_1_10 vss 6.5785e-17
C4713 core_carry_1_9 vss 6.5785e-17
C4714 core_carry_1_11 vss 3.65472e-17
C4715 core_carry_1_10 vss 3.65472e-17
C4716 core_carry_1_15 vss 6.156e-17
C4717 core_carry_1_14 vss 6.156e-17
C4718 core_carry_1_2 vss 1.66212e-16
C4719 core_carry_1_1 vss 1.66212e-16
C4720 core_carry_1_3 vss 9.234e-17
C4721 core_carry_1_2 vss 9.234e-17
C4722 core_carry_1_4 vss 1.2312e-17
C4723 core_carry_1_3 vss 1.2312e-17
C4724 core_carry_1_5 vss 1.2312e-16
C4725 core_carry_1_4 vss 1.2312e-16
C4726 core_carry_1_13 vss 8.14925e-17
C4727 core_carry_1_12 vss 8.14925e-17

R97_1 core_int_4_13 core_int_4_5 0.001
R97_2 core_int_4_12 core_int_4_22 0.001
R97_3 core_int_4_2 core_int_4_10 0.001
R97_4 core_int_4_11 core_int_4 0.001
R97_5 core_int_4_8 core_int_4_7 0.001
R97_6 core_int_4_9 core_int_4_7 0.001
R97_7 core_int_4_19 core_int_4_16 0.001
R97_8 core_int_4_17 core_int_4_14 0.001
R97_9 core_int_4_15 core_int_4_14 136.8
R97_10 core_int_4_17 core_int_4_16 0.324
R97_11 core_int_4_9 core_int_4_8 0.216
R97_12 core_int_4_10 core_int_4_9 0.216
R97_13 core_int_4_11 core_int_4_10 0.216
R97_14 core_int_4_19 core_int_4_18 0.432
R97_15 core_int_4_20 core_int_4_19 0.702
R97_16 core_int_4_21 core_int_4_20 0.054
R97_17 core_int_4_22 core_int_4_21 0.378
R97_18 core_int_4_2 core_int_4_1 0.648
R97_19 core_int_4_3 core_int_4_2 0.432
R97_20 core_int_4_4 core_int_4_3 0.054
R97_21 core_int_4_5 core_int_4_4 0.378
R97_22 core_int_4_13 core_int_4_12 5.184

C4728 core_int_4_15 vss 1.54536e-16
C4729 core_int_4_14 vss 1.54536e-16
C4730 core_int_4_17 vss 3.90485e-17
C4731 core_int_4_16 vss 3.90485e-17
C4732 core_int_4_9 vss 4.38566e-17
C4733 core_int_4_8 vss 4.38566e-17
C4734 core_int_4_10 vss 5.11661e-17
C4735 core_int_4_9 vss 5.11661e-17
C4736 core_int_4_11 vss 5.11661e-17
C4737 core_int_4_10 vss 5.11661e-17
C4738 core_int_4_19 vss 9.8496e-17
C4739 core_int_4_18 vss 9.8496e-17
C4740 core_int_4_20 vss 1.60056e-16
C4741 core_int_4_19 vss 1.60056e-16
C4742 core_int_4_21 vss 1.2312e-17
C4743 core_int_4_20 vss 1.2312e-17
C4744 core_int_4_22 vss 9.234e-17
C4745 core_int_4_21 vss 9.234e-17
C4746 core_int_4_2 vss 1.539e-16
C4747 core_int_4_1 vss 1.539e-16
C4748 core_int_4_3 vss 1.04652e-16
C4749 core_int_4_2 vss 1.04652e-16
C4750 core_int_4_4 vss 1.2312e-17
C4751 core_int_4_3 vss 1.2312e-17
C4752 core_int_4_5 vss 9.234e-17
C4753 core_int_4_4 vss 9.234e-17
C4754 core_int_4_13 vss 5.29701e-16
C4755 core_int_4_12 vss 5.29701e-16

R98_1 n3019_2 n3019_33 0.001
R98_2 n3019_20 n3019_6 0.001
R98_3 n3019_1 n3019_32 0.001
R98_4 n3019_29 n3019_5 0.001
R98_5 n3019_39 n3019_9 0.001
R98_6 n3019_38 n3019_9 0.001
R98_7 n3019_36 n3019_9 0.001
R98_8 n3019_37 n3019_9 0.001
R98_9 n3019_35 n3019_9 0.001
R98_10 n3019_26 n3019_10 0.001
R98_11 n3019_27 n3019_10 0.001
R98_12 n3019_28 n3019_10 0.001
R98_13 n3019_24 n3019_10 0.001
R98_14 n3019_25 n3019_12 0.001
R98_15 n3019_18 n3019_13 0.001
R98_16 n3019_17 n3019_13 0.001
R98_17 n3019_16 n3019_13 0.001
R98_18 n3019_11 n3019_15 0.001
R98_19 n3019_14 n3019_13 0.001
R98_20 n3019_6 n3019_5 7.2
R98_21 n3019_7 n3019_6 21.6
R98_22 n3019 n3019_7 0.001
R98_23 n3019_14 n3019_22 0.324
R98_24 n3019_15 n3019_14 0.108
R98_25 n3019_16 n3019_15 0.108
R98_26 n3019_17 n3019_16 0.108
R98_27 n3019_18 n3019_17 0.108
R98_28 n3019_19 n3019_18 0.001
R98_29 n3019_12 n3019_11 0.216
R98_30 n3019_20 n3019_29 0.108
R98_31 n3019_21 n3019_20 0.001
R98_32 n3019_23 n3019_22 0.324
R98_33 n3019_24 n3019_23 0.324
R98_34 n3019_25 n3019_24 0.108
R98_35 n3019_26 n3019_25 0.108
R98_36 n3019_27 n3019_26 0.108
R98_37 n3019_28 n3019_27 0.108
R98_38 n3019_29 n3019_28 0.108
R98_39 n3019_30 n3019_29 0.216
R98_40 n3019_31 n3019_30 0.108
R98_41 n3019_32 n3019_31 0.216
R98_42 n3019_35 n3019_32 0.108
R98_43 n3019_36 n3019_35 0.108
R98_44 n3019_37 n3019_36 0.108
R98_45 n3019_38 n3019_37 0.108
R98_46 n3019_39 n3019_38 0.108
R98_47 n3019_40 n3019_39 0.001
R98_48 n3019_33 n3019_32 0.108
R98_49 n3019_34 n3019_33 0.001
R98_50 n3019_2 n3019_1 7.2
R98_51 n3019_3 n3019_2 21.6
R98_52 n3019_4 n3019_3 0.001

C4756 n3019_6 vss 4.20552e-17
C4757 n3019_5 vss 4.20552e-17
C4758 n3019_7 vss 9.46242e-17
C4759 n3019_6 vss 9.46242e-17
C4760 n3019 vss 3.05111e-16
C4761 n3019_7 vss 3.05111e-16
C4762 n3019_14 vss 1.0959e-16
C4763 n3019_22 vss 1.0959e-16
C4764 n3019_15 vss 3.91392e-17
C4765 n3019_14 vss 3.91392e-17
C4766 n3019_16 vss 3.91392e-17
C4767 n3019_15 vss 3.91392e-17
C4768 n3019_17 vss 3.91392e-17
C4769 n3019_16 vss 3.91392e-17
C4770 n3019_18 vss 3.91392e-17
C4771 n3019_17 vss 3.91392e-17
C4772 n3019_19 vss 1.40901e-17
C4773 n3019_18 vss 1.40901e-17
C4774 n3019_12 vss 7.81488e-17
C4775 n3019_11 vss 7.81488e-17
C4776 n3019_20 vss 3.71822e-17
C4777 n3019_29 vss 3.71822e-17
C4778 n3019_21 vss 1.40901e-17
C4779 n3019_20 vss 1.40901e-17
C4780 n3019_23 vss 9.39341e-17
C4781 n3019_22 vss 9.39341e-17
C4782 n3019_24 vss 1.0959e-16
C4783 n3019_23 vss 1.0959e-16
C4784 n3019_25 vss 3.91392e-17
C4785 n3019_24 vss 3.91392e-17
C4786 n3019_26 vss 3.91392e-17
C4787 n3019_25 vss 3.91392e-17
C4788 n3019_27 vss 3.91392e-17
C4789 n3019_26 vss 3.91392e-17
C4790 n3019_28 vss 3.91392e-17
C4791 n3019_27 vss 3.91392e-17
C4792 n3019_29 vss 4.6967e-17
C4793 n3019_28 vss 4.6967e-17
C4794 n3019_30 vss 5.63604e-17
C4795 n3019_29 vss 5.63604e-17
C4796 n3019_31 vss 2.81802e-17
C4797 n3019_30 vss 2.81802e-17
C4798 n3019_32 vss 6.41883e-17
C4799 n3019_31 vss 6.41883e-17
C4800 n3019_35 vss 4.6967e-17
C4801 n3019_32 vss 4.6967e-17
C4802 n3019_36 vss 3.91392e-17
C4803 n3019_35 vss 3.91392e-17
C4804 n3019_37 vss 4.6967e-17
C4805 n3019_36 vss 4.6967e-17
C4806 n3019_38 vss 3.91392e-17
C4807 n3019_37 vss 3.91392e-17
C4808 n3019_39 vss 3.91392e-17
C4809 n3019_38 vss 3.91392e-17
C4810 n3019_40 vss 1.40901e-17
C4811 n3019_39 vss 1.40901e-17
C4812 n3019_33 vss 3.71822e-17
C4813 n3019_32 vss 3.71822e-17
C4814 n3019_34 vss 1.40901e-17
C4815 n3019_33 vss 1.40901e-17
C4816 n3019_2 vss 4.20552e-17
C4817 n3019_1 vss 4.20552e-17
C4818 n3019_3 vss 9.46242e-17
C4819 n3019_2 vss 9.46242e-17
C4820 n3019_4 vss 5.47139e-16
C4821 n3019_3 vss 5.47139e-16

R99_1 n3051_2 n3051_9 0.001
R99_2 n3051_6 n3051_1 0.001
R99_3 n3051_2 n3051_7 0.001
R99_4 n3051_4 n3051 0.001
R99_5 n3051_5 n3051_4 0.756
R99_6 n3051_6 n3051_5 0.108
R99_7 n3051_8 n3051_6 0.756
R99_8 n3051_8 n3051_7 0.108
R99_9 n3051_9 n3051_8 0.108

C4822 n3051_5 vss 8.14925e-17
C4823 n3051_4 vss 8.14925e-17
C4824 n3051_6 vss 2.37557e-17
C4825 n3051_5 vss 2.37557e-17
C4826 n3051_8 vss 8.14925e-17
C4827 n3051_6 vss 8.14925e-17
C4828 n3051_8 vss 2.19283e-17
C4829 n3051_7 vss 2.19283e-17
C4830 n3051_9 vss 2.19283e-17
C4831 n3051_8 vss 2.19283e-17

R100_1 n3062_1 n3062_4 0.001
R100_2 n3062_3 n3062 0.001
R100_3 n3062_4 n3062_3 0.756

C4832 n3062_4 vss 8.14925e-17
C4833 n3062_3 vss 8.14925e-17

R101_1 n3071_2 n3071_9 0.001
R101_2 n3071_6 n3071_1 0.001
R101_3 n3071_2 n3071_7 0.001
R101_4 n3071_4 n3071 0.001
R101_5 n3071_5 n3071_4 0.756
R101_6 n3071_6 n3071_5 0.108
R101_7 n3071_8 n3071_6 0.756
R101_8 n3071_8 n3071_7 0.108
R101_9 n3071_9 n3071_8 0.108

C4834 n3071_5 vss 8.14925e-17
C4835 n3071_4 vss 8.14925e-17
C4836 n3071_6 vss 2.37557e-17
C4837 n3071_5 vss 2.37557e-17
C4838 n3071_8 vss 8.14925e-17
C4839 n3071_6 vss 8.14925e-17
C4840 n3071_8 vss 2.19283e-17
C4841 n3071_7 vss 2.19283e-17
C4842 n3071_9 vss 2.19283e-17
C4843 n3071_8 vss 2.19283e-17

R102_1 n3082_1 n3082_4 0.001
R102_2 n3082_3 n3082 0.001
R102_3 n3082_4 n3082_3 0.756

C4844 n3082_4 vss 8.14925e-17
C4845 n3082_3 vss 8.14925e-17

R103_1 n3091_2 n3091_9 0.001
R103_2 n3091_6 n3091_1 0.001
R103_3 n3091_2 n3091_7 0.001
R103_4 n3091_4 n3091 0.001
R103_5 n3091_5 n3091_4 0.756
R103_6 n3091_6 n3091_5 0.108
R103_7 n3091_8 n3091_6 0.756
R103_8 n3091_8 n3091_7 0.108
R103_9 n3091_9 n3091_8 0.108

C4846 n3091_5 vss 8.14925e-17
C4847 n3091_4 vss 8.14925e-17
C4848 n3091_6 vss 2.37557e-17
C4849 n3091_5 vss 2.37557e-17
C4850 n3091_8 vss 8.14925e-17
C4851 n3091_6 vss 8.14925e-17
C4852 n3091_8 vss 2.19283e-17
C4853 n3091_7 vss 2.19283e-17
C4854 n3091_9 vss 2.19283e-17
C4855 n3091_8 vss 2.19283e-17

R104_1 n3102_5 n3102_2 0.001
R104_2 n3102_1 n3102_9 0.001
R104_3 n3102_4 n3102_2 0.001
R104_4 n3102_6 n3102 0.001
R104_5 n3102_7 n3102_4 0.108
R104_6 n3102_5 n3102_7 0.108
R104_7 n3102_8 n3102_6 0.756
R104_8 n3102_7 n3102_9 0.756
R104_9 n3102_9 n3102_8 0.108

C4856 n3102_7 vss 2.19283e-17
C4857 n3102_4 vss 2.19283e-17
C4858 n3102_5 vss 2.19283e-17
C4859 n3102_7 vss 2.19283e-17
C4860 n3102_8 vss 8.14925e-17
C4861 n3102_6 vss 8.14925e-17
C4862 n3102_7 vss 8.14925e-17
C4863 n3102_9 vss 8.14925e-17
C4864 n3102_9 vss 2.37557e-17
C4865 n3102_8 vss 2.37557e-17

R105_1 n3113_1 n3113_4 0.001
R105_2 n3113_3 n3113 0.001
R105_3 n3113_4 n3113_3 0.756

C4866 n3113_4 vss 8.14925e-17
C4867 n3113_3 vss 8.14925e-17

R106_1 core_mux_3 core_mux_3_6 0.001
R106_2 core_mux_3_4 core_mux_3_2 0.001
R106_3 core_mux_3_5 core_mux_3_12 0.001
R106_4 core_mux_3_3 core_mux_3_2 0.001
R106_5 core_mux_3_8 core_mux_3_21 0.001
R106_6 core_mux_3_9 core_mux_3_7 0.001
R106_7 core_mux_3_25 core_mux_3_15 0.001
R106_8 core_mux_3_18 core_mux_3_29 0.001
R106_9 core_mux_3_28 core_mux_3_23 0.001
R106_10 core_mux_3_15 core_mux_3_14 115.2
R106_11 core_mux_3_16 core_mux_3_15 43.2
R106_12 core_mux_3_25 core_mux_3_26 0.108
R106_13 core_mux_3_23 core_mux_3_22 115.2
R106_14 core_mux_3_24 core_mux_3_23 64.8
R106_15 core_mux_3_26 core_mux_3_27 1.62
R106_16 core_mux_3_28 core_mux_3_27 0.216
R106_17 core_mux_3_29 core_mux_3_28 0.216
R106_18 core_mux_3_18 core_mux_3_17 0.81
R106_19 core_mux_3_19 core_mux_3_18 0.324
R106_20 core_mux_3_20 core_mux_3_19 0.054
R106_21 core_mux_3_21 core_mux_3_20 0.918
R106_22 core_mux_3_8 core_mux_3_7 0.756
R106_23 core_mux_3_10 core_mux_3_9 0.108
R106_24 core_mux_3_11 core_mux_3_10 0.054
R106_25 core_mux_3_12 core_mux_3_11 0.648
R106_26 core_mux_3_13 core_mux_3_12 0.486
R106_27 core_mux_3_4 core_mux_3_3 0.216
R106_28 core_mux_3_5 core_mux_3_4 0.324
R106_29 core_mux_3_6 core_mux_3_5 0.216

C4868 core_mux_3_15 vss 1.25194e-16
C4869 core_mux_3_14 vss 1.25194e-16
C4870 core_mux_3_16 vss 5.086e-17
C4871 core_mux_3_15 vss 5.086e-17
C4872 core_mux_3_25 vss 2.92378e-17
C4873 core_mux_3_26 vss 2.92378e-17
C4874 core_mux_3_23 vss 1.25194e-16
C4875 core_mux_3_22 vss 1.25194e-16
C4876 core_mux_3_24 vss 7.43336e-17
C4877 core_mux_3_23 vss 7.43336e-17
C4878 core_mux_3_26 vss 1.69776e-16
C4879 core_mux_3_27 vss 1.69776e-16
C4880 core_mux_3_28 vss 2.71642e-17
C4881 core_mux_3_27 vss 2.71642e-17
C4882 core_mux_3_29 vss 4.38566e-17
C4883 core_mux_3_28 vss 4.38566e-17
C4884 core_mux_3_18 vss 1.8468e-16
C4885 core_mux_3_17 vss 1.8468e-16
C4886 core_mux_3_19 vss 7.3872e-17
C4887 core_mux_3_18 vss 7.3872e-17
C4888 core_mux_3_20 vss 1.2312e-17
C4889 core_mux_3_19 vss 1.2312e-17
C4890 core_mux_3_21 vss 2.1546e-16
C4891 core_mux_3_20 vss 2.1546e-16
C4892 core_mux_3_8 vss 8.14925e-17
C4893 core_mux_3_7 vss 8.14925e-17
C4894 core_mux_3_10 vss 3.078e-17
C4895 core_mux_3_9 vss 3.078e-17
C4896 core_mux_3_11 vss 1.2312e-17
C4897 core_mux_3_10 vss 1.2312e-17
C4898 core_mux_3_12 vss 1.47744e-16
C4899 core_mux_3_11 vss 1.47744e-16
C4900 core_mux_3_13 vss 1.10808e-16
C4901 core_mux_3_12 vss 1.10808e-16
C4902 core_mux_3_4 vss 4.38566e-17
C4903 core_mux_3_3 vss 4.38566e-17
C4904 core_mux_3_5 vss 5.84755e-17
C4905 core_mux_3_4 vss 5.84755e-17
C4906 core_mux_3_6 vss 4.38566e-17
C4907 core_mux_3_5 vss 4.38566e-17

R107_1 core_regout_3_3 core_regout_3_15 0.001
R107_2 core_regout_3_14 core_regout_3_17 0.001
R107_3 core_regout_3_16 core_regout_3_19 0.001
R107_4 core_regout_3_18 core_regout_3_29 0.001
R107_5 core_regout_3 core_regout_3_13 0.001
R107_6 core_regout_3 core_regout_3_11 0.001
R107_7 core_regout_3_26 core_regout_3_21 0.001
R107_8 core_regout_3_20 core_regout_3_23 0.001
R107_9 core_regout_3_10 core_regout_3_2 0.001
R107_10 core_regout_3_8 core_regout_3_2 0.001
R107_11 core_regout_3_9 core_regout_3_5 0.001
R107_12 core_regout_3_23 core_regout_3_22 72
R107_13 core_regout_3_24 core_regout_3_23 43.2
R107_14 core_regout_3_21 core_regout_3_20 0.108
R107_15 core_regout_3_26 core_regout_3_25 0.756
R107_16 core_regout_3_27 core_regout_3_26 0.324
R107_17 core_regout_3_28 core_regout_3_27 0.054
R107_18 core_regout_3_29 core_regout_3_28 0.108
R107_19 core_regout_3_19 core_regout_3_18 0.756
R107_20 core_regout_3_17 core_regout_3_16 0.108
R107_21 core_regout_3_15 core_regout_3_14 1.188
R107_22 core_regout_3_3 core_regout_3_7 0.27
R107_23 core_regout_3_5 core_regout_3_4 0.378
R107_24 core_regout_3_6 core_regout_3_5 0.702
R107_25 core_regout_3_7 core_regout_3_6 0.054
R107_26 core_regout_3_9 core_regout_3_8 0.108
R107_27 core_regout_3_10 core_regout_3_9 0.108
R107_28 core_regout_3_11 core_regout_3_10 0.648
R107_29 core_regout_3_12 core_regout_3_11 0.001
R107_30 core_regout_3_13 core_regout_3_12 0.001

C4908 core_regout_3_23 vss 8.21582e-17
C4909 core_regout_3_22 vss 8.21582e-17
C4910 core_regout_3_24 vss 5.086e-17
C4911 core_regout_3_23 vss 5.086e-17
C4912 core_regout_3_21 vss 3.65472e-17
C4913 core_regout_3_20 vss 3.65472e-17
C4914 core_regout_3_26 vss 1.78524e-16
C4915 core_regout_3_25 vss 1.78524e-16
C4916 core_regout_3_27 vss 8.0028e-17
C4917 core_regout_3_26 vss 8.0028e-17
C4918 core_regout_3_28 vss 1.2312e-17
C4919 core_regout_3_27 vss 1.2312e-17
C4920 core_regout_3_29 vss 3.078e-17
C4921 core_regout_3_28 vss 3.078e-17
C4922 core_regout_3_19 vss 8.14925e-17
C4923 core_regout_3_18 vss 8.14925e-17
C4924 core_regout_3_17 vss 3.078e-17
C4925 core_regout_3_16 vss 3.078e-17
C4926 core_regout_3_15 vss 1.22239e-16
C4927 core_regout_3_14 vss 1.22239e-16
C4928 core_regout_3_3 vss 6.156e-17
C4929 core_regout_3_7 vss 6.156e-17
C4930 core_regout_3_5 vss 9.234e-17
C4931 core_regout_3_4 vss 9.234e-17
C4932 core_regout_3_6 vss 1.66212e-16
C4933 core_regout_3_5 vss 1.66212e-16
C4934 core_regout_3_7 vss 1.2312e-17
C4935 core_regout_3_6 vss 1.2312e-17
C4936 core_regout_3_9 vss 2.19283e-17
C4937 core_regout_3_8 vss 2.19283e-17
C4938 core_regout_3_10 vss 2.19283e-17
C4939 core_regout_3_9 vss 2.19283e-17
C4940 core_regout_3_11 vss 7.47014e-17
C4941 core_regout_3_10 vss 7.47014e-17
C4942 core_regout_3_12 vss 1.3157e-17
C4943 core_regout_3_11 vss 1.3157e-17
C4944 core_regout_3_13 vss 1.60808e-17
C4945 core_regout_3_12 vss 1.60808e-17

R108_1 n3197_1 n3197_11 0.001
R108_2 n3197_7 n3197_5 0.001
R108_3 n3197_9 n3197_6 0.001
R108_4 n3197_4 n3197_2 72
R108_5 n3197 n3197_4 43.2
R108_6 n3197_5 n3197_4 7.2
R108_7 n3197_7 n3197_8 0.108
R108_8 n3197_9 n3197_8 0.756
R108_9 n3197_10 n3197_9 0.324
R108_10 n3197_11 n3197_10 0.648

C4946 n3197_4 vss 8.21582e-17
C4947 n3197_2 vss 8.21582e-17
C4948 n3197 vss 5.086e-17
C4949 n3197_4 vss 5.086e-17
C4950 n3197_5 vss 3.15414e-17
C4951 n3197_4 vss 3.15414e-17
C4952 n3197_7 vss 3.65472e-17
C4953 n3197_8 vss 3.65472e-17
C4954 n3197_9 vss 8.14925e-17
C4955 n3197_8 vss 8.14925e-17
C4956 n3197_10 vss 4.07462e-17
C4957 n3197_9 vss 4.07462e-17
C4958 n3197_11 vss 6.79104e-17
C4959 n3197_10 vss 6.79104e-17

R109_1 n3212 n3212_10 0.001
R109_2 n3212_7 n3212_4 0.001
R109_3 n3212_6 n3212_5 0.001
R109_4 n3212_2 n3212_4 144
R109_5 n3212_4 n3212_3 72
R109_6 n3212_7 n3212_6 0.216
R109_7 n3212_7 n3212_8 0.54
R109_8 n3212_9 n3212_8 0.648
R109_9 n3212_10 n3212_9 0.432

C4960 n3212_2 vss 1.6236e-16
C4961 n3212_4 vss 1.6236e-16
C4962 n3212_4 vss 7.8246e-17
C4963 n3212_3 vss 7.8246e-17
C4964 n3212_7 vss 3.22574e-17
C4965 n3212_6 vss 3.22574e-17
C4966 n3212_7 vss 5.60261e-17
C4967 n3212_8 vss 5.60261e-17
C4968 n3212_9 vss 7.47014e-17
C4969 n3212_8 vss 7.47014e-17
C4970 n3212_10 vss 4.75373e-17
C4971 n3212_9 vss 4.75373e-17

R110_1 n3223 n3223_12 0.001
R110_2 n3223_10 n3223_5 0.001
R110_3 n3223_8 n3223_6 0.001
R110_4 n3223_7 n3223_6 0.001
R110_5 n3223_2 n3223_3 72
R110_6 n3223_8 n3223_7 0.108
R110_7 n3223_4 n3223_3 64.8
R110_8 n3223_8 n3223_9 0.324
R110_9 n3223_5 n3223_4 21.6
R110_10 n3223_10 n3223_9 0.648
R110_11 n3223_11 n3223_10 0.324
R110_12 n3223_12 n3223_11 0.324

C4972 n3223_2 vss 8.21582e-17
C4973 n3223_3 vss 8.21582e-17
C4974 n3223_8 vss 3.10651e-17
C4975 n3223_7 vss 3.10651e-17
C4976 n3223_4 vss 7.04214e-17
C4977 n3223_3 vss 7.04214e-17
C4978 n3223_8 vss 4.07462e-17
C4979 n3223_9 vss 4.07462e-17
C4980 n3223_5 vss 2.34738e-17
C4981 n3223_4 vss 2.34738e-17
C4982 n3223_10 vss 7.47014e-17
C4983 n3223_9 vss 7.47014e-17
C4984 n3223_11 vss 3.39552e-17
C4985 n3223_10 vss 3.39552e-17
C4986 n3223_12 vss 4.07462e-17
C4987 n3223_11 vss 4.07462e-17

R111_1 core_l3_dff_s_1 core_l3_dff_s_6 0.001
R111_2 core_l3_dff_s_3 core_l3_dff_s_12 0.001
R111_3 core_l3_dff_s_4 core_l3_dff_s_2 0.001
R111_4 core_l3_dff_s core_l3_dff_s_9 180
R111_5 core_l3_dff_s_11 core_l3_dff_s_8 50.4
R111_6 core_l3_dff_s_11 core_l3_dff_s_9 43.2
R111_7 core_l3_dff_s_10 core_l3_dff_s_12 43.2
R111_8 core_l3_dff_s_12 core_l3_dff_s_11 28.8
R111_9 core_l3_dff_s_5 core_l3_dff_s_3 0.54
R111_10 core_l3_dff_s_5 core_l3_dff_s_4 0.648
R111_11 core_l3_dff_s_6 core_l3_dff_s_5 0.54

C4988 core_l3_dff_s vss 1.97571e-16
C4989 core_l3_dff_s_9 vss 1.97571e-16
C4990 core_l3_dff_s_11 vss 5.47722e-17
C4991 core_l3_dff_s_8 vss 5.47722e-17
C4992 core_l3_dff_s_11 vss 4.69476e-17
C4993 core_l3_dff_s_9 vss 4.69476e-17
C4994 core_l3_dff_s_10 vss 4.69476e-17
C4995 core_l3_dff_s_12 vss 4.69476e-17
C4996 core_l3_dff_s_12 vss 3.12984e-17
C4997 core_l3_dff_s_11 vss 3.12984e-17
C4998 core_l3_dff_s_5 vss 5.43283e-17
C4999 core_l3_dff_s_3 vss 5.43283e-17
C5000 core_l3_dff_s_5 vss 7.47014e-17
C5001 core_l3_dff_s_4 vss 7.47014e-17
C5002 core_l3_dff_s_6 vss 5.43283e-17
C5003 core_l3_dff_s_5 vss 5.43283e-17

R112_1 n3245 n3245_5 0.001
R112_2 n3245_3 n3245_2 0.001
R112_3 n3245_4 n3245_2 0.001
R112_4 n3245_4 n3245_3 0.108
R112_5 n3245_5 n3245_4 1.08

C5004 n3245_4 vss 3.10651e-17
C5005 n3245_3 vss 3.10651e-17
C5006 n3245_5 vss 1.18843e-16
C5007 n3245_4 vss 1.18843e-16

R113_1 n3252 n3252_5 0.001
R113_2 n3252_4 n3252_2 0.001
R113_3 n3252_3 n3252_2 0.001
R113_4 n3252_4 n3252_3 0.108
R113_5 n3252_5 n3252_4 1.188

C5008 n3252_4 vss 2.92378e-17
C5009 n3252_3 vss 2.92378e-17
C5010 n3252_5 vss 1.22239e-16
C5011 n3252_4 vss 1.22239e-16

R114_1 core_l3_dff_m core_l3_dff_m_12 0.001
R114_2 core_l3_dff_m_7 core_l3_dff_m_2 0.001
R114_3 core_l3_dff_m_6 core_l3_dff_m_4 0.001
R114_4 core_l3_dff_m_4 core_l3_dff_m_3 64.8
R114_5 core_l3_dff_m_5 core_l3_dff_m_4 93.6
R114_6 core_l3_dff_m_8 core_l3_dff_m_6 0.648
R114_7 core_l3_dff_m_8 core_l3_dff_m_7 0.216
R114_8 core_l3_dff_m_9 core_l3_dff_m_8 0.108
R114_9 core_l3_dff_m_10 core_l3_dff_m_9 0.648
R114_10 core_l3_dff_m_10 core_l3_dff_m_11 0.108
R114_11 core_l3_dff_m_12 core_l3_dff_m_11 0.216

C5012 core_l3_dff_m_4 vss 7.04214e-17
C5013 core_l3_dff_m_3 vss 7.04214e-17
C5014 core_l3_dff_m_5 vss 1.0172e-16
C5015 core_l3_dff_m_4 vss 1.0172e-16
C5016 core_l3_dff_m_8 vss 6.79104e-17
C5017 core_l3_dff_m_6 vss 6.79104e-17
C5018 core_l3_dff_m_8 vss 2.71642e-17
C5019 core_l3_dff_m_7 vss 2.71642e-17
C5020 core_l3_dff_m_9 vss 1.35821e-17
C5021 core_l3_dff_m_8 vss 1.35821e-17
C5022 core_l3_dff_m_10 vss 6.79104e-17
C5023 core_l3_dff_m_9 vss 6.79104e-17
C5024 core_l3_dff_m_10 vss 1.35821e-17
C5025 core_l3_dff_m_11 vss 1.35821e-17
C5026 core_l3_dff_m_12 vss 2.71642e-17
C5027 core_l3_dff_m_11 vss 2.71642e-17

R115_1 n3282 n3282_18 0.001
R115_2 n3282_17 n3282_7 0.001
R115_3 n3282_12 n3282_9 0.001
R115_4 n3282_15 n3282_14 0.001
R115_5 n3282_13 n3282_11 0.001
R115_6 n3282_6 n3282_4 0.001
R115_7 n3282_3 n3282_2 0.001
R115_8 n3282_10 n3282_9 43.2
R115_9 n3282_12 n3282_11 0.54
R115_10 n3282_6 n3282_5 36
R115_11 n3282_4 n3282_3 0.108
R115_12 n3282_14 n3282_13 57.6
R115_13 n3282_7 n3282_6 93.6
R115_14 n3282_16 n3282_15 0.54
R115_15 n3282_8 n3282_7 86.4
R115_16 n3282_17 n3282_16 0.972
R115_17 n3282_18 n3282_17 0.216

C5028 n3282_10 vss 5.086e-17
C5029 n3282_9 vss 5.086e-17
C5030 n3282_12 vss 5.43283e-17
C5031 n3282_11 vss 5.43283e-17
C5032 n3282_6 vss 3.9123e-17
C5033 n3282_5 vss 3.9123e-17
C5034 n3282_4 vss 2.92378e-17
C5035 n3282_3 vss 2.92378e-17
C5036 n3282_14 vss 6.25968e-17
C5037 n3282_13 vss 6.25968e-17
C5038 n3282_7 vss 1.0172e-16
C5039 n3282_6 vss 1.0172e-16
C5040 n3282_16 vss 5.43283e-17
C5041 n3282_15 vss 5.43283e-17
C5042 n3282_8 vss 9.97636e-17
C5043 n3282_7 vss 9.97636e-17
C5044 n3282_17 vss 1.00168e-16
C5045 n3282_16 vss 1.00168e-16
C5046 n3282_18 vss 2.71642e-17
C5047 n3282_17 vss 2.71642e-17

R116_1 core_int_5 core_int_5_7 0.001
R116_2 core_int_5_4 core_int_5_2 0.001
R116_3 core_int_5_5 core_int_5_13 0.001
R116_4 core_int_5_3 core_int_5_2 0.001
R116_5 core_int_5_9 core_int_5_22 0.001
R116_6 core_int_5_10 core_int_5_8 0.001
R116_7 core_int_5_26 core_int_5_16 0.001
R116_8 core_int_5_19 core_int_5_30 0.001
R116_9 core_int_5_29 core_int_5_24 0.001
R116_10 core_int_5_16 core_int_5_15 115.2
R116_11 core_int_5_17 core_int_5_16 43.2
R116_12 core_int_5_26 core_int_5_27 0.108
R116_13 core_int_5_24 core_int_5_23 115.2
R116_14 core_int_5_25 core_int_5_24 64.8
R116_15 core_int_5_27 core_int_5_28 1.62
R116_16 core_int_5_29 core_int_5_28 0.216
R116_17 core_int_5_30 core_int_5_29 0.216
R116_18 core_int_5_19 core_int_5_18 0.81
R116_19 core_int_5_20 core_int_5_19 0.324
R116_20 core_int_5_21 core_int_5_20 0.054
R116_21 core_int_5_22 core_int_5_21 0.81
R116_22 core_int_5_9 core_int_5_8 1.62
R116_23 core_int_5_11 core_int_5_10 0.27
R116_24 core_int_5_12 core_int_5_11 0.054
R116_25 core_int_5_13 core_int_5_12 0.594
R116_26 core_int_5_14 core_int_5_13 0.54
R116_27 core_int_5_4 core_int_5_3 0.216
R116_28 core_int_5_5 core_int_5_4 0.216
R116_29 core_int_5_6 core_int_5_5 0.108
R116_30 core_int_5_7 core_int_5_6 0.324

C5048 core_int_5_16 vss 1.25194e-16
C5049 core_int_5_15 vss 1.25194e-16
C5050 core_int_5_17 vss 5.086e-17
C5051 core_int_5_16 vss 5.086e-17
C5052 core_int_5_26 vss 2.92378e-17
C5053 core_int_5_27 vss 2.92378e-17
C5054 core_int_5_24 vss 1.25194e-16
C5055 core_int_5_23 vss 1.25194e-16
C5056 core_int_5_25 vss 7.43336e-17
C5057 core_int_5_24 vss 7.43336e-17
C5058 core_int_5_27 vss 1.69776e-16
C5059 core_int_5_28 vss 1.69776e-16
C5060 core_int_5_29 vss 2.71642e-17
C5061 core_int_5_28 vss 2.71642e-17
C5062 core_int_5_30 vss 4.38566e-17
C5063 core_int_5_29 vss 4.38566e-17
C5064 core_int_5_19 vss 1.8468e-16
C5065 core_int_5_18 vss 1.8468e-16
C5066 core_int_5_20 vss 7.3872e-17
C5067 core_int_5_19 vss 7.3872e-17
C5068 core_int_5_21 vss 1.2312e-17
C5069 core_int_5_20 vss 1.2312e-17
C5070 core_int_5_22 vss 1.8468e-16
C5071 core_int_5_21 vss 1.8468e-16
C5072 core_int_5_9 vss 1.62985e-16
C5073 core_int_5_8 vss 1.62985e-16
C5074 core_int_5_11 vss 6.156e-17
C5075 core_int_5_10 vss 6.156e-17
C5076 core_int_5_12 vss 1.2312e-17
C5077 core_int_5_11 vss 1.2312e-17
C5078 core_int_5_13 vss 1.35432e-16
C5079 core_int_5_12 vss 1.35432e-16
C5080 core_int_5_14 vss 1.2312e-16
C5081 core_int_5_13 vss 1.2312e-16
C5082 core_int_5_4 vss 4.38566e-17
C5083 core_int_5_3 vss 4.38566e-17
C5084 core_int_5_5 vss 4.38566e-17
C5085 core_int_5_4 vss 4.38566e-17
C5086 core_int_5_6 vss 3.65472e-17
C5087 core_int_5_5 vss 3.65472e-17
C5088 core_int_5_7 vss 4.07462e-17
C5089 core_int_5_6 vss 4.07462e-17

R117_1 bb_2_2 bb_2_6 0.001
R117_2 bb_2_4 bb_2_44 0.001
R117_3 bb_2_41 bb_2_8 0.001
R117_4 bb_2_7 bb_2_11 0.001
R117_5 bb_2_9 bb_2_20 0.001
R117_6 bb_2_19 bb_2_16 0.001
R117_7 bb_2_18 bb_2_24 0.001
R117_8 bb_2_38 bb_2_25 0.001
R117_9 bb_2_26 bb_2_29 0.001
R117_10 bb_2_32 bb_2_49 0.001
R117_11 bb_2_33 bb_2_31 0.001
R117_12 bb_2_47 bb_2_71 0.001
R117_13 bb_2_67 bb_2_50 0.001
R117_14 bb_2_68 bb_2_50 0.001
R117_15 bb_2_70 bb_2_50 0.001
R117_16 bb_2_69 bb_2_50 0.001
R117_17 bb_2_60 bb_2_51 0.001
R117_18 bb_2_59 bb_2_51 0.001
R117_19 bb_2_58 bb_2_51 0.001
R117_20 bb_2_53 bb_2_51 0.001
R117_21 bb_2_54 bb_2_51 0.001
R117_22 bb_2_55 bb_2_51 0.001
R117_23 bb_2_56 bb_2_51 0.001
R117_24 bb_2_57 bb_2_51 0.001
R117_25 bb_2_65 bb_2_51 0.001
R117_26 bb_2_66 bb_2_51 0.001
R117_27 bb_2_61 bb_2_51 0.001
R117_28 bb_2_62 bb_2_51 0.001
R117_29 bb_2_64 bb_2_51 0.001
R117_30 bb_2_63 bb_2_51 0.001
R117_31 bb_2_23 bb_2_21 115.2
R117_32 bb_2_22 bb_2_23 64.8
R117_33 bb_2_24 bb_2_23 7.2
R117_34 bb_2_17 bb_2_14 115.2
R117_35 bb_2_15 bb_2_17 43.2
R117_36 bb_2_53 bb_2_52 0.001
R117_37 bb_2_54 bb_2_53 0.108
R117_38 bb_2_55 bb_2_54 0.108
R117_39 bb_2_56 bb_2_55 0.108
R117_40 bb_2_57 bb_2_56 0.108
R117_41 bb_2_58 bb_2_57 0.108
R117_42 bb_2_59 bb_2_58 0.108
R117_43 bb_2_60 bb_2_59 0.108
R117_44 bb_2_61 bb_2_60 0.108
R117_45 bb_2_62 bb_2_61 0.108
R117_46 bb_2_63 bb_2_62 0.108
R117_47 bb_2_64 bb_2_63 0.108
R117_48 bb_2_65 bb_2_64 0.108
R117_49 bb_2_66 bb_2_65 0.108
R117_50 bb_2_67 bb_2_66 0.864
R117_51 bb_2_68 bb_2_67 0.108
R117_52 bb_2_69 bb_2_68 0.108
R117_53 bb_2_70 bb_2_69 0.108
R117_54 bb_2_71 bb_2_70 0.54
R117_55 bb_2_72 bb_2_71 0.001
R117_56 bb_2_17 bb_2_16 7.2
R117_57 bb_2_19 bb_2_18 0.756
R117_58 bb_2_47 bb_2_46 0.001
R117_59 bb_2_20 bb_2_19 0.108
R117_60 bb_2_48 bb_2_47 0.054
R117_61 bb_2_49 bb_2_48 5.832
R117_62 bb_2_30 bb_2_27 72
R117_63 bb_2_28 bb_2_30 50.4
R117_64 bb_2_9 bb_2_13 0.702
R117_65 bb_2_10 bb_2_9 0.378
R117_66 bb_2_32 bb_2_31 19.548
R117_67 bb_2_30 bb_2_29 7.2
R117_68 bb_2_12 bb_2_11 0.648
R117_69 bb_2_13 bb_2_12 0.054
R117_70 bb_2_34 bb_2_33 0.486
R117_71 bb_2_26 bb_2_25 0.324
R117_72 bb_2_8 bb_2_7 1.944
R117_73 bb_2_35 bb_2_34 0.054
R117_74 bb_2_36 bb_2_35 0.378
R117_75 bb_2_37 bb_2_36 0.054
R117_76 bb_2_38 bb_2_37 0.432
R117_77 bb_2_39 bb_2_38 0.594
R117_78 bb_2_40 bb_2_39 0.054
R117_79 bb_2_41 bb_2_40 0.378
R117_80 bb_2_42 bb_2_41 0.648
R117_81 bb_2_43 bb_2_42 0.054
R117_82 bb_2_44 bb_2_43 0.432
R117_83 bb_2_45 bb_2_44 0.702
R117_84 bb_2_4 bb_2_5 0.216
R117_85 bb_2_6 bb_2_5 0.216
R117_86 bb_2_2 bb_2_1 72
R117_87 bb_2 bb_2_2 50.4

C5090 bb_2_23 vss 1.25194e-16
C5091 bb_2_21 vss 1.25194e-16
C5092 bb_2_22 vss 7.43336e-17
C5093 bb_2_23 vss 7.43336e-17
C5094 bb_2_24 vss 3.15414e-17
C5095 bb_2_23 vss 3.15414e-17
C5096 bb_2_17 vss 1.25194e-16
C5097 bb_2_14 vss 1.25194e-16
C5098 bb_2_15 vss 5.086e-17
C5099 bb_2_17 vss 5.086e-17
C5100 bb_2_53 vss 1.40901e-17
C5101 bb_2_52 vss 1.40901e-17
C5102 bb_2_54 vss 3.13114e-17
C5103 bb_2_53 vss 3.13114e-17
C5104 bb_2_55 vss 3.13114e-17
C5105 bb_2_54 vss 3.13114e-17
C5106 bb_2_56 vss 3.13114e-17
C5107 bb_2_55 vss 3.13114e-17
C5108 bb_2_57 vss 3.13114e-17
C5109 bb_2_56 vss 3.13114e-17
C5110 bb_2_58 vss 3.13114e-17
C5111 bb_2_57 vss 3.13114e-17
C5112 bb_2_59 vss 3.13114e-17
C5113 bb_2_58 vss 3.13114e-17
C5114 bb_2_60 vss 3.13114e-17
C5115 bb_2_59 vss 3.13114e-17
C5116 bb_2_61 vss 3.13114e-17
C5117 bb_2_60 vss 3.13114e-17
C5118 bb_2_62 vss 3.13114e-17
C5119 bb_2_61 vss 3.13114e-17
C5120 bb_2_63 vss 3.13114e-17
C5121 bb_2_62 vss 3.13114e-17
C5122 bb_2_64 vss 3.13114e-17
C5123 bb_2_63 vss 3.13114e-17
C5124 bb_2_65 vss 3.13114e-17
C5125 bb_2_64 vss 3.13114e-17
C5126 bb_2_66 vss 3.13114e-17
C5127 bb_2_65 vss 3.13114e-17
C5128 bb_2_67 vss 2.42663e-16
C5129 bb_2_66 vss 2.42663e-16
C5130 bb_2_68 vss 3.91392e-17
C5131 bb_2_67 vss 3.91392e-17
C5132 bb_2_69 vss 3.91392e-17
C5133 bb_2_68 vss 3.91392e-17
C5134 bb_2_70 vss 3.91392e-17
C5135 bb_2_69 vss 3.91392e-17
C5136 bb_2_71 vss 1.64385e-16
C5137 bb_2_70 vss 1.64385e-16
C5138 bb_2_72 vss 2.1918e-17
C5139 bb_2_71 vss 2.1918e-17
C5140 bb_2_17 vss 3.15414e-17
C5141 bb_2_16 vss 3.15414e-17
C5142 bb_2_19 vss 8.14925e-17
C5143 bb_2_18 vss 8.14925e-17
C5144 bb_2_47 vss 1.30248e-17
C5145 bb_2_46 vss 1.30248e-17
C5146 bb_2_20 vss 3.65472e-17
C5147 bb_2_19 vss 3.65472e-17
C5148 bb_2_48 vss 1.95372e-17
C5149 bb_2_47 vss 1.95372e-17
C5150 bb_2_49 vss 2.11002e-15
C5151 bb_2_48 vss 2.11002e-15
C5152 bb_2_30 vss 8.21582e-17
C5153 bb_2_27 vss 8.21582e-17
C5154 bb_2_28 vss 5.86844e-17
C5155 bb_2_30 vss 5.86844e-17
C5156 bb_2_9 vss 1.66212e-16
C5157 bb_2_13 vss 1.66212e-16
C5158 bb_2_10 vss 9.234e-17
C5159 bb_2_9 vss 9.234e-17
C5160 bb_2_32 vss 1.97619e-15
C5161 bb_2_31 vss 1.97619e-15
C5162 bb_2_30 vss 3.15414e-17
C5163 bb_2_29 vss 3.15414e-17
C5164 bb_2_12 vss 1.539e-16
C5165 bb_2_11 vss 1.539e-16
C5166 bb_2_13 vss 1.2312e-17
C5167 bb_2_12 vss 1.2312e-17
C5168 bb_2_34 vss 1.16964e-16
C5169 bb_2_33 vss 1.16964e-16
C5170 bb_2_26 vss 3.39552e-17
C5171 bb_2_25 vss 3.39552e-17
C5172 bb_2_8 vss 2.03731e-16
C5173 bb_2_7 vss 2.03731e-16
C5174 bb_2_35 vss 1.2312e-17
C5175 bb_2_34 vss 1.2312e-17
C5176 bb_2_36 vss 9.234e-17
C5177 bb_2_35 vss 9.234e-17
C5178 bb_2_37 vss 1.2312e-17
C5179 bb_2_36 vss 1.2312e-17
C5180 bb_2_38 vss 1.04652e-16
C5181 bb_2_37 vss 1.04652e-16
C5182 bb_2_39 vss 1.41588e-16
C5183 bb_2_38 vss 1.41588e-16
C5184 bb_2_40 vss 1.2312e-17
C5185 bb_2_39 vss 1.2312e-17
C5186 bb_2_41 vss 9.234e-17
C5187 bb_2_40 vss 9.234e-17
C5188 bb_2_42 vss 1.539e-16
C5189 bb_2_41 vss 1.539e-16
C5190 bb_2_43 vss 1.2312e-17
C5191 bb_2_42 vss 1.2312e-17
C5192 bb_2_44 vss 9.8496e-17
C5193 bb_2_43 vss 9.8496e-17
C5194 bb_2_45 vss 1.60056e-16
C5195 bb_2_44 vss 1.60056e-16
C5196 bb_2_4 vss 2.54664e-17
C5197 bb_2_5 vss 2.54664e-17
C5198 bb_2_6 vss 2.71642e-17
C5199 bb_2_5 vss 2.71642e-17
C5200 bb_2_2 vss 8.21582e-17
C5201 bb_2_1 vss 8.21582e-17
C5202 bb_2 vss 5.86844e-17
C5203 bb_2_2 vss 5.86844e-17

R118_1 n3407_1 n3407_10 0.001
R118_2 n3407_9 n3407_5 0.001
R118_3 n3407_6 n3407_3 0.001
R118_4 n3407_8 n3407_5 0.001
R118_5 n3407_3 n3407_2 115.2
R118_6 n3407 n3407_3 43.2
R118_7 n3407_6 n3407_7 0.54
R118_8 n3407_9 n3407_7 2.376
R118_9 n3407_9 n3407_8 0.216
R118_10 n3407_11 n3407_9 0.756
R118_11 n3407_11 n3407_10 0.324

C5204 n3407_3 vss 1.25194e-16
C5205 n3407_2 vss 1.25194e-16
C5206 n3407 vss 5.086e-17
C5207 n3407_3 vss 5.086e-17
C5208 n3407_6 vss 5.43283e-17
C5209 n3407_7 vss 5.43283e-17
C5210 n3407_9 vss 2.44477e-16
C5211 n3407_7 vss 2.44477e-16
C5212 n3407_9 vss 3.83746e-17
C5213 n3407_8 vss 3.83746e-17
C5214 n3407_11 vss 8.65858e-17
C5215 n3407_9 vss 8.65858e-17
C5216 n3407_11 vss 4.07462e-17
C5217 n3407_10 vss 4.07462e-17

R119_1 n3422_7 n3422 0.001
R119_2 n3422_3 n3422_11 0.001
R119_3 n3422_6 n3422_5 0.001
R119_4 n3422_8 n3422_6 0.108
R119_5 n3422_9 n3422_7 0.108
R119_6 n3422_10 n3422_8 0.756
R119_7 n3422_9 n3422_10 0.216
R119_8 n3422_12 n3422_10 0.54
R119_9 n3422_12 n3422_11 0.108
R119_10 n3422_3 n3422_2 79.2
R119_11 n3422_4 n3422_3 43.2

C5218 n3422_8 vss 2.19283e-17
C5219 n3422_6 vss 2.19283e-17
C5220 n3422_9 vss 2.92378e-17
C5221 n3422_7 vss 2.92378e-17
C5222 n3422_10 vss 8.14925e-17
C5223 n3422_8 vss 8.14925e-17
C5224 n3422_9 vss 2.71642e-17
C5225 n3422_10 vss 2.71642e-17
C5226 n3422_12 vss 6.11194e-17
C5227 n3422_10 vss 6.11194e-17
C5228 n3422_12 vss 2.19283e-17
C5229 n3422_11 vss 2.19283e-17
C5230 n3422_3 vss 8.9983e-17
C5231 n3422_2 vss 8.9983e-17
C5232 n3422_4 vss 5.086e-17
C5233 n3422_3 vss 5.086e-17

R120_1 core_regout_2_2 core_regout_2_4 0.001
R120_2 core_regout_2_5 core_regout_2_11 0.001
R120_3 core_regout_2_7 core_regout_2_17 0.001
R120_4 core_regout_2_8 core_regout_2_6 0.001
R120_5 core_regout_2_20 core_regout_2_19 0.001
R120_6 core_regout_2_14 core_regout_2_24 0.001
R120_7 core_regout_2_23 core_regout_2_18 0.001
R120_8 core_regout_2_25 core_regout_2_18 0.001
R120_9 core_regout_2_21 core_regout_2_19 0.001
R120_10 core_regout_2_20 core_regout_2_22 0.001
R120_11 core_regout_2_21 core_regout_2_25 0.648
R120_12 core_regout_2_22 core_regout_2_21 0.001
R120_13 core_regout_2_24 core_regout_2_23 0.108
R120_14 core_regout_2_25 core_regout_2_24 0.108
R120_15 core_regout_2_14 core_regout_2_13 0.378
R120_16 core_regout_2_15 core_regout_2_14 0.702
R120_17 core_regout_2_16 core_regout_2_15 0.054
R120_18 core_regout_2_17 core_regout_2_16 0.648
R120_19 core_regout_2_7 core_regout_2_6 9.288
R120_20 core_regout_2_9 core_regout_2_8 0.378
R120_21 core_regout_2_10 core_regout_2_9 0.054
R120_22 core_regout_2_11 core_regout_2_10 0.702
R120_23 core_regout_2_12 core_regout_2_11 0.378
R120_24 core_regout_2_5 core_regout_2_4 0.108
R120_25 core_regout_2_2 core_regout_2_1 72
R120_26 core_regout_2 core_regout_2_2 43.2

C5234 core_regout_2_20 vss 1.60808e-17
C5235 core_regout_2_22 vss 1.60808e-17
C5236 core_regout_2_21 vss 7.47014e-17
C5237 core_regout_2_25 vss 7.47014e-17
C5238 core_regout_2_22 vss 1.3157e-17
C5239 core_regout_2_21 vss 1.3157e-17
C5240 core_regout_2_24 vss 2.19283e-17
C5241 core_regout_2_23 vss 2.19283e-17
C5242 core_regout_2_25 vss 2.19283e-17
C5243 core_regout_2_24 vss 2.19283e-17
C5244 core_regout_2_14 vss 9.234e-17
C5245 core_regout_2_13 vss 9.234e-17
C5246 core_regout_2_15 vss 1.66212e-16
C5247 core_regout_2_14 vss 1.66212e-16
C5248 core_regout_2_16 vss 1.2312e-17
C5249 core_regout_2_15 vss 1.2312e-17
C5250 core_regout_2_17 vss 1.539e-16
C5251 core_regout_2_16 vss 1.539e-16
C5252 core_regout_2_7 vss 9.37163e-16
C5253 core_regout_2_6 vss 9.37163e-16
C5254 core_regout_2_9 vss 9.234e-17
C5255 core_regout_2_8 vss 9.234e-17
C5256 core_regout_2_10 vss 1.2312e-17
C5257 core_regout_2_9 vss 1.2312e-17
C5258 core_regout_2_11 vss 1.66212e-16
C5259 core_regout_2_10 vss 1.66212e-16
C5260 core_regout_2_12 vss 9.234e-17
C5261 core_regout_2_11 vss 9.234e-17
C5262 core_regout_2_5 vss 3.65472e-17
C5263 core_regout_2_4 vss 3.65472e-17
C5264 core_regout_2_2 vss 8.21582e-17
C5265 core_regout_2_1 vss 8.21582e-17
C5266 core_regout_2 vss 5.086e-17
C5267 core_regout_2_2 vss 5.086e-17

R121_1 core_mux_2 core_mux_2_6 0.001
R121_2 core_mux_2_5 core_mux_2_45 0.001
R121_3 core_mux_2_23 core_mux_2_9 0.001
R121_4 core_mux_2_17 core_mux_2_12 0.001
R121_5 core_mux_2_32 core_mux_2_21 0.001
R121_6 core_mux_2_20 core_mux_2_15 0.001
R121_7 core_mux_2_3 core_mux_2_2 0.001
R121_8 core_mux_2_4 core_mux_2_2 0.001
R121_9 core_mux_2_24 core_mux_2_22 0.001
R121_10 core_mux_2_38 core_mux_2_31 0.001
R121_11 core_mux_2_30 core_mux_2_26 0.001
R121_12 core_mux_2_29 core_mux_2_34 0.001
R121_13 core_mux_2_41 core_mux_2_51 0.001
R121_14 core_mux_2_42 core_mux_2_40 0.001
R121_15 core_mux_2_39 core_mux_2_37 0.001
R121_16 core_mux_2_48 core_mux_2_52 0.001
R121_17 core_mux_2_53 core_mux_2_56 0.001
R121_18 core_mux_2_12 core_mux_2_11 115.2
R121_19 core_mux_2_13 core_mux_2_12 43.2
R121_20 core_mux_2_10 core_mux_2_7 72
R121_21 core_mux_2_8 core_mux_2_10 50.4
R121_22 core_mux_2_17 core_mux_2_18 0.108
R121_23 core_mux_2_15 core_mux_2_14 115.2
R121_24 core_mux_2_16 core_mux_2_15 64.8
R121_25 core_mux_2_10 core_mux_2_9 7.2
R121_26 core_mux_2_18 core_mux_2_19 1.62
R121_27 core_mux_2_20 core_mux_2_19 0.216
R121_28 core_mux_2_23 core_mux_2_22 0.324
R121_29 core_mux_2_21 core_mux_2_20 0.216
R121_30 core_mux_2_57 core_mux_2_54 72
R121_31 core_mux_2_55 core_mux_2_57 50.4
R121_32 core_mux_2_57 core_mux_2_56 7.2
R121_33 core_mux_2_24 core_mux_2_28 0.432
R121_34 core_mux_2_25 core_mux_2_24 0.648
R121_35 core_mux_2_32 core_mux_2_36 0.756
R121_36 core_mux_2_33 core_mux_2_32 0.378
R121_37 core_mux_2_27 core_mux_2_26 0.378
R121_38 core_mux_2_28 core_mux_2_27 0.054
R121_39 core_mux_2_35 core_mux_2_34 0.378
R121_40 core_mux_2_36 core_mux_2_35 0.054
R121_41 core_mux_2_53 core_mux_2_52 0.324
R121_42 core_mux_2_30 core_mux_2_29 2.376
R121_43 core_mux_2_31 core_mux_2_30 1.188
R121_44 core_mux_2_48 core_mux_2_47 0.486
R121_45 core_mux_2_49 core_mux_2_48 0.594
R121_46 core_mux_2_50 core_mux_2_49 0.054
R121_47 core_mux_2_51 core_mux_2_50 0.378
R121_48 core_mux_2_38 core_mux_2_37 0.27
R121_49 core_mux_2_40 core_mux_2_39 0.324
R121_50 core_mux_2_41 core_mux_2_40 0.756
R121_51 core_mux_2_43 core_mux_2_42 0.648
R121_52 core_mux_2_44 core_mux_2_43 0.054
R121_53 core_mux_2_45 core_mux_2_44 0.648
R121_54 core_mux_2_46 core_mux_2_45 0.486
R121_55 core_mux_2_4 core_mux_2_3 0.216
R121_56 core_mux_2_5 core_mux_2_4 0.324
R121_57 core_mux_2_6 core_mux_2_5 0.216

C5268 core_mux_2_12 vss 1.25194e-16
C5269 core_mux_2_11 vss 1.25194e-16
C5270 core_mux_2_13 vss 5.086e-17
C5271 core_mux_2_12 vss 5.086e-17
C5272 core_mux_2_10 vss 8.21582e-17
C5273 core_mux_2_7 vss 8.21582e-17
C5274 core_mux_2_8 vss 5.86844e-17
C5275 core_mux_2_10 vss 5.86844e-17
C5276 core_mux_2_17 vss 2.92378e-17
C5277 core_mux_2_18 vss 2.92378e-17
C5278 core_mux_2_15 vss 1.25194e-16
C5279 core_mux_2_14 vss 1.25194e-16
C5280 core_mux_2_16 vss 7.43336e-17
C5281 core_mux_2_15 vss 7.43336e-17
C5282 core_mux_2_10 vss 3.15414e-17
C5283 core_mux_2_9 vss 3.15414e-17
C5284 core_mux_2_18 vss 1.69776e-16
C5285 core_mux_2_19 vss 1.69776e-16
C5286 core_mux_2_20 vss 2.71642e-17
C5287 core_mux_2_19 vss 2.71642e-17
C5288 core_mux_2_23 vss 3.39552e-17
C5289 core_mux_2_22 vss 3.39552e-17
C5290 core_mux_2_21 vss 4.38566e-17
C5291 core_mux_2_20 vss 4.38566e-17
C5292 core_mux_2_57 vss 8.21582e-17
C5293 core_mux_2_54 vss 8.21582e-17
C5294 core_mux_2_55 vss 5.86844e-17
C5295 core_mux_2_57 vss 5.86844e-17
C5296 core_mux_2_57 vss 3.15414e-17
C5297 core_mux_2_56 vss 3.15414e-17
C5298 core_mux_2_24 vss 1.04652e-16
C5299 core_mux_2_28 vss 1.04652e-16
C5300 core_mux_2_25 vss 1.539e-16
C5301 core_mux_2_24 vss 1.539e-16
C5302 core_mux_2_32 vss 1.72368e-16
C5303 core_mux_2_36 vss 1.72368e-16
C5304 core_mux_2_33 vss 8.6184e-17
C5305 core_mux_2_32 vss 8.6184e-17
C5306 core_mux_2_27 vss 9.234e-17
C5307 core_mux_2_26 vss 9.234e-17
C5308 core_mux_2_28 vss 1.2312e-17
C5309 core_mux_2_27 vss 1.2312e-17
C5310 core_mux_2_35 vss 9.234e-17
C5311 core_mux_2_34 vss 9.234e-17
C5312 core_mux_2_36 vss 1.2312e-17
C5313 core_mux_2_35 vss 1.2312e-17
C5314 core_mux_2_53 vss 3.39552e-17
C5315 core_mux_2_52 vss 3.39552e-17
C5316 core_mux_2_30 vss 2.44477e-16
C5317 core_mux_2_29 vss 2.44477e-16
C5318 core_mux_2_31 vss 1.22239e-16
C5319 core_mux_2_30 vss 1.22239e-16
C5320 core_mux_2_48 vss 1.16964e-16
C5321 core_mux_2_47 vss 1.16964e-16
C5322 core_mux_2_49 vss 1.41588e-16
C5323 core_mux_2_48 vss 1.41588e-16
C5324 core_mux_2_50 vss 1.2312e-17
C5325 core_mux_2_49 vss 1.2312e-17
C5326 core_mux_2_51 vss 9.234e-17
C5327 core_mux_2_50 vss 9.234e-17
C5328 core_mux_2_38 vss 6.156e-17
C5329 core_mux_2_37 vss 6.156e-17
C5330 core_mux_2_40 vss 4.07462e-17
C5331 core_mux_2_39 vss 4.07462e-17
C5332 core_mux_2_41 vss 8.14925e-17
C5333 core_mux_2_40 vss 8.14925e-17
C5334 core_mux_2_43 vss 1.539e-16
C5335 core_mux_2_42 vss 1.539e-16
C5336 core_mux_2_44 vss 1.2312e-17
C5337 core_mux_2_43 vss 1.2312e-17
C5338 core_mux_2_45 vss 1.47744e-16
C5339 core_mux_2_44 vss 1.47744e-16
C5340 core_mux_2_46 vss 1.10808e-16
C5341 core_mux_2_45 vss 1.10808e-16
C5342 core_mux_2_4 vss 4.38566e-17
C5343 core_mux_2_3 vss 4.38566e-17
C5344 core_mux_2_5 vss 5.84755e-17
C5345 core_mux_2_4 vss 5.84755e-17
C5346 core_mux_2_6 vss 4.38566e-17
C5347 core_mux_2_5 vss 4.38566e-17

R122_1 core_int_6 core_int_6_6 0.001
R122_2 core_int_6_4 core_int_6_2 0.001
R122_3 core_int_6_5 core_int_6_10 0.001
R122_4 core_int_6_3 core_int_6_2 0.001
R122_5 core_int_6_7 core_int_6_13 0.001
R122_6 core_int_6_12 core_int_6_15 0.001
R122_7 core_int_6_14 core_int_6_17 0.001
R122_8 core_int_6_16 core_int_6_27 0.001
R122_9 core_int_6_24 core_int_6_22 0.001
R122_10 core_int_6_20 core_int_6_18 0.001
R122_11 core_int_6_19 core_int_6_18 136.8
R122_12 core_int_6_20 core_int_6_21 0.108
R122_13 core_int_6_22 core_int_6_21 0.108
R122_14 core_int_6_24 core_int_6_23 0.486
R122_15 core_int_6_25 core_int_6_24 0.648
R122_16 core_int_6_26 core_int_6_25 0.054
R122_17 core_int_6_27 core_int_6_26 0.27
R122_18 core_int_6_17 core_int_6_16 2.376
R122_19 core_int_6_15 core_int_6_14 0.54
R122_20 core_int_6_13 core_int_6_12 1.944
R122_21 core_int_6_8 core_int_6_7 0.27
R122_22 core_int_6_9 core_int_6_8 0.054
R122_23 core_int_6_10 core_int_6_9 0.594
R122_24 core_int_6_11 core_int_6_10 0.486
R122_25 core_int_6_4 core_int_6_3 0.216
R122_26 core_int_6_5 core_int_6_4 0.216
R122_27 core_int_6_6 core_int_6_5 0.216

C5348 core_int_6_19 vss 1.54536e-16
C5349 core_int_6_18 vss 1.54536e-16
C5350 core_int_6_20 vss 2.92378e-17
C5351 core_int_6_21 vss 2.92378e-17
C5352 core_int_6_22 vss 2.92378e-17
C5353 core_int_6_21 vss 2.92378e-17
C5354 core_int_6_24 vss 1.10808e-16
C5355 core_int_6_23 vss 1.10808e-16
C5356 core_int_6_25 vss 1.47744e-16
C5357 core_int_6_24 vss 1.47744e-16
C5358 core_int_6_26 vss 1.2312e-17
C5359 core_int_6_25 vss 1.2312e-17
C5360 core_int_6_27 vss 6.156e-17
C5361 core_int_6_26 vss 6.156e-17
C5362 core_int_6_17 vss 2.44477e-16
C5363 core_int_6_16 vss 2.44477e-16
C5364 core_int_6_15 vss 1.2312e-16
C5365 core_int_6_14 vss 1.2312e-16
C5366 core_int_6_13 vss 2.03731e-16
C5367 core_int_6_12 vss 2.03731e-16
C5368 core_int_6_8 vss 6.156e-17
C5369 core_int_6_7 vss 6.156e-17
C5370 core_int_6_9 vss 1.2312e-17
C5371 core_int_6_8 vss 1.2312e-17
C5372 core_int_6_10 vss 1.41588e-16
C5373 core_int_6_9 vss 1.41588e-16
C5374 core_int_6_11 vss 1.16964e-16
C5375 core_int_6_10 vss 1.16964e-16
C5376 core_int_6_4 vss 4.38566e-17
C5377 core_int_6_3 vss 4.38566e-17
C5378 core_int_6_5 vss 5.11661e-17
C5379 core_int_6_4 vss 5.11661e-17
C5380 core_int_6_6 vss 5.11661e-17
C5381 core_int_6_5 vss 5.11661e-17

R123_1 n3558_1 n3558_11 0.001
R123_2 n3558_7 n3558_5 0.001
R123_3 n3558_9 n3558_6 0.001
R123_4 n3558_4 n3558_2 72
R123_5 n3558 n3558_4 43.2
R123_6 n3558_5 n3558_4 7.2
R123_7 n3558_7 n3558_8 0.108
R123_8 n3558_9 n3558_8 0.756
R123_9 n3558_10 n3558_9 0.324
R123_10 n3558_11 n3558_10 0.648

C5382 n3558_4 vss 8.21582e-17
C5383 n3558_2 vss 8.21582e-17
C5384 n3558 vss 5.086e-17
C5385 n3558_4 vss 5.086e-17
C5386 n3558_5 vss 3.15414e-17
C5387 n3558_4 vss 3.15414e-17
C5388 n3558_7 vss 3.65472e-17
C5389 n3558_8 vss 3.65472e-17
C5390 n3558_9 vss 8.14925e-17
C5391 n3558_8 vss 8.14925e-17
C5392 n3558_10 vss 4.07462e-17
C5393 n3558_9 vss 4.07462e-17
C5394 n3558_11 vss 6.79104e-17
C5395 n3558_10 vss 6.79104e-17

R124_1 core_int_2 core_int_2_6 0.001
R124_2 core_int_2_3 core_int_2_2 0.001
R124_3 core_int_2_4 core_int_2_2 0.001
R124_4 core_int_2_5 core_int_2_10 0.001
R124_5 core_int_2_7 core_int_2_13 0.001
R124_6 core_int_2_12 core_int_2_23 0.001
R124_7 core_int_2_20 core_int_2_18 0.001
R124_8 core_int_2_16 core_int_2_14 0.001
R124_9 core_int_2_15 core_int_2_14 136.8
R124_10 core_int_2_16 core_int_2_17 0.108
R124_11 core_int_2_18 core_int_2_17 0.108
R124_12 core_int_2_20 core_int_2_19 0.486
R124_13 core_int_2_21 core_int_2_20 0.648
R124_14 core_int_2_22 core_int_2_21 0.054
R124_15 core_int_2_23 core_int_2_22 0.27
R124_16 core_int_2_13 core_int_2_12 1.188
R124_17 core_int_2_8 core_int_2_7 0.81
R124_18 core_int_2_9 core_int_2_8 0.054
R124_19 core_int_2_10 core_int_2_9 0.594
R124_20 core_int_2_11 core_int_2_10 0.486
R124_21 core_int_2_4 core_int_2_3 0.216
R124_22 core_int_2_5 core_int_2_4 0.216
R124_23 core_int_2_6 core_int_2_5 0.216

C5396 core_int_2_15 vss 1.54536e-16
C5397 core_int_2_14 vss 1.54536e-16
C5398 core_int_2_16 vss 2.92378e-17
C5399 core_int_2_17 vss 2.92378e-17
C5400 core_int_2_18 vss 2.92378e-17
C5401 core_int_2_17 vss 2.92378e-17
C5402 core_int_2_20 vss 1.10808e-16
C5403 core_int_2_19 vss 1.10808e-16
C5404 core_int_2_21 vss 1.47744e-16
C5405 core_int_2_20 vss 1.47744e-16
C5406 core_int_2_22 vss 1.2312e-17
C5407 core_int_2_21 vss 1.2312e-17
C5408 core_int_2_23 vss 6.156e-17
C5409 core_int_2_22 vss 6.156e-17
C5410 core_int_2_13 vss 1.22239e-16
C5411 core_int_2_12 vss 1.22239e-16
C5412 core_int_2_8 vss 1.8468e-16
C5413 core_int_2_7 vss 1.8468e-16
C5414 core_int_2_9 vss 1.2312e-17
C5415 core_int_2_8 vss 1.2312e-17
C5416 core_int_2_10 vss 1.41588e-16
C5417 core_int_2_9 vss 1.41588e-16
C5418 core_int_2_11 vss 1.16964e-16
C5419 core_int_2_10 vss 1.16964e-16
C5420 core_int_2_4 vss 4.38566e-17
C5421 core_int_2_3 vss 4.38566e-17
C5422 core_int_2_5 vss 5.11661e-17
C5423 core_int_2_4 vss 5.11661e-17
C5424 core_int_2_6 vss 5.11661e-17
C5425 core_int_2_5 vss 5.11661e-17

R125_1 n3595 n3595_11 0.001
R125_2 n3595_6 n3595_3 0.001
R125_3 n3595_7 n3595_5 0.001
R125_4 n3595_3 n3595_2 79.2
R125_5 n3595_4 n3595_3 43.2
R125_6 n3595_8 n3595_6 0.108
R125_7 n3595_9 n3595_7 0.108
R125_8 n3595_8 n3595_10 0.54
R125_9 n3595_10 n3595_9 0.756
R125_10 n3595_12 n3595_10 0.216
R125_11 n3595_12 n3595_11 0.108

C5426 n3595_3 vss 8.9983e-17
C5427 n3595_2 vss 8.9983e-17
C5428 n3595_4 vss 5.086e-17
C5429 n3595_3 vss 5.086e-17
C5430 n3595_8 vss 2.19283e-17
C5431 n3595_6 vss 2.19283e-17
C5432 n3595_9 vss 2.19283e-17
C5433 n3595_7 vss 2.19283e-17
C5434 n3595_8 vss 6.11194e-17
C5435 n3595_10 vss 6.11194e-17
C5436 n3595_10 vss 8.14925e-17
C5437 n3595_9 vss 8.14925e-17
C5438 n3595_12 vss 2.71642e-17
C5439 n3595_10 vss 2.71642e-17
C5440 n3595_12 vss 2.92378e-17
C5441 n3595_11 vss 2.92378e-17

R126_1 bb_1_1 bb_1_10 0.001
R126_2 bb_1_11 bb_1_7 0.001
R126_3 bb_1_9 bb_1_15 0.001
R126_4 bb_1_12 bb_1_30 0.001
R126_5 bb_1_28 bb_1_19 0.001
R126_6 bb_1_29 bb_1_47 0.001
R126_7 bb_1_17 bb_1_27 0.001
R126_8 bb_1_25 bb_1_23 0.001
R126_9 bb_1_44 bb_1_31 0.001
R126_10 bb_1_32 bb_1_35 0.001
R126_11 bb_1_38 bb_1_51 0.001
R126_12 bb_1_39 bb_1_37 0.001
R126_13 bb_1_49 bb_1_55 0.001
R126_14 bb_1_53 bb_1_77 0.001
R126_15 bb_1_74 bb_1_56 0.001
R126_16 bb_1_73 bb_1_56 0.001
R126_17 bb_1_76 bb_1_56 0.001
R126_18 bb_1_75 bb_1_56 0.001
R126_19 bb_1_50 bb_1_48 0.001
R126_20 bb_1_66 bb_1_57 0.001
R126_21 bb_1_65 bb_1_57 0.001
R126_22 bb_1_64 bb_1_57 0.001
R126_23 bb_1_59 bb_1_57 0.001
R126_24 bb_1_60 bb_1_57 0.001
R126_25 bb_1_61 bb_1_57 0.001
R126_26 bb_1_62 bb_1_57 0.001
R126_27 bb_1_63 bb_1_57 0.001
R126_28 bb_1_70 bb_1_57 0.001
R126_29 bb_1_69 bb_1_57 0.001
R126_30 bb_1_71 bb_1_57 0.001
R126_31 bb_1_72 bb_1_57 0.001
R126_32 bb_1_67 bb_1_57 0.001
R126_33 bb_1_68 bb_1_57 0.001
R126_34 bb_1_59 bb_1_58 0.001
R126_35 bb_1_60 bb_1_59 0.108
R126_36 bb_1_61 bb_1_60 0.108
R126_37 bb_1_62 bb_1_61 0.108
R126_38 bb_1_63 bb_1_62 0.108
R126_39 bb_1_64 bb_1_63 0.108
R126_40 bb_1_65 bb_1_64 0.108
R126_41 bb_1_66 bb_1_65 0.108
R126_42 bb_1_67 bb_1_66 0.108
R126_43 bb_1_68 bb_1_67 0.108
R126_44 bb_1_69 bb_1_68 0.108
R126_45 bb_1_70 bb_1_69 0.108
R126_46 bb_1_71 bb_1_70 0.108
R126_47 bb_1_72 bb_1_71 0.108
R126_48 bb_1_73 bb_1_72 0.864
R126_49 bb_1_74 bb_1_73 0.108
R126_50 bb_1_75 bb_1_74 0.108
R126_51 bb_1_76 bb_1_75 0.108
R126_52 bb_1_77 bb_1_76 0.54
R126_53 bb_1_78 bb_1_77 0.001
R126_54 bb_1_53 bb_1_52 0.001
R126_55 bb_1_54 bb_1_53 0.054
R126_56 bb_1_55 bb_1_54 0.162
R126_57 bb_1_49 bb_1_48 3.888
R126_58 bb_1_51 bb_1_50 5.454
R126_59 bb_1_23 bb_1_22 72
R126_60 bb_1_24 bb_1_23 50.4
R126_61 bb_1_36 bb_1_33 72
R126_62 bb_1_34 bb_1_36 50.4
R126_63 bb_1_38 bb_1_37 17.064
R126_64 bb_1_36 bb_1_35 7.2
R126_65 bb_1_25 bb_1_26 0.216
R126_66 bb_1_27 bb_1_26 0.216
R126_67 bb_1_40 bb_1_39 0.756
R126_68 bb_1_32 bb_1_31 0.324
R126_69 bb_1_41 bb_1_40 0.054
R126_70 bb_1_42 bb_1_41 0.378
R126_71 bb_1_43 bb_1_42 0.054
R126_72 bb_1_44 bb_1_43 0.432
R126_73 bb_1_45 bb_1_44 0.594
R126_74 bb_1_17 bb_1_21 0.432
R126_75 bb_1_18 bb_1_17 0.702
R126_76 bb_1_46 bb_1_45 0.054
R126_77 bb_1_47 bb_1_46 0.54
R126_78 bb_1_20 bb_1_19 0.54
R126_79 bb_1_21 bb_1_20 0.054
R126_80 bb_1_29 bb_1_28 2.376
R126_81 bb_1_30 bb_1_29 2.808
R126_82 bb_1_13 bb_1_12 0.54
R126_83 bb_1_14 bb_1_13 0.054
R126_84 bb_1_15 bb_1_14 0.702
R126_85 bb_1_16 bb_1_15 0.378
R126_86 bb_1_8 bb_1_5 115.2
R126_87 bb_1_6 bb_1_8 43.2
R126_88 bb_1_8 bb_1_7 7.2
R126_89 bb_1_9 bb_1_11 0.108
R126_90 bb_1_11 bb_1_10 0.756
R126_91 bb_1_1 bb_1_3 7.2
R126_92 bb_1_3 bb_1_2 115.2
R126_93 bb_1 bb_1_3 64.8

C5442 bb_1_59 vss 1.40901e-17
C5443 bb_1_58 vss 1.40901e-17
C5444 bb_1_60 vss 3.13114e-17
C5445 bb_1_59 vss 3.13114e-17
C5446 bb_1_61 vss 3.13114e-17
C5447 bb_1_60 vss 3.13114e-17
C5448 bb_1_62 vss 3.13114e-17
C5449 bb_1_61 vss 3.13114e-17
C5450 bb_1_63 vss 3.13114e-17
C5451 bb_1_62 vss 3.13114e-17
C5452 bb_1_64 vss 3.13114e-17
C5453 bb_1_63 vss 3.13114e-17
C5454 bb_1_65 vss 3.13114e-17
C5455 bb_1_64 vss 3.13114e-17
C5456 bb_1_66 vss 3.13114e-17
C5457 bb_1_65 vss 3.13114e-17
C5458 bb_1_67 vss 3.13114e-17
C5459 bb_1_66 vss 3.13114e-17
C5460 bb_1_68 vss 3.13114e-17
C5461 bb_1_67 vss 3.13114e-17
C5462 bb_1_69 vss 3.13114e-17
C5463 bb_1_68 vss 3.13114e-17
C5464 bb_1_70 vss 3.13114e-17
C5465 bb_1_69 vss 3.13114e-17
C5466 bb_1_71 vss 3.13114e-17
C5467 bb_1_70 vss 3.13114e-17
C5468 bb_1_72 vss 3.13114e-17
C5469 bb_1_71 vss 3.13114e-17
C5470 bb_1_73 vss 2.42663e-16
C5471 bb_1_72 vss 2.42663e-16
C5472 bb_1_74 vss 3.91392e-17
C5473 bb_1_73 vss 3.91392e-17
C5474 bb_1_75 vss 3.91392e-17
C5475 bb_1_74 vss 3.91392e-17
C5476 bb_1_76 vss 3.91392e-17
C5477 bb_1_75 vss 3.91392e-17
C5478 bb_1_77 vss 1.64385e-16
C5479 bb_1_76 vss 1.64385e-16
C5480 bb_1_78 vss 2.1918e-17
C5481 bb_1_77 vss 2.1918e-17
C5482 bb_1_53 vss 1.30248e-17
C5483 bb_1_52 vss 1.30248e-17
C5484 bb_1_54 vss 1.95372e-17
C5485 bb_1_53 vss 1.95372e-17
C5486 bb_1_55 vss 5.86116e-17
C5487 bb_1_54 vss 5.86116e-17
C5488 bb_1_49 vss 7.01706e-16
C5489 bb_1_48 vss 7.01706e-16
C5490 bb_1_51 vss 1.98629e-15
C5491 bb_1_50 vss 1.98629e-15
C5492 bb_1_23 vss 8.21582e-17
C5493 bb_1_22 vss 8.21582e-17
C5494 bb_1_24 vss 5.86844e-17
C5495 bb_1_23 vss 5.86844e-17
C5496 bb_1_36 vss 8.21582e-17
C5497 bb_1_33 vss 8.21582e-17
C5498 bb_1_34 vss 5.86844e-17
C5499 bb_1_36 vss 5.86844e-17
C5500 bb_1_38 vss 1.71813e-15
C5501 bb_1_37 vss 1.71813e-15
C5502 bb_1_36 vss 3.15414e-17
C5503 bb_1_35 vss 3.15414e-17
C5504 bb_1_25 vss 2.71642e-17
C5505 bb_1_26 vss 2.71642e-17
C5506 bb_1_27 vss 2.54664e-17
C5507 bb_1_26 vss 2.54664e-17
C5508 bb_1_40 vss 1.78524e-16
C5509 bb_1_39 vss 1.78524e-16
C5510 bb_1_32 vss 3.39552e-17
C5511 bb_1_31 vss 3.39552e-17
C5512 bb_1_41 vss 1.2312e-17
C5513 bb_1_40 vss 1.2312e-17
C5514 bb_1_42 vss 9.234e-17
C5515 bb_1_41 vss 9.234e-17
C5516 bb_1_43 vss 1.2312e-17
C5517 bb_1_42 vss 1.2312e-17
C5518 bb_1_44 vss 1.04652e-16
C5519 bb_1_43 vss 1.04652e-16
C5520 bb_1_45 vss 1.41588e-16
C5521 bb_1_44 vss 1.41588e-16
C5522 bb_1_17 vss 9.8496e-17
C5523 bb_1_21 vss 9.8496e-17
C5524 bb_1_18 vss 1.60056e-16
C5525 bb_1_17 vss 1.60056e-16
C5526 bb_1_46 vss 1.2312e-17
C5527 bb_1_45 vss 1.2312e-17
C5528 bb_1_47 vss 1.2312e-16
C5529 bb_1_46 vss 1.2312e-16
C5530 bb_1_20 vss 1.2312e-16
C5531 bb_1_19 vss 1.2312e-16
C5532 bb_1_21 vss 1.2312e-17
C5533 bb_1_20 vss 1.2312e-17
C5534 bb_1_29 vss 2.44477e-16
C5535 bb_1_28 vss 2.44477e-16
C5536 bb_1_30 vss 2.85224e-16
C5537 bb_1_29 vss 2.85224e-16
C5538 bb_1_13 vss 1.2312e-16
C5539 bb_1_12 vss 1.2312e-16
C5540 bb_1_14 vss 1.2312e-17
C5541 bb_1_13 vss 1.2312e-17
C5542 bb_1_15 vss 1.66212e-16
C5543 bb_1_14 vss 1.66212e-16
C5544 bb_1_16 vss 9.234e-17
C5545 bb_1_15 vss 9.234e-17
C5546 bb_1_8 vss 1.25194e-16
C5547 bb_1_5 vss 1.25194e-16
C5548 bb_1_6 vss 5.086e-17
C5549 bb_1_8 vss 5.086e-17
C5550 bb_1_8 vss 3.15414e-17
C5551 bb_1_7 vss 3.15414e-17
C5552 bb_1_9 vss 3.65472e-17
C5553 bb_1_11 vss 3.65472e-17
C5554 bb_1_11 vss 8.14925e-17
C5555 bb_1_10 vss 8.14925e-17
C5556 bb_1_1 vss 3.15414e-17
C5557 bb_1_3 vss 3.15414e-17
C5558 bb_1_3 vss 1.25194e-16
C5559 bb_1_2 vss 1.25194e-16
C5560 bb_1 vss 7.43336e-17
C5561 bb_1_3 vss 7.43336e-17

R127_1 core_mux_1 core_mux_1_6 0.001
R127_2 core_mux_1_4 core_mux_1_2 0.001
R127_3 core_mux_1_5 core_mux_1_27 0.001
R127_4 core_mux_1_13 core_mux_1_8 0.001
R127_5 core_mux_1_43 core_mux_1_17 0.001
R127_6 core_mux_1_16 core_mux_1_11 0.001
R127_7 core_mux_1_32 core_mux_1_18 0.001
R127_8 core_mux_1_19 core_mux_1_22 0.001
R127_9 core_mux_1_3 core_mux_1_2 0.001
R127_10 core_mux_1_24 core_mux_1_31 0.001
R127_11 core_mux_1_30 core_mux_1_49 0.001
R127_12 core_mux_1_29 core_mux_1_34 0.001
R127_13 core_mux_1_46 core_mux_1_37 0.001
R127_14 core_mux_1_38 core_mux_1_41 0.001
R127_15 core_mux_1_8 core_mux_1_7 115.2
R127_16 core_mux_1_9 core_mux_1_8 43.2
R127_17 core_mux_1_13 core_mux_1_14 0.108
R127_18 core_mux_1_11 core_mux_1_10 115.2
R127_19 core_mux_1_12 core_mux_1_11 64.8
R127_20 core_mux_1_42 core_mux_1_39 72
R127_21 core_mux_1_40 core_mux_1_42 50.4
R127_22 core_mux_1_23 core_mux_1_20 72
R127_23 core_mux_1_21 core_mux_1_23 50.4
R127_24 core_mux_1_14 core_mux_1_15 1.62
R127_25 core_mux_1_42 core_mux_1_41 7.2
R127_26 core_mux_1_23 core_mux_1_22 7.2
R127_27 core_mux_1_16 core_mux_1_15 0.216
R127_28 core_mux_1_17 core_mux_1_16 0.216
R127_29 core_mux_1_38 core_mux_1_37 0.324
R127_30 core_mux_1_19 core_mux_1_18 0.324
R127_31 core_mux_1_43 core_mux_1_51 0.756
R127_32 core_mux_1_44 core_mux_1_43 0.378
R127_33 core_mux_1_46 core_mux_1_45 0.486
R127_34 core_mux_1_47 core_mux_1_46 0.594
R127_35 core_mux_1_32 core_mux_1_36 0.432
R127_36 core_mux_1_33 core_mux_1_32 0.648
R127_37 core_mux_1_48 core_mux_1_47 0.054
R127_38 core_mux_1_49 core_mux_1_48 0.81
R127_39 core_mux_1_50 core_mux_1_49 0.27
R127_40 core_mux_1_51 core_mux_1_50 0.054
R127_41 core_mux_1_35 core_mux_1_34 0.27
R127_42 core_mux_1_36 core_mux_1_35 0.054
R127_43 core_mux_1_30 core_mux_1_29 4.86
R127_44 core_mux_1_31 core_mux_1_30 2.376
R127_45 core_mux_1_25 core_mux_1_24 0.27
R127_46 core_mux_1_26 core_mux_1_25 0.054
R127_47 core_mux_1_27 core_mux_1_26 0.648
R127_48 core_mux_1_28 core_mux_1_27 0.486
R127_49 core_mux_1_4 core_mux_1_3 0.216
R127_50 core_mux_1_5 core_mux_1_4 0.324
R127_51 core_mux_1_6 core_mux_1_5 0.216

C5562 core_mux_1_8 vss 1.25194e-16
C5563 core_mux_1_7 vss 1.25194e-16
C5564 core_mux_1_9 vss 5.086e-17
C5565 core_mux_1_8 vss 5.086e-17
C5566 core_mux_1_13 vss 2.92378e-17
C5567 core_mux_1_14 vss 2.92378e-17
C5568 core_mux_1_11 vss 1.25194e-16
C5569 core_mux_1_10 vss 1.25194e-16
C5570 core_mux_1_12 vss 7.43336e-17
C5571 core_mux_1_11 vss 7.43336e-17
C5572 core_mux_1_42 vss 8.21582e-17
C5573 core_mux_1_39 vss 8.21582e-17
C5574 core_mux_1_40 vss 5.86844e-17
C5575 core_mux_1_42 vss 5.86844e-17
C5576 core_mux_1_23 vss 8.21582e-17
C5577 core_mux_1_20 vss 8.21582e-17
C5578 core_mux_1_21 vss 5.86844e-17
C5579 core_mux_1_23 vss 5.86844e-17
C5580 core_mux_1_14 vss 1.69776e-16
C5581 core_mux_1_15 vss 1.69776e-16
C5582 core_mux_1_42 vss 3.15414e-17
C5583 core_mux_1_41 vss 3.15414e-17
C5584 core_mux_1_23 vss 3.15414e-17
C5585 core_mux_1_22 vss 3.15414e-17
C5586 core_mux_1_16 vss 2.71642e-17
C5587 core_mux_1_15 vss 2.71642e-17
C5588 core_mux_1_17 vss 4.38566e-17
C5589 core_mux_1_16 vss 4.38566e-17
C5590 core_mux_1_38 vss 3.39552e-17
C5591 core_mux_1_37 vss 3.39552e-17
C5592 core_mux_1_19 vss 3.39552e-17
C5593 core_mux_1_18 vss 3.39552e-17
C5594 core_mux_1_43 vss 1.72368e-16
C5595 core_mux_1_51 vss 1.72368e-16
C5596 core_mux_1_44 vss 8.6184e-17
C5597 core_mux_1_43 vss 8.6184e-17
C5598 core_mux_1_46 vss 1.16964e-16
C5599 core_mux_1_45 vss 1.16964e-16
C5600 core_mux_1_47 vss 1.41588e-16
C5601 core_mux_1_46 vss 1.41588e-16
C5602 core_mux_1_32 vss 1.04652e-16
C5603 core_mux_1_36 vss 1.04652e-16
C5604 core_mux_1_33 vss 1.539e-16
C5605 core_mux_1_32 vss 1.539e-16
C5606 core_mux_1_48 vss 1.2312e-17
C5607 core_mux_1_47 vss 1.2312e-17
C5608 core_mux_1_49 vss 1.8468e-16
C5609 core_mux_1_48 vss 1.8468e-16
C5610 core_mux_1_50 vss 6.156e-17
C5611 core_mux_1_49 vss 6.156e-17
C5612 core_mux_1_51 vss 1.2312e-17
C5613 core_mux_1_50 vss 1.2312e-17
C5614 core_mux_1_35 vss 6.156e-17
C5615 core_mux_1_34 vss 6.156e-17
C5616 core_mux_1_36 vss 1.2312e-17
C5617 core_mux_1_35 vss 1.2312e-17
C5618 core_mux_1_30 vss 4.88955e-16
C5619 core_mux_1_29 vss 4.88955e-16
C5620 core_mux_1_31 vss 2.44477e-16
C5621 core_mux_1_30 vss 2.44477e-16
C5622 core_mux_1_25 vss 6.156e-17
C5623 core_mux_1_24 vss 6.156e-17
C5624 core_mux_1_26 vss 1.2312e-17
C5625 core_mux_1_25 vss 1.2312e-17
C5626 core_mux_1_27 vss 1.47744e-16
C5627 core_mux_1_26 vss 1.47744e-16
C5628 core_mux_1_28 vss 1.10808e-16
C5629 core_mux_1_27 vss 1.10808e-16
C5630 core_mux_1_4 vss 4.38566e-17
C5631 core_mux_1_3 vss 4.38566e-17
C5632 core_mux_1_5 vss 5.84755e-17
C5633 core_mux_1_4 vss 5.84755e-17
C5634 core_mux_1_6 vss 4.38566e-17
C5635 core_mux_1_5 vss 4.38566e-17

R128_1 n3746_1 n3746_10 0.001
R128_2 n3746_9 n3746_5 0.001
R128_3 n3746_6 n3746_3 0.001
R128_4 n3746_8 n3746_5 0.001
R128_5 n3746_3 n3746_2 115.2
R128_6 n3746 n3746_3 43.2
R128_7 n3746_6 n3746_7 0.54
R128_8 n3746_9 n3746_7 2.376
R128_9 n3746_9 n3746_8 0.216
R128_10 n3746_11 n3746_9 0.756
R128_11 n3746_11 n3746_10 0.324

C5636 n3746_3 vss 1.25194e-16
C5637 n3746_2 vss 1.25194e-16
C5638 n3746 vss 5.086e-17
C5639 n3746_3 vss 5.086e-17
C5640 n3746_6 vss 5.43283e-17
C5641 n3746_7 vss 5.43283e-17
C5642 n3746_9 vss 2.44477e-16
C5643 n3746_7 vss 2.44477e-16
C5644 n3746_9 vss 3.83746e-17
C5645 n3746_8 vss 3.83746e-17
C5646 n3746_11 vss 8.65858e-17
C5647 n3746_9 vss 8.65858e-17
C5648 n3746_11 vss 4.07462e-17
C5649 n3746_10 vss 4.07462e-17

R129_1 core_mux_0 core_mux_0_6 0.001
R129_2 core_mux_0_4 core_mux_0_2 0.001
R129_3 core_mux_0_5 core_mux_0_12 0.001
R129_4 core_mux_0_3 core_mux_0_2 0.001
R129_5 core_mux_0_8 core_mux_0_27 0.001
R129_6 core_mux_0_9 core_mux_0_7 0.001
R129_7 core_mux_0_15 core_mux_0_35 0.001
R129_8 core_mux_0_26 core_mux_0_14 0.001
R129_9 core_mux_0_39 core_mux_0_29 0.001
R129_10 core_mux_0_32 core_mux_0_43 0.001
R129_11 core_mux_0_42 core_mux_0_37 0.001
R129_12 core_mux_0_23 core_mux_0_16 0.001
R129_13 core_mux_0_17 core_mux_0_20 0.001
R129_14 core_mux_0_29 core_mux_0_28 115.2
R129_15 core_mux_0_30 core_mux_0_29 43.2
R129_16 core_mux_0_39 core_mux_0_40 0.108
R129_17 core_mux_0_37 core_mux_0_36 115.2
R129_18 core_mux_0_38 core_mux_0_37 64.8
R129_19 core_mux_0_40 core_mux_0_41 1.62
R129_20 core_mux_0_42 core_mux_0_41 0.216
R129_21 core_mux_0_43 core_mux_0_42 0.216
R129_22 core_mux_0_21 core_mux_0_18 72
R129_23 core_mux_0_19 core_mux_0_21 50.4
R129_24 core_mux_0_32 core_mux_0_31 0.81
R129_25 core_mux_0_33 core_mux_0_32 0.324
R129_26 core_mux_0_21 core_mux_0_20 7.2
R129_27 core_mux_0_34 core_mux_0_33 0.054
R129_28 core_mux_0_35 core_mux_0_34 0.378
R129_29 core_mux_0_17 core_mux_0_16 0.324
R129_30 core_mux_0_15 core_mux_0_14 2.376
R129_31 core_mux_0_23 core_mux_0_22 0.486
R129_32 core_mux_0_24 core_mux_0_23 0.594
R129_33 core_mux_0_25 core_mux_0_24 0.054
R129_34 core_mux_0_26 core_mux_0_25 0.378
R129_35 core_mux_0_27 core_mux_0_26 0.378
R129_36 core_mux_0_8 core_mux_0_7 1.188
R129_37 core_mux_0_10 core_mux_0_9 0.27
R129_38 core_mux_0_11 core_mux_0_10 0.054
R129_39 core_mux_0_12 core_mux_0_11 0.648
R129_40 core_mux_0_13 core_mux_0_12 0.486
R129_41 core_mux_0_4 core_mux_0_3 0.216
R129_42 core_mux_0_5 core_mux_0_4 0.324
R129_43 core_mux_0_6 core_mux_0_5 0.216

C5650 core_mux_0_29 vss 1.25194e-16
C5651 core_mux_0_28 vss 1.25194e-16
C5652 core_mux_0_30 vss 5.086e-17
C5653 core_mux_0_29 vss 5.086e-17
C5654 core_mux_0_39 vss 2.92378e-17
C5655 core_mux_0_40 vss 2.92378e-17
C5656 core_mux_0_37 vss 1.25194e-16
C5657 core_mux_0_36 vss 1.25194e-16
C5658 core_mux_0_38 vss 7.43336e-17
C5659 core_mux_0_37 vss 7.43336e-17
C5660 core_mux_0_40 vss 1.69776e-16
C5661 core_mux_0_41 vss 1.69776e-16
C5662 core_mux_0_42 vss 2.71642e-17
C5663 core_mux_0_41 vss 2.71642e-17
C5664 core_mux_0_43 vss 4.38566e-17
C5665 core_mux_0_42 vss 4.38566e-17
C5666 core_mux_0_21 vss 8.21582e-17
C5667 core_mux_0_18 vss 8.21582e-17
C5668 core_mux_0_19 vss 5.86844e-17
C5669 core_mux_0_21 vss 5.86844e-17
C5670 core_mux_0_32 vss 1.8468e-16
C5671 core_mux_0_31 vss 1.8468e-16
C5672 core_mux_0_33 vss 7.3872e-17
C5673 core_mux_0_32 vss 7.3872e-17
C5674 core_mux_0_21 vss 3.15414e-17
C5675 core_mux_0_20 vss 3.15414e-17
C5676 core_mux_0_34 vss 1.2312e-17
C5677 core_mux_0_33 vss 1.2312e-17
C5678 core_mux_0_35 vss 9.234e-17
C5679 core_mux_0_34 vss 9.234e-17
C5680 core_mux_0_17 vss 3.39552e-17
C5681 core_mux_0_16 vss 3.39552e-17
C5682 core_mux_0_15 vss 2.44477e-16
C5683 core_mux_0_14 vss 2.44477e-16
C5684 core_mux_0_23 vss 1.16964e-16
C5685 core_mux_0_22 vss 1.16964e-16
C5686 core_mux_0_24 vss 1.41588e-16
C5687 core_mux_0_23 vss 1.41588e-16
C5688 core_mux_0_25 vss 1.2312e-17
C5689 core_mux_0_24 vss 1.2312e-17
C5690 core_mux_0_26 vss 9.234e-17
C5691 core_mux_0_25 vss 9.234e-17
C5692 core_mux_0_27 vss 9.234e-17
C5693 core_mux_0_26 vss 9.234e-17
C5694 core_mux_0_8 vss 1.22239e-16
C5695 core_mux_0_7 vss 1.22239e-16
C5696 core_mux_0_10 vss 6.156e-17
C5697 core_mux_0_9 vss 6.156e-17
C5698 core_mux_0_11 vss 1.2312e-17
C5699 core_mux_0_10 vss 1.2312e-17
C5700 core_mux_0_12 vss 1.47744e-16
C5701 core_mux_0_11 vss 1.47744e-16
C5702 core_mux_0_13 vss 1.10808e-16
C5703 core_mux_0_12 vss 1.10808e-16
C5704 core_mux_0_4 vss 4.38566e-17
C5705 core_mux_0_3 vss 4.38566e-17
C5706 core_mux_0_5 vss 5.84755e-17
C5707 core_mux_0_4 vss 5.84755e-17
C5708 core_mux_0_6 vss 4.38566e-17
C5709 core_mux_0_5 vss 4.38566e-17

R130_1 n3810_1 n3810_11 0.001
R130_2 n3810_7 n3810_5 0.001
R130_3 n3810_9 n3810_6 0.001
R130_4 n3810_4 n3810_2 72
R130_5 n3810 n3810_4 43.2
R130_6 n3810_5 n3810_4 7.2
R130_7 n3810_7 n3810_8 0.108
R130_8 n3810_9 n3810_8 0.756
R130_9 n3810_10 n3810_9 0.324
R130_10 n3810_11 n3810_10 0.648

C5710 n3810_4 vss 8.21582e-17
C5711 n3810_2 vss 8.21582e-17
C5712 n3810 vss 5.086e-17
C5713 n3810_4 vss 5.086e-17
C5714 n3810_5 vss 3.15414e-17
C5715 n3810_4 vss 3.15414e-17
C5716 n3810_7 vss 3.65472e-17
C5717 n3810_8 vss 3.65472e-17
C5718 n3810_9 vss 8.14925e-17
C5719 n3810_8 vss 8.14925e-17
C5720 n3810_10 vss 4.07462e-17
C5721 n3810_9 vss 4.07462e-17
C5722 n3810_11 vss 6.79104e-17
C5723 n3810_10 vss 6.79104e-17

R131_1 core_nsel_1 core_nsel_46 0.001
R131_2 core_nsel_45 core_nsel_20 0.001
R131_3 core_nsel_43 core_nsel_30 0.001
R131_4 core_nsel_44 core_nsel_41 0.001
R131_5 core_nsel_42 core_nsel_56 0.001
R131_6 core_nsel_7 core_nsel_3 0.001
R131_7 core_nsel_17 core_nsel_12 0.001
R131_8 core_nsel_27 core_nsel_22 0.001
R131_9 core_nsel_36 core_nsel_31 0.001
R131_10 core_nsel_53 core_nsel_48 0.001
R131_11 core_nsel_9 core_nsel_6 0.001
R131_12 core_nsel_11 core_nsel_14 0.001
R131_13 core_nsel_38 core_nsel_35 0.001
R131_14 core_nsel_21 core_nsel_24 0.001
R131_15 core_nsel_47 core_nsel_50 0.001
R131_16 core_nsel_34 core_nsel_32 0.001
R131_17 core_nsel_33 core_nsel_32 0.001
R131_18 core_nsel_14 core_nsel_13 72
R131_19 core_nsel_15 core_nsel_14 43.2
R131_20 core_nsel_24 core_nsel_23 72
R131_21 core_nsel_25 core_nsel_24 43.2
R131_22 core_nsel_50 core_nsel_49 72
R131_23 core_nsel_51 core_nsel_50 43.2
R131_24 core_nsel_12 core_nsel_11 0.108
R131_25 core_nsel_34 core_nsel_33 0.216
R131_26 core_nsel_35 core_nsel_34 0.216
R131_27 core_nsel_36 core_nsel_35 0.108
R131_28 core_nsel_22 core_nsel_21 0.108
R131_29 core_nsel_48 core_nsel_47 0.108
R131_30 core_nsel_17 core_nsel_16 0.756
R131_31 core_nsel_18 core_nsel_17 0.324
R131_32 core_nsel_38 core_nsel_37 0.648
R131_33 core_nsel_39 core_nsel_38 0.432
R131_34 core_nsel_27 core_nsel_26 0.756
R131_35 core_nsel_28 core_nsel_27 0.324
R131_36 core_nsel_53 core_nsel_52 0.756
R131_37 core_nsel_54 core_nsel_53 0.324
R131_38 core_nsel_19 core_nsel_18 0.054
R131_39 core_nsel_20 core_nsel_19 0.108
R131_40 core_nsel_40 core_nsel_39 0.054
R131_41 core_nsel_41 core_nsel_40 0.108
R131_42 core_nsel_29 core_nsel_28 0.054
R131_43 core_nsel_30 core_nsel_29 0.108
R131_44 core_nsel_55 core_nsel_54 0.054
R131_45 core_nsel_56 core_nsel_55 0.108
R131_46 core_nsel_43 core_nsel_42 12.528
R131_47 core_nsel_44 core_nsel_43 1.188
R131_48 core_nsel_45 core_nsel_44 9.72
R131_49 core_nsel_46 core_nsel_45 2.808
R131_50 core_nsel_1 core_nsel_5 0.108
R131_51 core_nsel_3 core_nsel_2 0.756
R131_52 core_nsel_4 core_nsel_3 0.324
R131_53 core_nsel_5 core_nsel_4 0.054
R131_54 core_nsel_7 core_nsel_6 0.108
R131_55 core_nsel_9 core_nsel_8 72
R131_56 core_nsel core_nsel_9 43.2

C5724 core_nsel_14 vss 8.21582e-17
C5725 core_nsel_13 vss 8.21582e-17
C5726 core_nsel_15 vss 5.086e-17
C5727 core_nsel_14 vss 5.086e-17
C5728 core_nsel_24 vss 8.21582e-17
C5729 core_nsel_23 vss 8.21582e-17
C5730 core_nsel_25 vss 5.086e-17
C5731 core_nsel_24 vss 5.086e-17
C5732 core_nsel_50 vss 8.21582e-17
C5733 core_nsel_49 vss 8.21582e-17
C5734 core_nsel_51 vss 5.086e-17
C5735 core_nsel_50 vss 5.086e-17
C5736 core_nsel_12 vss 3.65472e-17
C5737 core_nsel_11 vss 3.65472e-17
C5738 core_nsel_34 vss 4.38566e-17
C5739 core_nsel_33 vss 4.38566e-17
C5740 core_nsel_35 vss 5.11661e-17
C5741 core_nsel_34 vss 5.11661e-17
C5742 core_nsel_36 vss 3.65472e-17
C5743 core_nsel_35 vss 3.65472e-17
C5744 core_nsel_22 vss 3.65472e-17
C5745 core_nsel_21 vss 3.65472e-17
C5746 core_nsel_48 vss 3.65472e-17
C5747 core_nsel_47 vss 3.65472e-17
C5748 core_nsel_17 vss 1.78524e-16
C5749 core_nsel_16 vss 1.78524e-16
C5750 core_nsel_18 vss 8.0028e-17
C5751 core_nsel_17 vss 8.0028e-17
C5752 core_nsel_38 vss 1.539e-16
C5753 core_nsel_37 vss 1.539e-16
C5754 core_nsel_39 vss 1.04652e-16
C5755 core_nsel_38 vss 1.04652e-16
C5756 core_nsel_27 vss 1.78524e-16
C5757 core_nsel_26 vss 1.78524e-16
C5758 core_nsel_28 vss 8.0028e-17
C5759 core_nsel_27 vss 8.0028e-17
C5760 core_nsel_53 vss 1.78524e-16
C5761 core_nsel_52 vss 1.78524e-16
C5762 core_nsel_54 vss 8.0028e-17
C5763 core_nsel_53 vss 8.0028e-17
C5764 core_nsel_19 vss 1.2312e-17
C5765 core_nsel_18 vss 1.2312e-17
C5766 core_nsel_20 vss 3.078e-17
C5767 core_nsel_19 vss 3.078e-17
C5768 core_nsel_40 vss 1.2312e-17
C5769 core_nsel_39 vss 1.2312e-17
C5770 core_nsel_41 vss 3.078e-17
C5771 core_nsel_40 vss 3.078e-17
C5772 core_nsel_29 vss 1.2312e-17
C5773 core_nsel_28 vss 1.2312e-17
C5774 core_nsel_30 vss 3.078e-17
C5775 core_nsel_29 vss 3.078e-17
C5776 core_nsel_55 vss 1.2312e-17
C5777 core_nsel_54 vss 1.2312e-17
C5778 core_nsel_56 vss 3.078e-17
C5779 core_nsel_55 vss 3.078e-17
C5780 core_nsel_43 vss 1.26313e-15
C5781 core_nsel_42 vss 1.26313e-15
C5782 core_nsel_44 vss 1.22239e-16
C5783 core_nsel_43 vss 1.22239e-16
C5784 core_nsel_45 vss 9.7791e-16
C5785 core_nsel_44 vss 9.7791e-16
C5786 core_nsel_46 vss 2.85224e-16
C5787 core_nsel_45 vss 2.85224e-16
C5788 core_nsel_1 vss 3.078e-17
C5789 core_nsel_5 vss 3.078e-17
C5790 core_nsel_3 vss 1.78524e-16
C5791 core_nsel_2 vss 1.78524e-16
C5792 core_nsel_4 vss 8.0028e-17
C5793 core_nsel_3 vss 8.0028e-17
C5794 core_nsel_5 vss 1.2312e-17
C5795 core_nsel_4 vss 1.2312e-17
C5796 core_nsel_7 vss 3.65472e-17
C5797 core_nsel_6 vss 3.65472e-17
C5798 core_nsel_9 vss 8.21582e-17
C5799 core_nsel_8 vss 8.21582e-17
C5800 core_nsel vss 5.086e-17
C5801 core_nsel_9 vss 5.086e-17

R132_1 core_regout_0_2 core_regout_0_4 0.001
R132_2 core_regout_0_5 core_regout_0_11 0.001
R132_3 core_regout_0_7 core_regout_0_17 0.001
R132_4 core_regout_0_8 core_regout_0_6 0.001
R132_5 core_regout_0_20 core_regout_0_19 0.001
R132_6 core_regout_0_14 core_regout_0_24 0.001
R132_7 core_regout_0_23 core_regout_0_18 0.001
R132_8 core_regout_0_25 core_regout_0_18 0.001
R132_9 core_regout_0_21 core_regout_0_19 0.001
R132_10 core_regout_0_20 core_regout_0_22 0.001
R132_11 core_regout_0_21 core_regout_0_25 0.648
R132_12 core_regout_0_22 core_regout_0_21 0.001
R132_13 core_regout_0_24 core_regout_0_23 0.108
R132_14 core_regout_0_25 core_regout_0_24 0.108
R132_15 core_regout_0_14 core_regout_0_13 0.378
R132_16 core_regout_0_15 core_regout_0_14 0.702
R132_17 core_regout_0_16 core_regout_0_15 0.054
R132_18 core_regout_0_17 core_regout_0_16 0.918
R132_19 core_regout_0_7 core_regout_0_6 5.184
R132_20 core_regout_0_9 core_regout_0_8 0.108
R132_21 core_regout_0_10 core_regout_0_9 0.054
R132_22 core_regout_0_11 core_regout_0_10 0.702
R132_23 core_regout_0_12 core_regout_0_11 0.378
R132_24 core_regout_0_5 core_regout_0_4 0.108
R132_25 core_regout_0_2 core_regout_0_1 72
R132_26 core_regout_0 core_regout_0_2 43.2

C5802 core_regout_0_20 vss 1.60808e-17
C5803 core_regout_0_22 vss 1.60808e-17
C5804 core_regout_0_21 vss 7.47014e-17
C5805 core_regout_0_25 vss 7.47014e-17
C5806 core_regout_0_22 vss 1.3157e-17
C5807 core_regout_0_21 vss 1.3157e-17
C5808 core_regout_0_24 vss 2.19283e-17
C5809 core_regout_0_23 vss 2.19283e-17
C5810 core_regout_0_25 vss 2.19283e-17
C5811 core_regout_0_24 vss 2.19283e-17
C5812 core_regout_0_14 vss 9.234e-17
C5813 core_regout_0_13 vss 9.234e-17
C5814 core_regout_0_15 vss 1.66212e-16
C5815 core_regout_0_14 vss 1.66212e-16
C5816 core_regout_0_16 vss 1.2312e-17
C5817 core_regout_0_15 vss 1.2312e-17
C5818 core_regout_0_17 vss 2.1546e-16
C5819 core_regout_0_16 vss 2.1546e-16
C5820 core_regout_0_7 vss 5.29701e-16
C5821 core_regout_0_6 vss 5.29701e-16
C5822 core_regout_0_9 vss 3.078e-17
C5823 core_regout_0_8 vss 3.078e-17
C5824 core_regout_0_10 vss 1.2312e-17
C5825 core_regout_0_9 vss 1.2312e-17
C5826 core_regout_0_11 vss 1.66212e-16
C5827 core_regout_0_10 vss 1.66212e-16
C5828 core_regout_0_12 vss 9.234e-17
C5829 core_regout_0_11 vss 9.234e-17
C5830 core_regout_0_5 vss 3.65472e-17
C5831 core_regout_0_4 vss 3.65472e-17
C5832 core_regout_0_2 vss 8.21582e-17
C5833 core_regout_0_1 vss 8.21582e-17
C5834 core_regout_0 vss 5.086e-17
C5835 core_regout_0_2 vss 5.086e-17

R133_1 n3914_1 n3914_11 0.001
R133_2 n3914_7 n3914_5 0.001
R133_3 n3914_9 n3914_6 0.001
R133_4 n3914_4 n3914_2 72
R133_5 n3914 n3914_4 43.2
R133_6 n3914_5 n3914_4 7.2
R133_7 n3914_7 n3914_8 0.108
R133_8 n3914_9 n3914_8 0.756
R133_9 n3914_10 n3914_9 0.324
R133_10 n3914_11 n3914_10 0.648

C5836 n3914_4 vss 8.21582e-17
C5837 n3914_2 vss 8.21582e-17
C5838 n3914 vss 5.086e-17
C5839 n3914_4 vss 5.086e-17
C5840 n3914_5 vss 3.15414e-17
C5841 n3914_4 vss 3.15414e-17
C5842 n3914_7 vss 3.65472e-17
C5843 n3914_8 vss 3.65472e-17
C5844 n3914_9 vss 8.14925e-17
C5845 n3914_8 vss 8.14925e-17
C5846 n3914_10 vss 4.07462e-17
C5847 n3914_9 vss 4.07462e-17
C5848 n3914_11 vss 6.79104e-17
C5849 n3914_10 vss 6.79104e-17

R134_1 core_int_1_7 core_int_1_18 0.001
R134_2 core_int_1_17 core_int_1_20 0.001
R134_3 core_int_1_19 core_int_1_22 0.001
R134_4 core_int_1_21 core_int_1_28 0.001
R134_5 core_int_1_30 core_int_1_23 0.001
R134_6 core_int_1_2 core_int_1_16 0.001
R134_7 core_int_1_13 core_int_1_5 0.001
R134_8 core_int_1_12 core_int_1_9 0.001
R134_9 core_int_1_25 core_int_1_33 0.001
R134_10 core_int_1_31 core_int_1_29 0.001
R134_11 core_int_1_32 core_int_1_29 0.001
R134_12 core_int_1_30 core_int_1_34 0.324
R134_13 core_int_1_32 core_int_1_31 0.216
R134_14 core_int_1_33 core_int_1_32 0.216
R134_15 core_int_1_34 core_int_1_33 0.108
R134_16 core_int_1_25 core_int_1_24 0.648
R134_17 core_int_1_26 core_int_1_25 0.486
R134_18 core_int_1_27 core_int_1_26 0.054
R134_19 core_int_1_28 core_int_1_27 0.27
R134_20 core_int_1_22 core_int_1_21 3.564
R134_21 core_int_1_20 core_int_1_19 0.108
R134_22 core_int_1_18 core_int_1_17 6.048
R134_23 core_int_1_7 core_int_1_11 0.378
R134_24 core_int_1_9 core_int_1_8 0.81
R134_25 core_int_1_10 core_int_1_9 0.324
R134_26 core_int_1_11 core_int_1_10 0.054
R134_27 core_int_1_5 core_int_1_4 115.2
R134_28 core_int_1 core_int_1_5 64.8
R134_29 core_int_1_12 core_int_1_13 0.216
R134_30 core_int_1_13 core_int_1_14 0.216
R134_31 core_int_1_15 core_int_1_14 1.62
R134_32 core_int_1_16 core_int_1_15 0.108
R134_33 core_int_1_2 core_int_1_1 115.2
R134_34 core_int_1_3 core_int_1_2 43.2

C5850 core_int_1_30 vss 4.07462e-17
C5851 core_int_1_34 vss 4.07462e-17
C5852 core_int_1_32 vss 4.38566e-17
C5853 core_int_1_31 vss 4.38566e-17
C5854 core_int_1_33 vss 4.38566e-17
C5855 core_int_1_32 vss 4.38566e-17
C5856 core_int_1_34 vss 3.65472e-17
C5857 core_int_1_33 vss 3.65472e-17
C5858 core_int_1_25 vss 1.47744e-16
C5859 core_int_1_24 vss 1.47744e-16
C5860 core_int_1_26 vss 1.10808e-16
C5861 core_int_1_25 vss 1.10808e-16
C5862 core_int_1_27 vss 1.2312e-17
C5863 core_int_1_26 vss 1.2312e-17
C5864 core_int_1_28 vss 6.156e-17
C5865 core_int_1_27 vss 6.156e-17
C5866 core_int_1_22 vss 3.66716e-16
C5867 core_int_1_21 vss 3.66716e-16
C5868 core_int_1_20 vss 3.078e-17
C5869 core_int_1_19 vss 3.078e-17
C5870 core_int_1_18 vss 6.11194e-16
C5871 core_int_1_17 vss 6.11194e-16
C5872 core_int_1_7 vss 9.234e-17
C5873 core_int_1_11 vss 9.234e-17
C5874 core_int_1_9 vss 1.8468e-16
C5875 core_int_1_8 vss 1.8468e-16
C5876 core_int_1_10 vss 7.3872e-17
C5877 core_int_1_9 vss 7.3872e-17
C5878 core_int_1_11 vss 1.2312e-17
C5879 core_int_1_10 vss 1.2312e-17
C5880 core_int_1_5 vss 1.25194e-16
C5881 core_int_1_4 vss 1.25194e-16
C5882 core_int_1 vss 7.43336e-17
C5883 core_int_1_5 vss 7.43336e-17
C5884 core_int_1_12 vss 4.38566e-17
C5885 core_int_1_13 vss 4.38566e-17
C5886 core_int_1_13 vss 2.71642e-17
C5887 core_int_1_14 vss 2.71642e-17
C5888 core_int_1_15 vss 1.69776e-16
C5889 core_int_1_14 vss 1.69776e-16
C5890 core_int_1_16 vss 2.92378e-17
C5891 core_int_1_15 vss 2.92378e-17
C5892 core_int_1_2 vss 1.25194e-16
C5893 core_int_1_1 vss 1.25194e-16
C5894 core_int_1_3 vss 5.086e-17
C5895 core_int_1_2 vss 5.086e-17

R135_1 core_carry_0_1 core_carry_0_6 0.001
R135_2 core_carry_0_7 core_carry_0_15 0.001
R135_3 core_carry_0_5 core_carry_0_11 0.001
R135_4 core_carry_0_12 core_carry_0_42 0.001
R135_5 core_carry_0_41 core_carry_0_27 0.001
R135_6 core_carry_0_40 core_carry_0_32 0.001
R135_7 core_carry_0_39 core_carry_0_47 0.001
R135_8 core_carry_0_22 core_carry_0_17 0.001
R135_9 core_carry_0_24 core_carry_0_21 0.001
R135_10 core_carry_0_19 core_carry_0_18 0.001
R135_11 core_carry_0_20 core_carry_0_18 0.001
R135_12 core_carry_0_29 core_carry_0_38 0.001
R135_13 core_carry_0_44 core_carry_0_53 0.001
R135_14 core_carry_0_51 core_carry_0_49 0.001
R135_15 core_carry_0_36 core_carry_0_34 0.001
R135_16 core_carry_0_34 core_carry_0_33 72
R135_17 core_carry_0_35 core_carry_0_34 50.4
R135_18 core_carry_0_49 core_carry_0_48 72
R135_19 core_carry_0_50 core_carry_0_49 50.4
R135_20 core_carry_0_36 core_carry_0_37 0.216
R135_21 core_carry_0_51 core_carry_0_52 0.216
R135_22 core_carry_0_38 core_carry_0_37 0.216
R135_23 core_carry_0_53 core_carry_0_52 0.216
R135_24 core_carry_0_20 core_carry_0_19 0.216
R135_25 core_carry_0_21 core_carry_0_20 0.216
R135_26 core_carry_0_22 core_carry_0_21 0.216
R135_27 core_carry_0_24 core_carry_0_23 0.648
R135_28 core_carry_0_25 core_carry_0_24 0.432
R135_29 core_carry_0_29 core_carry_0_28 0.486
R135_30 core_carry_0_30 core_carry_0_29 0.648
R135_31 core_carry_0_44 core_carry_0_43 0.486
R135_32 core_carry_0_45 core_carry_0_44 0.648
R135_33 core_carry_0_26 core_carry_0_25 0.054
R135_34 core_carry_0_27 core_carry_0_26 0.27
R135_35 core_carry_0_31 core_carry_0_30 0.054
R135_36 core_carry_0_32 core_carry_0_31 0.27
R135_37 core_carry_0_46 core_carry_0_45 0.054
R135_38 core_carry_0_47 core_carry_0_46 0.27
R135_39 core_carry_0_40 core_carry_0_39 1.62
R135_40 core_carry_0_41 core_carry_0_40 6.804
R135_41 core_carry_0_42 core_carry_0_41 2.376
R135_42 core_carry_0_10 core_carry_0_8 115.2
R135_43 core_carry_0 core_carry_0_10 64.8
R135_44 core_carry_0_13 core_carry_0_12 0.81
R135_45 core_carry_0_11 core_carry_0_10 7.2
R135_46 core_carry_0_14 core_carry_0_13 0.054
R135_47 core_carry_0_15 core_carry_0_14 0.702
R135_48 core_carry_0_16 core_carry_0_15 0.378
R135_49 core_carry_0_6 core_carry_0_5 0.756
R135_50 core_carry_0_7 core_carry_0_6 0.108
R135_51 core_carry_0_3 core_carry_0_1 7.2
R135_52 core_carry_0_3 core_carry_0_2 115.2
R135_53 core_carry_0_4 core_carry_0_3 43.2

C5896 core_carry_0_34 vss 8.21582e-17
C5897 core_carry_0_33 vss 8.21582e-17
C5898 core_carry_0_35 vss 5.86844e-17
C5899 core_carry_0_34 vss 5.86844e-17
C5900 core_carry_0_49 vss 8.21582e-17
C5901 core_carry_0_48 vss 8.21582e-17
C5902 core_carry_0_50 vss 5.86844e-17
C5903 core_carry_0_49 vss 5.86844e-17
C5904 core_carry_0_36 vss 2.71642e-17
C5905 core_carry_0_37 vss 2.71642e-17
C5906 core_carry_0_51 vss 2.71642e-17
C5907 core_carry_0_52 vss 2.71642e-17
C5908 core_carry_0_38 vss 2.54664e-17
C5909 core_carry_0_37 vss 2.54664e-17
C5910 core_carry_0_53 vss 2.54664e-17
C5911 core_carry_0_52 vss 2.54664e-17
C5912 core_carry_0_20 vss 4.38566e-17
C5913 core_carry_0_19 vss 4.38566e-17
C5914 core_carry_0_21 vss 5.11661e-17
C5915 core_carry_0_20 vss 5.11661e-17
C5916 core_carry_0_22 vss 5.11661e-17
C5917 core_carry_0_21 vss 5.11661e-17
C5918 core_carry_0_24 vss 1.539e-16
C5919 core_carry_0_23 vss 1.539e-16
C5920 core_carry_0_25 vss 1.04652e-16
C5921 core_carry_0_24 vss 1.04652e-16
C5922 core_carry_0_29 vss 1.10808e-16
C5923 core_carry_0_28 vss 1.10808e-16
C5924 core_carry_0_30 vss 1.47744e-16
C5925 core_carry_0_29 vss 1.47744e-16
C5926 core_carry_0_44 vss 1.10808e-16
C5927 core_carry_0_43 vss 1.10808e-16
C5928 core_carry_0_45 vss 1.47744e-16
C5929 core_carry_0_44 vss 1.47744e-16
C5930 core_carry_0_26 vss 1.2312e-17
C5931 core_carry_0_25 vss 1.2312e-17
C5932 core_carry_0_27 vss 6.156e-17
C5933 core_carry_0_26 vss 6.156e-17
C5934 core_carry_0_31 vss 1.2312e-17
C5935 core_carry_0_30 vss 1.2312e-17
C5936 core_carry_0_32 vss 6.156e-17
C5937 core_carry_0_31 vss 6.156e-17
C5938 core_carry_0_46 vss 1.2312e-17
C5939 core_carry_0_45 vss 1.2312e-17
C5940 core_carry_0_47 vss 6.156e-17
C5941 core_carry_0_46 vss 6.156e-17
C5942 core_carry_0_40 vss 1.62985e-16
C5943 core_carry_0_39 vss 1.62985e-16
C5944 core_carry_0_41 vss 6.92686e-16
C5945 core_carry_0_40 vss 6.92686e-16
C5946 core_carry_0_42 vss 2.44477e-16
C5947 core_carry_0_41 vss 2.44477e-16
C5948 core_carry_0_10 vss 1.25194e-16
C5949 core_carry_0_8 vss 1.25194e-16
C5950 core_carry_0 vss 7.43336e-17
C5951 core_carry_0_10 vss 7.43336e-17
C5952 core_carry_0_13 vss 1.8468e-16
C5953 core_carry_0_12 vss 1.8468e-16
C5954 core_carry_0_11 vss 3.15414e-17
C5955 core_carry_0_10 vss 3.15414e-17
C5956 core_carry_0_14 vss 1.2312e-17
C5957 core_carry_0_13 vss 1.2312e-17
C5958 core_carry_0_15 vss 1.66212e-16
C5959 core_carry_0_14 vss 1.66212e-16
C5960 core_carry_0_16 vss 9.234e-17
C5961 core_carry_0_15 vss 9.234e-17
C5962 core_carry_0_6 vss 8.14925e-17
C5963 core_carry_0_5 vss 8.14925e-17
C5964 core_carry_0_7 vss 3.65472e-17
C5965 core_carry_0_6 vss 3.65472e-17
C5966 core_carry_0_3 vss 3.15414e-17
C5967 core_carry_0_1 vss 3.15414e-17
C5968 core_carry_0_3 vss 1.25194e-16
C5969 core_carry_0_2 vss 1.25194e-16
C5970 core_carry_0_4 vss 5.086e-17
C5971 core_carry_0_3 vss 5.086e-17

R136_1 core_regout_1_15 core_regout_1_2 0.001
R136_2 core_regout_1_1 core_regout_1_12 0.001
R136_3 core_regout_1 core_regout_1_23 0.001
R136_4 core_regout_1 core_regout_1_25 0.001
R136_5 core_regout_1_9 core_regout_1_4 0.001
R136_6 core_regout_1_3 core_regout_1_6 0.001
R136_7 core_regout_1_22 core_regout_1_14 0.001
R136_8 core_regout_1_20 core_regout_1_14 0.001
R136_9 core_regout_1_21 core_regout_1_17 0.001
R136_10 core_regout_1_6 core_regout_1_5 72
R136_11 core_regout_1_7 core_regout_1_6 43.2
R136_12 core_regout_1_4 core_regout_1_3 0.108
R136_13 core_regout_1_9 core_regout_1_8 0.756
R136_14 core_regout_1_10 core_regout_1_9 0.324
R136_15 core_regout_1_11 core_regout_1_10 0.054
R136_16 core_regout_1_12 core_regout_1_11 0.27
R136_17 core_regout_1_2 core_regout_1_1 8.1
R136_18 core_regout_1_15 core_regout_1_19 0.27
R136_19 core_regout_1_17 core_regout_1_16 0.378
R136_20 core_regout_1_18 core_regout_1_17 0.702
R136_21 core_regout_1_19 core_regout_1_18 0.054
R136_22 core_regout_1_21 core_regout_1_20 0.108
R136_23 core_regout_1_22 core_regout_1_21 0.108
R136_24 core_regout_1_23 core_regout_1_22 0.648
R136_25 core_regout_1_24 core_regout_1_23 0.001
R136_26 core_regout_1_25 core_regout_1_24 0.001

C5972 core_regout_1_6 vss 8.21582e-17
C5973 core_regout_1_5 vss 8.21582e-17
C5974 core_regout_1_7 vss 5.086e-17
C5975 core_regout_1_6 vss 5.086e-17
C5976 core_regout_1_4 vss 3.65472e-17
C5977 core_regout_1_3 vss 3.65472e-17
C5978 core_regout_1_9 vss 1.78524e-16
C5979 core_regout_1_8 vss 1.78524e-16
C5980 core_regout_1_10 vss 8.0028e-17
C5981 core_regout_1_9 vss 8.0028e-17
C5982 core_regout_1_11 vss 1.2312e-17
C5983 core_regout_1_10 vss 1.2312e-17
C5984 core_regout_1_12 vss 6.156e-17
C5985 core_regout_1_11 vss 6.156e-17
C5986 core_regout_1_2 vss 8.14925e-16
C5987 core_regout_1_1 vss 8.14925e-16
C5988 core_regout_1_15 vss 6.156e-17
C5989 core_regout_1_19 vss 6.156e-17
C5990 core_regout_1_17 vss 9.234e-17
C5991 core_regout_1_16 vss 9.234e-17
C5992 core_regout_1_18 vss 1.66212e-16
C5993 core_regout_1_17 vss 1.66212e-16
C5994 core_regout_1_19 vss 1.2312e-17
C5995 core_regout_1_18 vss 1.2312e-17
C5996 core_regout_1_21 vss 2.19283e-17
C5997 core_regout_1_20 vss 2.19283e-17
C5998 core_regout_1_22 vss 2.19283e-17
C5999 core_regout_1_21 vss 2.19283e-17
C6000 core_regout_1_23 vss 7.47014e-17
C6001 core_regout_1_22 vss 7.47014e-17
C6002 core_regout_1_24 vss 1.3157e-17
C6003 core_regout_1_23 vss 1.3157e-17
C6004 core_regout_1_25 vss 1.60808e-17
C6005 core_regout_1_24 vss 1.60808e-17

R137_1 n4048_1 n4048_10 0.001
R137_2 n4048_9 n4048_5 0.001
R137_3 n4048_6 n4048_3 0.001
R137_4 n4048_8 n4048_5 0.001
R137_5 n4048_3 n4048_2 115.2
R137_6 n4048 n4048_3 43.2
R137_7 n4048_6 n4048_7 0.54
R137_8 n4048_9 n4048_7 2.376
R137_9 n4048_9 n4048_8 0.216
R137_10 n4048_11 n4048_9 0.756
R137_11 n4048_11 n4048_10 0.324

C6006 n4048_3 vss 1.25194e-16
C6007 n4048_2 vss 1.25194e-16
C6008 n4048 vss 5.086e-17
C6009 n4048_3 vss 5.086e-17
C6010 n4048_6 vss 5.43283e-17
C6011 n4048_7 vss 5.43283e-17
C6012 n4048_9 vss 2.44477e-16
C6013 n4048_7 vss 2.44477e-16
C6014 n4048_9 vss 3.83746e-17
C6015 n4048_8 vss 3.83746e-17
C6016 n4048_11 vss 8.65858e-17
C6017 n4048_9 vss 8.65858e-17
C6018 n4048_11 vss 4.07462e-17
C6019 n4048_10 vss 4.07462e-17

R138_1 n4065 n4065_12 0.001
R138_2 n4065_10 n4065_5 0.001
R138_3 n4065_8 n4065_6 0.001
R138_4 n4065_7 n4065_6 0.001
R138_5 n4065_2 n4065_3 72
R138_6 n4065_8 n4065_7 0.108
R138_7 n4065_4 n4065_3 64.8
R138_8 n4065_8 n4065_9 0.324
R138_9 n4065_5 n4065_4 21.6
R138_10 n4065_10 n4065_9 0.648
R138_11 n4065_11 n4065_10 0.324
R138_12 n4065_12 n4065_11 0.324

C6020 n4065_2 vss 8.21582e-17
C6021 n4065_3 vss 8.21582e-17
C6022 n4065_8 vss 3.10651e-17
C6023 n4065_7 vss 3.10651e-17
C6024 n4065_4 vss 7.04214e-17
C6025 n4065_3 vss 7.04214e-17
C6026 n4065_8 vss 4.07462e-17
C6027 n4065_9 vss 4.07462e-17
C6028 n4065_5 vss 2.34738e-17
C6029 n4065_4 vss 2.34738e-17
C6030 n4065_10 vss 7.47014e-17
C6031 n4065_9 vss 7.47014e-17
C6032 n4065_11 vss 3.39552e-17
C6033 n4065_10 vss 3.39552e-17
C6034 n4065_12 vss 4.07462e-17
C6035 n4065_11 vss 4.07462e-17

R139_1 n4080 n4080_10 0.001
R139_2 n4080_7 n4080_3 0.001
R139_3 n4080_6 n4080_5 0.001
R139_4 n4080_3 n4080_2 72
R139_5 n4080_4 n4080_3 144
R139_6 n4080_7 n4080_6 0.216
R139_7 n4080_7 n4080_8 0.54
R139_8 n4080_9 n4080_8 0.648
R139_9 n4080_10 n4080_9 0.432

C6036 n4080_3 vss 7.8246e-17
C6037 n4080_2 vss 7.8246e-17
C6038 n4080_4 vss 1.6236e-16
C6039 n4080_3 vss 1.6236e-16
C6040 n4080_7 vss 3.22574e-17
C6041 n4080_6 vss 3.22574e-17
C6042 n4080_7 vss 5.60261e-17
C6043 n4080_8 vss 5.60261e-17
C6044 n4080_9 vss 7.47014e-17
C6045 n4080_8 vss 7.47014e-17
C6046 n4080_10 vss 4.75373e-17
C6047 n4080_9 vss 4.75373e-17

R140_1 n4085 n4085_5 0.001
R140_2 n4085_3 n4085_2 0.001
R140_3 n4085_4 n4085_2 0.001
R140_4 n4085_4 n4085_3 0.108
R140_5 n4085_5 n4085_4 1.08

C6048 n4085_4 vss 3.10651e-17
C6049 n4085_3 vss 3.10651e-17
C6050 n4085_5 vss 1.18843e-16
C6051 n4085_4 vss 1.18843e-16

R141_1 core_l1_dff_s_1 core_l1_dff_s_6 0.001
R141_2 core_l1_dff_s_3 core_l1_dff_s_12 0.001
R141_3 core_l1_dff_s_4 core_l1_dff_s_2 0.001
R141_4 core_l1_dff_s core_l1_dff_s_9 180
R141_5 core_l1_dff_s_11 core_l1_dff_s_8 50.4
R141_6 core_l1_dff_s_11 core_l1_dff_s_9 43.2
R141_7 core_l1_dff_s_10 core_l1_dff_s_12 43.2
R141_8 core_l1_dff_s_12 core_l1_dff_s_11 28.8
R141_9 core_l1_dff_s_5 core_l1_dff_s_3 0.54
R141_10 core_l1_dff_s_5 core_l1_dff_s_4 0.648
R141_11 core_l1_dff_s_6 core_l1_dff_s_5 0.54

C6052 core_l1_dff_s vss 1.97571e-16
C6053 core_l1_dff_s_9 vss 1.97571e-16
C6054 core_l1_dff_s_11 vss 5.47722e-17
C6055 core_l1_dff_s_8 vss 5.47722e-17
C6056 core_l1_dff_s_11 vss 4.69476e-17
C6057 core_l1_dff_s_9 vss 4.69476e-17
C6058 core_l1_dff_s_10 vss 4.69476e-17
C6059 core_l1_dff_s_12 vss 4.69476e-17
C6060 core_l1_dff_s_12 vss 3.12984e-17
C6061 core_l1_dff_s_11 vss 3.12984e-17
C6062 core_l1_dff_s_5 vss 5.43283e-17
C6063 core_l1_dff_s_3 vss 5.43283e-17
C6064 core_l1_dff_s_5 vss 7.47014e-17
C6065 core_l1_dff_s_4 vss 7.47014e-17
C6066 core_l1_dff_s_6 vss 5.43283e-17
C6067 core_l1_dff_s_5 vss 5.43283e-17

R142_1 n4115 n4115_18 0.001
R142_2 n4115_17 n4115_7 0.001
R142_3 n4115_12 n4115_9 0.001
R142_4 n4115_15 n4115_14 0.001
R142_5 n4115_13 n4115_11 0.001
R142_6 n4115_6 n4115_4 0.001
R142_7 n4115_3 n4115_2 0.001
R142_8 n4115_10 n4115_9 43.2
R142_9 n4115_12 n4115_11 0.54
R142_10 n4115_6 n4115_5 36
R142_11 n4115_4 n4115_3 0.108
R142_12 n4115_14 n4115_13 57.6
R142_13 n4115_7 n4115_6 93.6
R142_14 n4115_16 n4115_15 0.54
R142_15 n4115_8 n4115_7 86.4
R142_16 n4115_17 n4115_16 0.972
R142_17 n4115_18 n4115_17 0.216

C6068 n4115_10 vss 5.086e-17
C6069 n4115_9 vss 5.086e-17
C6070 n4115_12 vss 5.43283e-17
C6071 n4115_11 vss 5.43283e-17
C6072 n4115_6 vss 3.9123e-17
C6073 n4115_5 vss 3.9123e-17
C6074 n4115_4 vss 2.92378e-17
C6075 n4115_3 vss 2.92378e-17
C6076 n4115_14 vss 6.25968e-17
C6077 n4115_13 vss 6.25968e-17
C6078 n4115_7 vss 1.0172e-16
C6079 n4115_6 vss 1.0172e-16
C6080 n4115_16 vss 5.43283e-17
C6081 n4115_15 vss 5.43283e-17
C6082 n4115_8 vss 9.97636e-17
C6083 n4115_7 vss 9.97636e-17
C6084 n4115_17 vss 1.00168e-16
C6085 n4115_16 vss 1.00168e-16
C6086 n4115_18 vss 2.71642e-17
C6087 n4115_17 vss 2.71642e-17

R143_1 n4126 n4126_5 0.001
R143_2 n4126_4 n4126_2 0.001
R143_3 n4126_3 n4126_2 0.001
R143_4 n4126_4 n4126_3 0.108
R143_5 n4126_5 n4126_4 1.188

C6088 n4126_4 vss 2.92378e-17
C6089 n4126_3 vss 2.92378e-17
C6090 n4126_5 vss 1.22239e-16
C6091 n4126_4 vss 1.22239e-16

R144_1 core_l1_dff_m core_l1_dff_m_12 0.001
R144_2 core_l1_dff_m_7 core_l1_dff_m_2 0.001
R144_3 core_l1_dff_m_6 core_l1_dff_m_4 0.001
R144_4 core_l1_dff_m_4 core_l1_dff_m_3 64.8
R144_5 core_l1_dff_m_5 core_l1_dff_m_4 93.6
R144_6 core_l1_dff_m_8 core_l1_dff_m_6 0.648
R144_7 core_l1_dff_m_8 core_l1_dff_m_7 0.216
R144_8 core_l1_dff_m_9 core_l1_dff_m_8 0.108
R144_9 core_l1_dff_m_10 core_l1_dff_m_9 0.648
R144_10 core_l1_dff_m_10 core_l1_dff_m_11 0.108
R144_11 core_l1_dff_m_12 core_l1_dff_m_11 0.216

C6092 core_l1_dff_m_4 vss 7.04214e-17
C6093 core_l1_dff_m_3 vss 7.04214e-17
C6094 core_l1_dff_m_5 vss 1.0172e-16
C6095 core_l1_dff_m_4 vss 1.0172e-16
C6096 core_l1_dff_m_8 vss 6.79104e-17
C6097 core_l1_dff_m_6 vss 6.79104e-17
C6098 core_l1_dff_m_8 vss 2.71642e-17
C6099 core_l1_dff_m_7 vss 2.71642e-17
C6100 core_l1_dff_m_9 vss 1.35821e-17
C6101 core_l1_dff_m_8 vss 1.35821e-17
C6102 core_l1_dff_m_10 vss 6.79104e-17
C6103 core_l1_dff_m_9 vss 6.79104e-17
C6104 core_l1_dff_m_10 vss 1.35821e-17
C6105 core_l1_dff_m_11 vss 1.35821e-17
C6106 core_l1_dff_m_12 vss 2.71642e-17
C6107 core_l1_dff_m_11 vss 2.71642e-17

R3_1 a_2_50 a_2_1 0.001
R3_2 a_2_48 a_2_1 0.001
R3_3 a_2_49 a_2_1 0.001
R3_4 a_2_47 a_2_1 0.001
R3_5 a_2_46 a_2_1 0.001
R3_6 a_2_45 a_2_1 0.001
R3_7 a_2_44 a_2_1 0.001
R3_8 a_2_43 a_2_1 0.001
R3_9 a_2_41 a_2_2 0.001
R3_10 a_2_42 a_2_2 0.001
R3_11 a_2_39 a_2_2 0.001
R3_12 a_2_40 a_2_2 0.001
R3_13 a_2_36 a_2_2 0.001
R3_14 a_2_37 a_2_2 0.001
R3_15 a_2_38 a_2_2 0.001
R3_16 a_2_35 a_2_2 0.001
R3_17 a_2_34 a_2_2 0.001
R3_18 a_2_33 a_2_2 0.001
R3_19 a_2_32 a_2_2 0.001
R3_20 a_2_30 a_2_2 0.001
R3_21 a_2_31 a_2_2 0.001
R3_22 a_2_28 a_2_2 0.001
R3_23 a_2_29 a_2_2 0.001
R3_24 a_2_27 a_2_2 0.001
R3_25 a_2_26 a_2_2 0.001
R3_26 a_2_24 a_2_2 0.001
R3_27 a_2_25 a_2_2 0.001
R3_28 a_2_23 a_2_2 0.001
R3_29 a_2_79 a_2_3 0.001
R3_30 a_2_77 a_2_3 0.001
R3_31 a_2_78 a_2_3 0.001
R3_32 a_2_76 a_2_3 0.001
R3_33 a_2_75 a_2_3 0.001
R3_34 a_2_73 a_2_3 0.001
R3_35 a_2_74 a_2_3 0.001
R3_36 a_2_72 a_2_3 0.001
R3_37 a_2_70 a_2_4 0.001
R3_38 a_2_71 a_2_4 0.001
R3_39 a_2_68 a_2_4 0.001
R3_40 a_2_69 a_2_4 0.001
R3_41 a_2_66 a_2_4 0.001
R3_42 a_2_65 a_2_4 0.001
R3_43 a_2_67 a_2_4 0.001
R3_44 a_2_63 a_2_4 0.001
R3_45 a_2_64 a_2_4 0.001
R3_46 a_2_62 a_2_4 0.001
R3_47 a_2_61 a_2_4 0.001
R3_48 a_2_59 a_2_4 0.001
R3_49 a_2_60 a_2_4 0.001
R3_50 a_2_58 a_2_4 0.001
R3_51 a_2_57 a_2_4 0.001
R3_52 a_2_55 a_2_4 0.001
R3_53 a_2_56 a_2_4 0.001
R3_54 a_2_54 a_2_4 0.001
R3_55 a_2_53 a_2_4 0.001
R3_56 a_2_52 a_2_4 0.001
R3_57 a_2_14 a_2_5 0.001
R3_58 a_2_13 a_2_8 0.001
R3_59 a_2 a_2_11 0.001
R3_60 a_2_6 a_2_5 21.6
R3_61 a_2_8 a_2_7 7.2
R3_62 a_2_9 a_2_8 7.2
R3_63 a_2_10 a_2_9 14.4
R3_64 a_2_13 a_2_12 0.001
R3_65 a_2_16 a_2_13 0.216
R3_66 a_2_14 a_2_16 0.216
R3_67 a_2_15 a_2_14 0.001
R3_68 a_2_16 a_2_17 0.324
R3_69 a_2_18 a_2_17 2.268
R3_70 a_2_19 a_2_18 1.08
R3_71 a_2_20 a_2_19 0.001
R3_72 a_2_21 a_2_20 0.001
R3_73 a_2_51 a_2_21 0.216
R3_74 a_2_23 a_2_22 0.001
R3_75 a_2_24 a_2_23 0.108
R3_76 a_2_25 a_2_24 0.108
R3_77 a_2_26 a_2_25 0.108
R3_78 a_2_27 a_2_26 0.108
R3_79 a_2_28 a_2_27 0.108
R3_80 a_2_29 a_2_28 0.108
R3_81 a_2_30 a_2_29 0.108
R3_82 a_2_31 a_2_30 0.108
R3_83 a_2_32 a_2_31 0.108
R3_84 a_2_33 a_2_32 0.108
R3_85 a_2_34 a_2_33 0.108
R3_86 a_2_35 a_2_34 0.108
R3_87 a_2_36 a_2_35 0.108
R3_88 a_2_37 a_2_36 0.108
R3_89 a_2_38 a_2_37 0.108
R3_90 a_2_39 a_2_38 0.108
R3_91 a_2_40 a_2_39 0.108
R3_92 a_2_41 a_2_40 0.108
R3_93 a_2_42 a_2_41 0.108
R3_94 a_2_43 a_2_42 0.864
R3_95 a_2_44 a_2_43 0.108
R3_96 a_2_45 a_2_44 0.108
R3_97 a_2_46 a_2_45 0.108
R3_98 a_2_47 a_2_46 0.108
R3_99 a_2_48 a_2_47 0.108
R3_100 a_2_49 a_2_48 0.108
R3_101 a_2_50 a_2_49 0.108
R3_102 a_2_81 a_2_50 0.54
R3_103 a_2_52 a_2_51 0.001
R3_104 a_2_53 a_2_52 0.108
R3_105 a_2_54 a_2_53 0.108
R3_106 a_2_55 a_2_54 0.108
R3_107 a_2_56 a_2_55 0.108
R3_108 a_2_57 a_2_56 0.108
R3_109 a_2_58 a_2_57 0.108
R3_110 a_2_59 a_2_58 0.108
R3_111 a_2_60 a_2_59 0.108
R3_112 a_2_61 a_2_60 0.108
R3_113 a_2_62 a_2_61 0.108
R3_114 a_2_63 a_2_62 0.108
R3_115 a_2_64 a_2_63 0.108
R3_116 a_2_65 a_2_64 0.108
R3_117 a_2_66 a_2_65 0.108
R3_118 a_2_67 a_2_66 0.108
R3_119 a_2_68 a_2_67 0.108
R3_120 a_2_69 a_2_68 0.108
R3_121 a_2_70 a_2_69 0.108
R3_122 a_2_71 a_2_70 0.108
R3_123 a_2_72 a_2_71 0.864
R3_124 a_2_73 a_2_72 0.108
R3_125 a_2_74 a_2_73 0.108
R3_126 a_2_75 a_2_74 0.108
R3_127 a_2_76 a_2_75 0.108
R3_128 a_2_77 a_2_76 0.108
R3_129 a_2_78 a_2_77 0.108
R3_130 a_2_79 a_2_78 0.108
R3_131 a_2_82 a_2_79 0.54
R3_132 a_2_82 a_2_80 0.001
R3_133 a_2_81 a_2_82 0.108
R3_134 a_2_83 a_2_82 0.54
R3_135 a_2_84 a_2_83 0.001
R3_136 a_2 a_2_84 0.001

C6108 a_2_6 vss 9.46242e-17
C6109 a_2_5 vss 9.46242e-17
C6110 a_2_8 vss 3.15414e-17
C6111 a_2_7 vss 3.15414e-17
C6112 a_2_9 vss 3.15414e-17
C6113 a_2_8 vss 3.15414e-17
C6114 a_2_10 vss 6.30828e-17
C6115 a_2_9 vss 6.30828e-17
C6116 a_2_13 vss 1.40901e-17
C6117 a_2_12 vss 1.40901e-17
C6118 a_2_16 vss 7.82784e-17
C6119 a_2_13 vss 7.82784e-17
C6120 a_2_14 vss 7.04506e-17
C6121 a_2_16 vss 7.04506e-17
C6122 a_2_15 vss 1.40901e-17
C6123 a_2_14 vss 1.40901e-17
C6124 a_2_16 vss 9.39341e-17
C6125 a_2_17 vss 9.39341e-17
C6126 a_2_18 vss 6.18399e-16
C6127 a_2_17 vss 6.18399e-16
C6128 a_2_19 vss 2.97458e-16
C6129 a_2_18 vss 2.97458e-16
C6130 a_2_20 vss 2.50491e-17
C6131 a_2_19 vss 2.50491e-17
C6132 a_2_21 vss 1.25245e-17
C6133 a_2_20 vss 1.25245e-17
C6134 a_2_51 vss 8.14095e-17
C6135 a_2_21 vss 8.14095e-17
C6136 a_2_23 vss 1.40901e-17
C6137 a_2_22 vss 1.40901e-17
C6138 a_2_24 vss 3.13114e-17
C6139 a_2_23 vss 3.13114e-17
C6140 a_2_25 vss 3.13114e-17
C6141 a_2_24 vss 3.13114e-17
C6142 a_2_26 vss 3.13114e-17
C6143 a_2_25 vss 3.13114e-17
C6144 a_2_27 vss 3.13114e-17
C6145 a_2_26 vss 3.13114e-17
C6146 a_2_28 vss 3.13114e-17
C6147 a_2_27 vss 3.13114e-17
C6148 a_2_29 vss 3.13114e-17
C6149 a_2_28 vss 3.13114e-17
C6150 a_2_30 vss 3.13114e-17
C6151 a_2_29 vss 3.13114e-17
C6152 a_2_31 vss 3.13114e-17
C6153 a_2_30 vss 3.13114e-17
C6154 a_2_32 vss 3.13114e-17
C6155 a_2_31 vss 3.13114e-17
C6156 a_2_33 vss 3.13114e-17
C6157 a_2_32 vss 3.13114e-17
C6158 a_2_34 vss 3.13114e-17
C6159 a_2_33 vss 3.13114e-17
C6160 a_2_35 vss 3.13114e-17
C6161 a_2_34 vss 3.13114e-17
C6162 a_2_36 vss 3.13114e-17
C6163 a_2_35 vss 3.13114e-17
C6164 a_2_37 vss 3.13114e-17
C6165 a_2_36 vss 3.13114e-17
C6166 a_2_38 vss 3.13114e-17
C6167 a_2_37 vss 3.13114e-17
C6168 a_2_39 vss 3.13114e-17
C6169 a_2_38 vss 3.13114e-17
C6170 a_2_40 vss 3.13114e-17
C6171 a_2_39 vss 3.13114e-17
C6172 a_2_41 vss 3.13114e-17
C6173 a_2_40 vss 3.13114e-17
C6174 a_2_42 vss 3.13114e-17
C6175 a_2_41 vss 3.13114e-17
C6176 a_2_43 vss 2.42663e-16
C6177 a_2_42 vss 2.42663e-16
C6178 a_2_44 vss 3.13114e-17
C6179 a_2_43 vss 3.13114e-17
C6180 a_2_45 vss 3.13114e-17
C6181 a_2_44 vss 3.13114e-17
C6182 a_2_46 vss 3.13114e-17
C6183 a_2_45 vss 3.13114e-17
C6184 a_2_47 vss 3.13114e-17
C6185 a_2_46 vss 3.13114e-17
C6186 a_2_48 vss 3.13114e-17
C6187 a_2_47 vss 3.13114e-17
C6188 a_2_49 vss 3.13114e-17
C6189 a_2_48 vss 3.13114e-17
C6190 a_2_50 vss 3.13114e-17
C6191 a_2_49 vss 3.13114e-17
C6192 a_2_81 vss 1.40901e-16
C6193 a_2_50 vss 1.40901e-16
C6194 a_2_52 vss 1.40901e-17
C6195 a_2_51 vss 1.40901e-17
C6196 a_2_53 vss 3.13114e-17
C6197 a_2_52 vss 3.13114e-17
C6198 a_2_54 vss 3.13114e-17
C6199 a_2_53 vss 3.13114e-17
C6200 a_2_55 vss 3.13114e-17
C6201 a_2_54 vss 3.13114e-17
C6202 a_2_56 vss 3.13114e-17
C6203 a_2_55 vss 3.13114e-17
C6204 a_2_57 vss 3.13114e-17
C6205 a_2_56 vss 3.13114e-17
C6206 a_2_58 vss 3.13114e-17
C6207 a_2_57 vss 3.13114e-17
C6208 a_2_59 vss 3.13114e-17
C6209 a_2_58 vss 3.13114e-17
C6210 a_2_60 vss 3.13114e-17
C6211 a_2_59 vss 3.13114e-17
C6212 a_2_61 vss 3.13114e-17
C6213 a_2_60 vss 3.13114e-17
C6214 a_2_62 vss 3.13114e-17
C6215 a_2_61 vss 3.13114e-17
C6216 a_2_63 vss 3.13114e-17
C6217 a_2_62 vss 3.13114e-17
C6218 a_2_64 vss 3.13114e-17
C6219 a_2_63 vss 3.13114e-17
C6220 a_2_65 vss 3.13114e-17
C6221 a_2_64 vss 3.13114e-17
C6222 a_2_66 vss 3.13114e-17
C6223 a_2_65 vss 3.13114e-17
C6224 a_2_67 vss 3.13114e-17
C6225 a_2_66 vss 3.13114e-17
C6226 a_2_68 vss 3.13114e-17
C6227 a_2_67 vss 3.13114e-17
C6228 a_2_69 vss 3.13114e-17
C6229 a_2_68 vss 3.13114e-17
C6230 a_2_70 vss 3.13114e-17
C6231 a_2_69 vss 3.13114e-17
C6232 a_2_71 vss 3.13114e-17
C6233 a_2_70 vss 3.13114e-17
C6234 a_2_72 vss 2.42663e-16
C6235 a_2_71 vss 2.42663e-16
C6236 a_2_73 vss 3.13114e-17
C6237 a_2_72 vss 3.13114e-17
C6238 a_2_74 vss 3.13114e-17
C6239 a_2_73 vss 3.13114e-17
C6240 a_2_75 vss 3.13114e-17
C6241 a_2_74 vss 3.13114e-17
C6242 a_2_76 vss 3.13114e-17
C6243 a_2_75 vss 3.13114e-17
C6244 a_2_77 vss 3.13114e-17
C6245 a_2_76 vss 3.13114e-17
C6246 a_2_78 vss 3.13114e-17
C6247 a_2_77 vss 3.13114e-17
C6248 a_2_79 vss 3.13114e-17
C6249 a_2_78 vss 3.13114e-17
C6250 a_2_82 vss 1.40901e-16
C6251 a_2_79 vss 1.40901e-16
C6252 a_2_82 vss 6.34418e-17
C6253 a_2_80 vss 6.34418e-17
C6254 a_2_81 vss 1.42197e-16
C6255 a_2_82 vss 1.42197e-16
C6256 a_2_83 vss 6.8969e-16
C6257 a_2_82 vss 6.8969e-16
C6258 a_2_84 vss 3.48676e-17
C6259 a_2_83 vss 3.48676e-17
C6260 a_2 vss 4.3846e-15
C6261 a_2_84 vss 4.3846e-15

R145_1 selsel_45 selsel_10 0.001
R145_2 selsel_44 selsel_20 0.001
R145_3 selsel_42 selsel_30 0.001
R145_4 selsel_43 selsel_40 0.001
R145_5 selsel_41 selsel_56 0.001
R145_6 selsel_51 selsel_60 0.001
R145_7 selsel_59 selsel_62 0.001
R145_8 selsel_7 selsel_2 0.001
R145_9 selsel_17 selsel_12 0.001
R145_10 selsel_27 selsel_22 0.001
R145_11 selsel_53 selsel_47 0.001
R145_12 selsel_1 selsel_4 0.001
R145_13 selsel_11 selsel_14 0.001
R145_14 selsel_37 selsel_31 0.001
R145_15 selsel_21 selsel_24 0.001
R145_16 selsel_32 selsel_34 0.001
R145_17 selsel_46 selsel_49 0.001
R145_18 selsel_61 selsel_89 0.001
R145_19 selsel_87 selsel_64 0.001
R145_20 selsel_84 selsel_66 0.001
R145_21 selsel_86 selsel_66 0.001
R145_22 selsel_83 selsel_66 0.001
R145_23 selsel_85 selsel_66 0.001
R145_24 selsel_72 selsel_67 0.001
R145_25 selsel_69 selsel_67 0.001
R145_26 selsel_70 selsel_67 0.001
R145_27 selsel_71 selsel_67 0.001
R145_28 selsel_73 selsel_67 0.001
R145_29 selsel_76 selsel_67 0.001
R145_30 selsel_75 selsel_67 0.001
R145_31 selsel_74 selsel_67 0.001
R145_32 selsel_79 selsel_67 0.001
R145_33 selsel_77 selsel_67 0.001
R145_34 selsel_78 selsel_67 0.001
R145_35 selsel_80 selsel_67 0.001
R145_36 selsel_81 selsel_67 0.001
R145_37 selsel_82 selsel_67 0.001
R145_38 selsel_64 selsel_63 0.001
R145_39 selsel_65 selsel_64 0.054
R145_40 selsel_69 selsel_68 0.001
R145_41 selsel_70 selsel_69 0.108
R145_42 selsel_71 selsel_70 0.108
R145_43 selsel_72 selsel_71 0.108
R145_44 selsel_73 selsel_72 0.108
R145_45 selsel_74 selsel_73 0.108
R145_46 selsel_75 selsel_74 0.108
R145_47 selsel_76 selsel_75 0.108
R145_48 selsel_77 selsel_76 0.108
R145_49 selsel_78 selsel_77 0.108
R145_50 selsel_79 selsel_78 0.108
R145_51 selsel_80 selsel_79 0.108
R145_52 selsel_81 selsel_80 0.108
R145_53 selsel_82 selsel_81 0.108
R145_54 selsel_83 selsel_82 0.864
R145_55 selsel_84 selsel_83 0.108
R145_56 selsel_85 selsel_84 0.108
R145_57 selsel_86 selsel_85 0.108
R145_58 selsel_87 selsel_86 0.54
R145_59 selsel_88 selsel_87 0.001
R145_60 selsel_89 selsel_88 9.72
R145_61 selsel_14 selsel_13 72
R145_62 selsel_15 selsel_14 43.2
R145_63 selsel_34 selsel_33 64.8
R145_64 selsel_35 selsel_34 50.4
R145_65 selsel_24 selsel_23 72
R145_66 selsel_25 selsel_24 43.2
R145_67 selsel_49 selsel_48 72
R145_68 selsel_50 selsel_49 43.2
R145_69 selsel_62 selsel_61 4.644
R145_70 selsel_4 selsel_3 72
R145_71 selsel selsel_4 43.2
R145_72 selsel_12 selsel_11 0.108
R145_73 selsel_32 selsel_31 0.324
R145_74 selsel_22 selsel_21 0.108
R145_75 selsel_60 selsel_59 2.052
R145_76 selsel_47 selsel_46 0.108
R145_77 selsel_2 selsel_1 0.108
R145_78 selsel_17 selsel_16 0.756
R145_79 selsel_18 selsel_17 0.324
R145_80 selsel_37 selsel_36 0.486
R145_81 selsel_38 selsel_37 0.648
R145_82 selsel_27 selsel_26 0.756
R145_83 selsel_28 selsel_27 0.324
R145_84 selsel_51 selsel_58 0.108
R145_85 selsel_53 selsel_52 0.756
R145_86 selsel_54 selsel_53 0.324
R145_87 selsel_19 selsel_18 0.054
R145_88 selsel_20 selsel_19 0.54
R145_89 selsel_39 selsel_38 0.054
R145_90 selsel_40 selsel_39 0.54
R145_91 selsel_29 selsel_28 0.054
R145_92 selsel_30 selsel_29 0.54
R145_93 selsel_55 selsel_54 0.054
R145_94 selsel_56 selsel_55 0.54
R145_95 selsel_57 selsel_56 0.108
R145_96 selsel_58 selsel_57 0.054
R145_97 selsel_7 selsel_6 0.756
R145_98 selsel_8 selsel_7 0.324
R145_99 selsel_9 selsel_8 0.054
R145_100 selsel_10 selsel_9 0.54
R145_101 selsel_42 selsel_41 12.528
R145_102 selsel_43 selsel_42 1.62
R145_103 selsel_44 selsel_43 9.288
R145_104 selsel_45 selsel_44 2.808

C6262 selsel_64 vss 1.30248e-17
C6263 selsel_63 vss 1.30248e-17
C6264 selsel_65 vss 1.95372e-17
C6265 selsel_64 vss 1.95372e-17
C6266 selsel_69 vss 1.40901e-17
C6267 selsel_68 vss 1.40901e-17
C6268 selsel_70 vss 3.13114e-17
C6269 selsel_69 vss 3.13114e-17
C6270 selsel_71 vss 3.13114e-17
C6271 selsel_70 vss 3.13114e-17
C6272 selsel_72 vss 3.13114e-17
C6273 selsel_71 vss 3.13114e-17
C6274 selsel_73 vss 3.13114e-17
C6275 selsel_72 vss 3.13114e-17
C6276 selsel_74 vss 3.13114e-17
C6277 selsel_73 vss 3.13114e-17
C6278 selsel_75 vss 3.13114e-17
C6279 selsel_74 vss 3.13114e-17
C6280 selsel_76 vss 3.13114e-17
C6281 selsel_75 vss 3.13114e-17
C6282 selsel_77 vss 3.13114e-17
C6283 selsel_76 vss 3.13114e-17
C6284 selsel_78 vss 3.13114e-17
C6285 selsel_77 vss 3.13114e-17
C6286 selsel_79 vss 3.13114e-17
C6287 selsel_78 vss 3.13114e-17
C6288 selsel_80 vss 3.13114e-17
C6289 selsel_79 vss 3.13114e-17
C6290 selsel_81 vss 3.13114e-17
C6291 selsel_80 vss 3.13114e-17
C6292 selsel_82 vss 3.13114e-17
C6293 selsel_81 vss 3.13114e-17
C6294 selsel_83 vss 2.42663e-16
C6295 selsel_82 vss 2.42663e-16
C6296 selsel_84 vss 3.91392e-17
C6297 selsel_83 vss 3.91392e-17
C6298 selsel_85 vss 3.91392e-17
C6299 selsel_84 vss 3.91392e-17
C6300 selsel_86 vss 3.91392e-17
C6301 selsel_85 vss 3.91392e-17
C6302 selsel_87 vss 1.64385e-16
C6303 selsel_86 vss 1.64385e-16
C6304 selsel_88 vss 2.1918e-17
C6305 selsel_87 vss 2.1918e-17
C6306 selsel_89 vss 9.79268e-16
C6307 selsel_88 vss 9.79268e-16
C6308 selsel_14 vss 8.21582e-17
C6309 selsel_13 vss 8.21582e-17
C6310 selsel_15 vss 5.086e-17
C6311 selsel_14 vss 5.086e-17
C6312 selsel_34 vss 7.43336e-17
C6313 selsel_33 vss 7.43336e-17
C6314 selsel_35 vss 5.86844e-17
C6315 selsel_34 vss 5.86844e-17
C6316 selsel_24 vss 8.21582e-17
C6317 selsel_23 vss 8.21582e-17
C6318 selsel_25 vss 5.086e-17
C6319 selsel_24 vss 5.086e-17
C6320 selsel_49 vss 8.21582e-17
C6321 selsel_48 vss 8.21582e-17
C6322 selsel_50 vss 5.086e-17
C6323 selsel_49 vss 5.086e-17
C6324 selsel_62 vss 1.05883e-15
C6325 selsel_61 vss 1.05883e-15
C6326 selsel_4 vss 8.21582e-17
C6327 selsel_3 vss 8.21582e-17
C6328 selsel vss 5.086e-17
C6329 selsel_4 vss 5.086e-17
C6330 selsel_12 vss 3.65472e-17
C6331 selsel_11 vss 3.65472e-17
C6332 selsel_32 vss 3.39552e-17
C6333 selsel_31 vss 3.39552e-17
C6334 selsel_22 vss 3.65472e-17
C6335 selsel_21 vss 3.65472e-17
C6336 selsel_60 vss 2.10522e-16
C6337 selsel_59 vss 2.10522e-16
C6338 selsel_47 vss 3.65472e-17
C6339 selsel_46 vss 3.65472e-17
C6340 selsel_2 vss 3.65472e-17
C6341 selsel_1 vss 3.65472e-17
C6342 selsel_17 vss 1.78524e-16
C6343 selsel_16 vss 1.78524e-16
C6344 selsel_18 vss 8.0028e-17
C6345 selsel_17 vss 8.0028e-17
C6346 selsel_37 vss 1.10808e-16
C6347 selsel_36 vss 1.10808e-16
C6348 selsel_38 vss 1.47744e-16
C6349 selsel_37 vss 1.47744e-16
C6350 selsel_27 vss 1.78524e-16
C6351 selsel_26 vss 1.78524e-16
C6352 selsel_28 vss 8.0028e-17
C6353 selsel_27 vss 8.0028e-17
C6354 selsel_51 vss 2.4624e-17
C6355 selsel_58 vss 2.4624e-17
C6356 selsel_53 vss 1.78524e-16
C6357 selsel_52 vss 1.78524e-16
C6358 selsel_54 vss 8.0028e-17
C6359 selsel_53 vss 8.0028e-17
C6360 selsel_19 vss 1.2312e-17
C6361 selsel_18 vss 1.2312e-17
C6362 selsel_20 vss 1.2312e-16
C6363 selsel_19 vss 1.2312e-16
C6364 selsel_39 vss 1.2312e-17
C6365 selsel_38 vss 1.2312e-17
C6366 selsel_40 vss 1.2312e-16
C6367 selsel_39 vss 1.2312e-16
C6368 selsel_29 vss 1.2312e-17
C6369 selsel_28 vss 1.2312e-17
C6370 selsel_30 vss 1.2312e-16
C6371 selsel_29 vss 1.2312e-16
C6372 selsel_55 vss 1.2312e-17
C6373 selsel_54 vss 1.2312e-17
C6374 selsel_56 vss 1.2312e-16
C6375 selsel_55 vss 1.2312e-16
C6376 selsel_57 vss 3.078e-17
C6377 selsel_56 vss 3.078e-17
C6378 selsel_58 vss 1.2312e-17
C6379 selsel_57 vss 1.2312e-17
C6380 selsel_7 vss 1.78524e-16
C6381 selsel_6 vss 1.78524e-16
C6382 selsel_8 vss 8.0028e-17
C6383 selsel_7 vss 8.0028e-17
C6384 selsel_9 vss 1.2312e-17
C6385 selsel_8 vss 1.2312e-17
C6386 selsel_10 vss 1.2312e-16
C6387 selsel_9 vss 1.2312e-16
C6388 selsel_42 vss 1.26313e-15
C6389 selsel_41 vss 1.26313e-15
C6390 selsel_43 vss 1.62985e-16
C6391 selsel_42 vss 1.62985e-16
C6392 selsel_44 vss 9.37163e-16
C6393 selsel_43 vss 9.37163e-16
C6394 selsel_45 vss 2.85224e-16
C6395 selsel_44 vss 2.85224e-16

R146_1 ss_1_16 ss_1_2 0.001
R146_2 ss_1_15 ss_1_29 0.001
R146_3 ss_1_26 ss_1_31 0.001
R146_4 ss_1_23 ss_1_17 0.001
R146_5 ss_1_18 ss_1_21 0.001
R146_6 ss_1_30 ss_1_36 0.001
R146_7 ss_1_33 ss_1_42 0.001
R146_8 ss_1_40 ss_1_37 0.001
R146_9 ss_1_41 ss_1_37 0.001
R146_10 ss_1_39 ss_1_38 0.001
R146_11 ss_1_1 ss_1_4 0.001
R146_12 ss_1_3 ss_1_6 0.001
R146_13 ss_1_5 ss_1_8 0.001
R146_14 ss_1_7 ss_1_10 0.001
R146_15 ss_1_9 ss_1_14 0.001
R146_16 ss_1_13 ss_1_12 0.001
R146_17 ss_1_12 ss_1_11 475.2
R146_18 ss_1_39 ss_1_43 0.324
R146_19 ss_1_14 ss_1_13 0.324
R146_20 ss_1_41 ss_1_40 0.216
R146_21 ss_1_42 ss_1_41 0.216
R146_22 ss_1_43 ss_1_42 0.108
R146_23 ss_1_10 ss_1_9 0.162
R146_24 ss_1 ss_1_21 50.4
R146_25 ss_1_21 ss_1_20 108
R146_26 ss_1_33 ss_1_32 0.648
R146_27 ss_1_34 ss_1_33 0.486
R146_28 ss_1_35 ss_1_34 0.054
R146_29 ss_1_36 ss_1_35 0.108
R146_30 ss_1_8 ss_1_7 0.864
R146_31 ss_1_18 ss_1_17 0.216
R146_32 ss_1_31 ss_1_30 7.668
R146_33 ss_1_6 ss_1_5 5.94
R146_34 ss_1_23 ss_1_22 0.594
R146_35 ss_1_24 ss_1_23 0.486
R146_36 ss_1_25 ss_1_24 0.054
R146_37 ss_1_26 ss_1_25 0.108
R146_38 ss_1_27 ss_1_26 0.54
R146_39 ss_1_4 ss_1_3 37.044
R146_40 ss_1_28 ss_1_27 0.054
R146_41 ss_1_29 ss_1_28 0.108
R146_42 ss_1_2 ss_1_1 4.86
R146_43 ss_1_16 ss_1_15 0.54

C6396 ss_1_12 vss 5.18379e-16
C6397 ss_1_11 vss 5.18379e-16
C6398 ss_1_39 vss 4.07462e-17
C6399 ss_1_43 vss 4.07462e-17
C6400 ss_1_14 vss 7.30944e-17
C6401 ss_1_13 vss 7.30944e-17
C6402 ss_1_41 vss 4.38566e-17
C6403 ss_1_40 vss 4.38566e-17
C6404 ss_1_42 vss 4.38566e-17
C6405 ss_1_41 vss 4.38566e-17
C6406 ss_1_43 vss 3.65472e-17
C6407 ss_1_42 vss 3.65472e-17
C6408 ss_1_10 vss 6.5124e-17
C6409 ss_1_9 vss 6.5124e-17
C6410 ss_1 vss 5.86844e-17
C6411 ss_1_21 vss 5.86844e-17
C6412 ss_1_21 vss 1.21281e-16
C6413 ss_1_20 vss 1.21281e-16
C6414 ss_1_33 vss 1.47744e-16
C6415 ss_1_32 vss 1.47744e-16
C6416 ss_1_34 vss 1.10808e-16
C6417 ss_1_33 vss 1.10808e-16
C6418 ss_1_35 vss 1.2312e-17
C6419 ss_1_34 vss 1.2312e-17
C6420 ss_1_36 vss 3.078e-17
C6421 ss_1_35 vss 3.078e-17
C6422 ss_1_8 vss 1.53498e-16
C6423 ss_1_7 vss 1.53498e-16
C6424 ss_1_18 vss 2.71642e-17
C6425 ss_1_17 vss 2.71642e-17
C6426 ss_1_31 vss 7.74179e-16
C6427 ss_1_30 vss 7.74179e-16
C6428 ss_1_6 vss 2.14909e-15
C6429 ss_1_5 vss 2.14909e-15
C6430 ss_1_23 vss 1.41588e-16
C6431 ss_1_22 vss 1.41588e-16
C6432 ss_1_24 vss 1.16964e-16
C6433 ss_1_23 vss 1.16964e-16
C6434 ss_1_25 vss 1.2312e-17
C6435 ss_1_24 vss 1.2312e-17
C6436 ss_1_26 vss 3.078e-17
C6437 ss_1_25 vss 3.078e-17
C6438 ss_1_27 vss 1.2312e-16
C6439 ss_1_26 vss 1.2312e-16
C6440 ss_1_4 vss 3.72828e-15
C6441 ss_1_3 vss 3.72828e-15
C6442 ss_1_28 vss 1.2312e-17
C6443 ss_1_27 vss 1.2312e-17
C6444 ss_1_29 vss 2.4624e-17
C6445 ss_1_28 vss 2.4624e-17
C6446 ss_1_2 vss 1.10808e-15
C6447 ss_1_1 vss 1.10808e-15
C6448 ss_1_16 vss 5.43283e-17
C6449 ss_1_15 vss 5.43283e-17

R147_1 aa_3_2 aa_3_18 0.001
R147_2 aa_3_1 aa_3_14 0.001
R147_3 aa_3_9 aa_3_4 0.001
R147_4 aa_3_3 aa_3_6 0.001
R147_5 aa_3_16 aa_3_22 0.001
R147_6 aa_3_17 aa_3_15 0.001
R147_7 aa_3_29 aa_3_19 0.001
R147_8 aa_3_31 aa_3_19 0.001
R147_9 aa_3_32 aa_3_19 0.001
R147_10 aa_3_30 aa_3_19 0.001
R147_11 aa_3_36 aa_3_20 0.001
R147_12 aa_3_34 aa_3_20 0.001
R147_13 aa_3_33 aa_3_20 0.001
R147_14 aa_3_38 aa_3_20 0.001
R147_15 aa_3_37 aa_3_20 0.001
R147_16 aa_3_35 aa_3_20 0.001
R147_17 aa_3_39 aa_3_20 0.001
R147_18 aa_3_40 aa_3_20 0.001
R147_19 aa_3_41 aa_3_20 0.001
R147_20 aa_3_46 aa_3_20 0.001
R147_21 aa_3_45 aa_3_20 0.001
R147_22 aa_3_44 aa_3_20 0.001
R147_23 aa_3_43 aa_3_20 0.001
R147_24 aa_3_42 aa_3_20 0.001
R147_25 aa_3_21 aa_3_26 0.001
R147_26 aa_3_28 aa_3_24 0.001
R147_27 aa_3_24 aa_3_23 0.054
R147_28 aa_3_25 aa_3_24 0.001
R147_29 aa_3_29 aa_3_28 0.54
R147_30 aa_3_30 aa_3_29 0.108
R147_31 aa_3_31 aa_3_30 0.108
R147_32 aa_3_32 aa_3_31 0.108
R147_33 aa_3_33 aa_3_32 0.864
R147_34 aa_3_34 aa_3_33 0.108
R147_35 aa_3_35 aa_3_34 0.108
R147_36 aa_3_36 aa_3_35 0.108
R147_37 aa_3_37 aa_3_36 0.108
R147_38 aa_3_38 aa_3_37 0.108
R147_39 aa_3_39 aa_3_38 0.108
R147_40 aa_3_40 aa_3_39 0.108
R147_41 aa_3_41 aa_3_40 0.108
R147_42 aa_3_42 aa_3_41 0.108
R147_43 aa_3_43 aa_3_42 0.108
R147_44 aa_3_44 aa_3_43 0.108
R147_45 aa_3_45 aa_3_44 0.108
R147_46 aa_3_46 aa_3_45 0.108
R147_47 aa_3_47 aa_3_46 0.001
R147_48 aa_3_6 aa_3_5 72
R147_49 aa_3 aa_3_6 43.2
R147_50 aa_3_27 aa_3_26 0.864
R147_51 aa_3_28 aa_3_27 0.001
R147_52 aa_3_22 aa_3_21 2.484
R147_53 aa_3_4 aa_3_3 0.108
R147_54 aa_3_16 aa_3_15 9.72
R147_55 aa_3_9 aa_3_8 0.756
R147_56 aa_3_10 aa_3_9 0.324
R147_57 aa_3_11 aa_3_10 0.054
R147_58 aa_3_12 aa_3_11 0.648
R147_59 aa_3_18 aa_3_17 4.59
R147_60 aa_3_13 aa_3_12 0.054
R147_61 aa_3_14 aa_3_13 0.216
R147_62 aa_3_2 aa_3_1 35.208

C6450 aa_3_24 vss 1.95372e-17
C6451 aa_3_23 vss 1.95372e-17
C6452 aa_3_25 vss 1.30248e-17
C6453 aa_3_24 vss 1.30248e-17
C6454 aa_3_29 vss 1.64385e-16
C6455 aa_3_28 vss 1.64385e-16
C6456 aa_3_30 vss 3.91392e-17
C6457 aa_3_29 vss 3.91392e-17
C6458 aa_3_31 vss 3.91392e-17
C6459 aa_3_30 vss 3.91392e-17
C6460 aa_3_32 vss 3.91392e-17
C6461 aa_3_31 vss 3.91392e-17
C6462 aa_3_33 vss 2.42663e-16
C6463 aa_3_32 vss 2.42663e-16
C6464 aa_3_34 vss 3.13114e-17
C6465 aa_3_33 vss 3.13114e-17
C6466 aa_3_35 vss 3.13114e-17
C6467 aa_3_34 vss 3.13114e-17
C6468 aa_3_36 vss 3.13114e-17
C6469 aa_3_35 vss 3.13114e-17
C6470 aa_3_37 vss 3.13114e-17
C6471 aa_3_36 vss 3.13114e-17
C6472 aa_3_38 vss 3.13114e-17
C6473 aa_3_37 vss 3.13114e-17
C6474 aa_3_39 vss 3.13114e-17
C6475 aa_3_38 vss 3.13114e-17
C6476 aa_3_40 vss 3.13114e-17
C6477 aa_3_39 vss 3.13114e-17
C6478 aa_3_41 vss 3.13114e-17
C6479 aa_3_40 vss 3.13114e-17
C6480 aa_3_42 vss 3.13114e-17
C6481 aa_3_41 vss 3.13114e-17
C6482 aa_3_43 vss 3.13114e-17
C6483 aa_3_42 vss 3.13114e-17
C6484 aa_3_44 vss 3.13114e-17
C6485 aa_3_43 vss 3.13114e-17
C6486 aa_3_45 vss 3.13114e-17
C6487 aa_3_44 vss 3.13114e-17
C6488 aa_3_46 vss 3.13114e-17
C6489 aa_3_45 vss 3.13114e-17
C6490 aa_3_47 vss 1.40901e-17
C6491 aa_3_46 vss 1.40901e-17
C6492 aa_3_6 vss 8.21582e-17
C6493 aa_3_5 vss 8.21582e-17
C6494 aa_3 vss 5.086e-17
C6495 aa_3_6 vss 5.086e-17
C6496 aa_3_27 vss 9.64328e-17
C6497 aa_3_26 vss 9.64328e-17
C6498 aa_3_28 vss 2.1918e-17
C6499 aa_3_27 vss 2.1918e-17
C6500 aa_3_22 vss 5.72508e-16
C6501 aa_3_21 vss 5.72508e-16
C6502 aa_3_4 vss 3.65472e-17
C6503 aa_3_3 vss 3.65472e-17
C6504 aa_3_16 vss 9.84701e-16
C6505 aa_3_15 vss 9.84701e-16
C6506 aa_3_9 vss 1.78524e-16
C6507 aa_3_8 vss 1.78524e-16
C6508 aa_3_10 vss 8.0028e-17
C6509 aa_3_9 vss 8.0028e-17
C6510 aa_3_11 vss 1.2312e-17
C6511 aa_3_10 vss 1.2312e-17
C6512 aa_3_12 vss 1.539e-16
C6513 aa_3_11 vss 1.539e-16
C6514 aa_3_18 vss 1.04652e-15
C6515 aa_3_17 vss 1.04652e-15
C6516 aa_3_13 vss 1.2312e-17
C6517 aa_3_12 vss 1.2312e-17
C6518 aa_3_14 vss 5.5404e-17
C6519 aa_3_13 vss 5.5404e-17
C6520 aa_3_2 vss 3.55171e-15
C6521 aa_3_1 vss 3.55171e-15

R148_1 aa_2_2 aa_2_21 0.001
R148_2 aa_2_1 aa_2_14 0.001
R148_3 aa_2_9 aa_2_4 0.001
R148_4 aa_2_3 aa_2_6 0.001
R148_5 aa_2_34 aa_2_15 0.001
R148_6 aa_2_33 aa_2_15 0.001
R148_7 aa_2_31 aa_2_15 0.001
R148_8 aa_2_32 aa_2_15 0.001
R148_9 aa_2_30 aa_2_15 0.001
R148_10 aa_2_29 aa_2_15 0.001
R148_11 aa_2_38 aa_2_15 0.001
R148_12 aa_2_35 aa_2_15 0.001
R148_13 aa_2_36 aa_2_15 0.001
R148_14 aa_2_37 aa_2_15 0.001
R148_15 aa_2_42 aa_2_15 0.001
R148_16 aa_2_41 aa_2_15 0.001
R148_17 aa_2_40 aa_2_15 0.001
R148_18 aa_2_39 aa_2_15 0.001
R148_19 aa_2_25 aa_2_19 0.001
R148_20 aa_2_24 aa_2_17 0.001
R148_21 aa_2_26 aa_2_19 0.001
R148_22 aa_2_27 aa_2_19 0.001
R148_23 aa_2_28 aa_2_19 0.001
R148_24 aa_2_20 aa_2_22 0.001
R148_25 aa_2_6 aa_2_5 72
R148_26 aa_2 aa_2_6 43.2
R148_27 aa_2_17 aa_2_16 0.054
R148_28 aa_2_18 aa_2_17 0.001
R148_29 aa_2_4 aa_2_3 0.108
R148_30 aa_2_25 aa_2_24 0.54
R148_31 aa_2_26 aa_2_25 0.108
R148_32 aa_2_27 aa_2_26 0.108
R148_33 aa_2_28 aa_2_27 0.108
R148_34 aa_2_29 aa_2_28 0.864
R148_35 aa_2_30 aa_2_29 0.108
R148_36 aa_2_31 aa_2_30 0.108
R148_37 aa_2_32 aa_2_31 0.108
R148_38 aa_2_33 aa_2_32 0.108
R148_39 aa_2_34 aa_2_33 0.108
R148_40 aa_2_35 aa_2_34 0.108
R148_41 aa_2_36 aa_2_35 0.108
R148_42 aa_2_37 aa_2_36 0.108
R148_43 aa_2_38 aa_2_37 0.108
R148_44 aa_2_39 aa_2_38 0.108
R148_45 aa_2_40 aa_2_39 0.108
R148_46 aa_2_41 aa_2_40 0.108
R148_47 aa_2_42 aa_2_41 0.108
R148_48 aa_2_43 aa_2_42 0.001
R148_49 aa_2_23 aa_2_22 10.368
R148_50 aa_2_24 aa_2_23 0.001
R148_51 aa_2_9 aa_2_8 0.756
R148_52 aa_2_10 aa_2_9 0.324
R148_53 aa_2_11 aa_2_10 0.054
R148_54 aa_2_12 aa_2_11 0.648
R148_55 aa_2_21 aa_2_20 2.592
R148_56 aa_2_13 aa_2_12 0.054
R148_57 aa_2_14 aa_2_13 0.378
R148_58 aa_2_2 aa_2_1 23.004

C6522 aa_2_6 vss 8.21582e-17
C6523 aa_2_5 vss 8.21582e-17
C6524 aa_2 vss 5.086e-17
C6525 aa_2_6 vss 5.086e-17
C6526 aa_2_17 vss 1.95372e-17
C6527 aa_2_16 vss 1.95372e-17
C6528 aa_2_18 vss 1.30248e-17
C6529 aa_2_17 vss 1.30248e-17
C6530 aa_2_4 vss 3.65472e-17
C6531 aa_2_3 vss 3.65472e-17
C6532 aa_2_25 vss 1.64385e-16
C6533 aa_2_24 vss 1.64385e-16
C6534 aa_2_26 vss 3.91392e-17
C6535 aa_2_25 vss 3.91392e-17
C6536 aa_2_27 vss 3.91392e-17
C6537 aa_2_26 vss 3.91392e-17
C6538 aa_2_28 vss 3.91392e-17
C6539 aa_2_27 vss 3.91392e-17
C6540 aa_2_29 vss 2.42663e-16
C6541 aa_2_28 vss 2.42663e-16
C6542 aa_2_30 vss 3.13114e-17
C6543 aa_2_29 vss 3.13114e-17
C6544 aa_2_31 vss 3.13114e-17
C6545 aa_2_30 vss 3.13114e-17
C6546 aa_2_32 vss 3.13114e-17
C6547 aa_2_31 vss 3.13114e-17
C6548 aa_2_33 vss 3.13114e-17
C6549 aa_2_32 vss 3.13114e-17
C6550 aa_2_34 vss 3.13114e-17
C6551 aa_2_33 vss 3.13114e-17
C6552 aa_2_35 vss 3.13114e-17
C6553 aa_2_34 vss 3.13114e-17
C6554 aa_2_36 vss 3.13114e-17
C6555 aa_2_35 vss 3.13114e-17
C6556 aa_2_37 vss 3.13114e-17
C6557 aa_2_36 vss 3.13114e-17
C6558 aa_2_38 vss 3.13114e-17
C6559 aa_2_37 vss 3.13114e-17
C6560 aa_2_39 vss 3.13114e-17
C6561 aa_2_38 vss 3.13114e-17
C6562 aa_2_40 vss 3.13114e-17
C6563 aa_2_39 vss 3.13114e-17
C6564 aa_2_41 vss 3.13114e-17
C6565 aa_2_40 vss 3.13114e-17
C6566 aa_2_42 vss 3.13114e-17
C6567 aa_2_41 vss 3.13114e-17
C6568 aa_2_43 vss 1.40901e-17
C6569 aa_2_42 vss 1.40901e-17
C6570 aa_2_23 vss 1.04718e-15
C6571 aa_2_22 vss 1.04718e-15
C6572 aa_2_24 vss 2.1918e-17
C6573 aa_2_23 vss 2.1918e-17
C6574 aa_2_9 vss 1.78524e-16
C6575 aa_2_8 vss 1.78524e-16
C6576 aa_2_10 vss 8.0028e-17
C6577 aa_2_9 vss 8.0028e-17
C6578 aa_2_11 vss 1.2312e-17
C6579 aa_2_10 vss 1.2312e-17
C6580 aa_2_12 vss 1.539e-16
C6581 aa_2_11 vss 1.539e-16
C6582 aa_2_21 vss 5.90976e-16
C6583 aa_2_20 vss 5.90976e-16
C6584 aa_2_13 vss 1.2312e-17
C6585 aa_2_12 vss 1.2312e-17
C6586 aa_2_14 vss 8.6184e-17
C6587 aa_2_13 vss 8.6184e-17
C6588 aa_2_2 vss 2.32254e-15
C6589 aa_2_1 vss 2.32254e-15

R149_1 ss_3_2 ss_3_28 0.001
R149_2 ss_3_10 ss_3_1 0.001
R149_3 ss_3_4 ss_3_7 0.001
R149_4 ss_3_8 ss_3_5 0.001
R149_5 ss_3_6 ss_3_14 0.001
R149_6 ss_3_12 ss_3_9 0.001
R149_7 ss_3_13 ss_3_11 0.001
R149_8 ss_3_23 ss_3_15 0.001
R149_9 ss_3_16 ss_3_19 0.001
R149_10 ss_3_20 ss_3_30 0.001
R149_11 ss_3_29 ss_3_35 0.001
R149_12 ss_3_32 ss_3_41 0.001
R149_13 ss_3_39 ss_3_36 0.001
R149_14 ss_3_40 ss_3_36 0.001
R149_15 ss_3_38 ss_3_37 0.001
R149_16 ss_3_38 ss_3_42 0.324
R149_17 ss_3_40 ss_3_39 0.216
R149_18 ss_3_41 ss_3_40 0.216
R149_19 ss_3_42 ss_3_41 0.108
R149_20 ss_3_32 ss_3_31 0.648
R149_21 ss_3_33 ss_3_32 0.486
R149_22 ss_3_34 ss_3_33 0.054
R149_23 ss_3_35 ss_3_34 0.27
R149_24 ss_3 ss_3_19 50.4
R149_25 ss_3_19 ss_3_18 108
R149_26 ss_3_30 ss_3_29 3.996
R149_27 ss_3_16 ss_3_15 0.216
R149_28 ss_3_21 ss_3_20 0.81
R149_29 ss_3_22 ss_3_21 0.054
R149_30 ss_3_23 ss_3_22 0.54
R149_31 ss_3_24 ss_3_23 0.486
R149_32 ss_3_25 ss_3_24 0.054
R149_33 ss_3_26 ss_3_25 0.648
R149_34 ss_3_27 ss_3_26 0.054
R149_35 ss_3_28 ss_3_27 0.378
R149_36 ss_3_2 ss_3_1 8.424
R149_37 ss_3_10 ss_3_9 0.648
R149_38 ss_3_12 ss_3_11 5.184
R149_39 ss_3_14 ss_3_13 1.35
R149_40 ss_3_6 ss_3_8 0.54
R149_41 ss_3_4 ss_3_3 475.2
R149_42 ss_3_8 ss_3_7 0.324

C6590 ss_3_38 vss 4.07462e-17
C6591 ss_3_42 vss 4.07462e-17
C6592 ss_3_40 vss 4.38566e-17
C6593 ss_3_39 vss 4.38566e-17
C6594 ss_3_41 vss 4.38566e-17
C6595 ss_3_40 vss 4.38566e-17
C6596 ss_3_42 vss 3.65472e-17
C6597 ss_3_41 vss 3.65472e-17
C6598 ss_3_32 vss 1.47744e-16
C6599 ss_3_31 vss 1.47744e-16
C6600 ss_3_33 vss 1.10808e-16
C6601 ss_3_32 vss 1.10808e-16
C6602 ss_3_34 vss 1.2312e-17
C6603 ss_3_33 vss 1.2312e-17
C6604 ss_3_35 vss 6.156e-17
C6605 ss_3_34 vss 6.156e-17
C6606 ss_3 vss 5.86844e-17
C6607 ss_3_19 vss 5.86844e-17
C6608 ss_3_19 vss 1.21281e-16
C6609 ss_3_18 vss 1.21281e-16
C6610 ss_3_30 vss 4.07462e-16
C6611 ss_3_29 vss 4.07462e-16
C6612 ss_3_16 vss 2.71642e-17
C6613 ss_3_15 vss 2.71642e-17
C6614 ss_3_21 vss 1.8468e-16
C6615 ss_3_20 vss 1.8468e-16
C6616 ss_3_22 vss 1.2312e-17
C6617 ss_3_21 vss 1.2312e-17
C6618 ss_3_23 vss 1.29276e-16
C6619 ss_3_22 vss 1.29276e-16
C6620 ss_3_24 vss 1.16964e-16
C6621 ss_3_23 vss 1.16964e-16
C6622 ss_3_25 vss 1.2312e-17
C6623 ss_3_24 vss 1.2312e-17
C6624 ss_3_26 vss 1.539e-16
C6625 ss_3_25 vss 1.539e-16
C6626 ss_3_27 vss 1.2312e-17
C6627 ss_3_26 vss 1.2312e-17
C6628 ss_3_28 vss 8.6184e-17
C6629 ss_3_27 vss 8.6184e-17
C6630 ss_3_2 vss 8.55671e-16
C6631 ss_3_1 vss 8.55671e-16
C6632 ss_3_10 vss 1.539e-16
C6633 ss_3_9 vss 1.539e-16
C6634 ss_3_12 vss 9.1368e-16
C6635 ss_3_11 vss 9.1368e-16
C6636 ss_3_14 vss 3.078e-16
C6637 ss_3_13 vss 3.078e-16
C6638 ss_3_6 vss 1.09642e-16
C6639 ss_3_8 vss 1.09642e-16
C6640 ss_3_4 vss 5.18379e-16
C6641 ss_3_3 vss 5.18379e-16
C6642 ss_3_8 vss 7.30944e-17
C6643 ss_3_7 vss 7.30944e-17

R150_1 n4533 n4533_26 0.001
R150_2 n4533 n4533_27 0.001
R150_3 n4533 n4533_28 0.001
R150_4 n4533 n4533_24 0.001
R150_5 n4533 n4533_25 0.001
R150_6 n4533 n4533_23 0.001
R150_7 n4533 n4533_22 0.001
R150_8 n4533_20 n4533_2 0.001
R150_9 n4533_16 n4533_2 0.001
R150_10 n4533_17 n4533_2 0.001
R150_11 n4533_18 n4533_2 0.001
R150_12 n4533_19 n4533_2 0.001
R150_13 n4533_13 n4533_2 0.001
R150_14 n4533_15 n4533_2 0.001
R150_15 n4533_14 n4533_2 0.001
R150_16 n4533_10 n4533_2 0.001
R150_17 n4533_12 n4533_2 0.001
R150_18 n4533_11 n4533_2 0.001
R150_19 n4533_7 n4533_2 0.001
R150_20 n4533_8 n4533_2 0.001
R150_21 n4533_6 n4533_2 0.001
R150_22 n4533_9 n4533_2 0.001
R150_23 n4533_21 n4533_5 0.001
R150_24 n4533_3 n4533_4 453.6
R150_25 n4533_5 n4533_4 14.4
R150_26 n4533_7 n4533_6 0.108
R150_27 n4533_8 n4533_7 0.108
R150_28 n4533_9 n4533_8 0.108
R150_29 n4533_10 n4533_9 0.108
R150_30 n4533_11 n4533_10 0.108
R150_31 n4533_12 n4533_11 0.108
R150_32 n4533_13 n4533_12 0.108
R150_33 n4533_14 n4533_13 0.108
R150_34 n4533_15 n4533_14 0.108
R150_35 n4533_16 n4533_15 0.108
R150_36 n4533_17 n4533_16 0.108
R150_37 n4533_18 n4533_17 0.108
R150_38 n4533_19 n4533_18 0.108
R150_39 n4533_20 n4533_19 0.108
R150_40 n4533_21 n4533_20 0.108
R150_41 n4533_22 n4533_21 0.756
R150_42 n4533_23 n4533_22 0.108
R150_43 n4533_24 n4533_23 0.108
R150_44 n4533_25 n4533_24 0.108
R150_45 n4533_26 n4533_25 0.108
R150_46 n4533_27 n4533_26 0.108
R150_47 n4533_28 n4533_27 0.108

C6644 n4533_3 vss 4.98819e-16
C6645 n4533_4 vss 4.98819e-16
C6646 n4533_5 vss 8.41104e-17
C6647 n4533_4 vss 8.41104e-17
C6648 n4533_7 vss 2.92378e-17
C6649 n4533_6 vss 2.92378e-17
C6650 n4533_8 vss 2.92378e-17
C6651 n4533_7 vss 2.92378e-17
C6652 n4533_9 vss 2.92378e-17
C6653 n4533_8 vss 2.92378e-17
C6654 n4533_10 vss 2.92378e-17
C6655 n4533_9 vss 2.92378e-17
C6656 n4533_11 vss 2.92378e-17
C6657 n4533_10 vss 2.92378e-17
C6658 n4533_12 vss 2.92378e-17
C6659 n4533_11 vss 2.92378e-17
C6660 n4533_13 vss 2.92378e-17
C6661 n4533_12 vss 2.92378e-17
C6662 n4533_14 vss 2.92378e-17
C6663 n4533_13 vss 2.92378e-17
C6664 n4533_15 vss 2.92378e-17
C6665 n4533_14 vss 2.92378e-17
C6666 n4533_16 vss 2.92378e-17
C6667 n4533_15 vss 2.92378e-17
C6668 n4533_17 vss 2.92378e-17
C6669 n4533_16 vss 2.92378e-17
C6670 n4533_18 vss 2.92378e-17
C6671 n4533_17 vss 2.92378e-17
C6672 n4533_19 vss 2.92378e-17
C6673 n4533_18 vss 2.92378e-17
C6674 n4533_20 vss 2.92378e-17
C6675 n4533_19 vss 2.92378e-17
C6676 n4533_21 vss 3.65472e-17
C6677 n4533_20 vss 3.65472e-17
C6678 n4533_22 vss 1.46189e-16
C6679 n4533_21 vss 1.46189e-16
C6680 n4533_23 vss 2.92378e-17
C6681 n4533_22 vss 2.92378e-17
C6682 n4533_24 vss 2.92378e-17
C6683 n4533_23 vss 2.92378e-17
C6684 n4533_25 vss 2.92378e-17
C6685 n4533_24 vss 2.92378e-17
C6686 n4533_26 vss 2.92378e-17
C6687 n4533_25 vss 2.92378e-17
C6688 n4533_27 vss 2.92378e-17
C6689 n4533_26 vss 2.92378e-17
C6690 n4533_28 vss 2.92378e-17
C6691 n4533_27 vss 2.92378e-17

R151_1 n4572 n4572_37 0.001
R151_2 n4572 n4572_35 0.001
R151_3 n4572 n4572_36 0.001
R151_4 n4572 n4572_33 0.001
R151_5 n4572 n4572_32 0.001
R151_6 n4572 n4572_31 0.001
R151_7 n4572 n4572_34 0.001
R151_8 n4572_29 n4572_2 0.001
R151_9 n4572_26 n4572_2 0.001
R151_10 n4572_25 n4572_2 0.001
R151_11 n4572_28 n4572_2 0.001
R151_12 n4572_27 n4572_2 0.001
R151_13 n4572_23 n4572_2 0.001
R151_14 n4572_24 n4572_2 0.001
R151_15 n4572_22 n4572_2 0.001
R151_16 n4572_21 n4572_2 0.001
R151_17 n4572_19 n4572_2 0.001
R151_18 n4572_20 n4572_2 0.001
R151_19 n4572_16 n4572_2 0.001
R151_20 n4572_15 n4572_2 0.001
R151_21 n4572_18 n4572_2 0.001
R151_22 n4572_17 n4572_2 0.001
R151_23 n4572_14 n4572_12 0.001
R151_24 n4572_4 n4572_3 43.2
R151_25 n4572_11 n4572_4 21.6
R151_26 n4572_5 n4572_11 21.6
R151_27 n4572_6 n4572_5 43.2
R151_28 n4572_8 n4572_7 43.2
R151_29 n4572_13 n4572_8 21.6
R151_30 n4572_9 n4572_13 21.6
R151_31 n4572_10 n4572_9 43.2
R151_32 n4572_12 n4572_11 28.8
R151_33 n4572_13 n4572_12 28.8
R151_34 n4572_30 n4572_14 0.648
R151_35 n4572_16 n4572_15 0.108
R151_36 n4572_17 n4572_16 0.108
R151_37 n4572_18 n4572_17 0.108
R151_38 n4572_19 n4572_18 0.108
R151_39 n4572_20 n4572_19 0.108
R151_40 n4572_21 n4572_20 0.108
R151_41 n4572_22 n4572_21 0.108
R151_42 n4572_23 n4572_22 0.108
R151_43 n4572_24 n4572_23 0.108
R151_44 n4572_25 n4572_24 0.108
R151_45 n4572_26 n4572_25 0.108
R151_46 n4572_27 n4572_26 0.108
R151_47 n4572_28 n4572_27 0.108
R151_48 n4572_29 n4572_28 0.108
R151_49 n4572_30 n4572_29 0.432
R151_50 n4572_31 n4572_30 0.54
R151_51 n4572_32 n4572_31 0.108
R151_52 n4572_33 n4572_32 0.108
R151_53 n4572_34 n4572_33 0.108
R151_54 n4572_35 n4572_34 0.108
R151_55 n4572_36 n4572_35 0.108
R151_56 n4572_37 n4572_36 0.108

C6692 n4572_4 vss 4.69476e-17
C6693 n4572_3 vss 4.69476e-17
C6694 n4572_11 vss 2.34738e-17
C6695 n4572_4 vss 2.34738e-17
C6696 n4572_5 vss 2.34738e-17
C6697 n4572_11 vss 2.34738e-17
C6698 n4572_6 vss 4.69476e-17
C6699 n4572_5 vss 4.69476e-17
C6700 n4572_8 vss 4.69476e-17
C6701 n4572_7 vss 4.69476e-17
C6702 n4572_13 vss 2.34738e-17
C6703 n4572_8 vss 2.34738e-17
C6704 n4572_9 vss 2.34738e-17
C6705 n4572_13 vss 2.34738e-17
C6706 n4572_10 vss 4.69476e-17
C6707 n4572_9 vss 4.69476e-17
C6708 n4572_12 vss 7.33536e-17
C6709 n4572_11 vss 7.33536e-17
C6710 n4572_13 vss 8.25228e-17
C6711 n4572_12 vss 8.25228e-17
C6712 n4572_30 vss 1.3157e-16
C6713 n4572_14 vss 1.3157e-16
C6714 n4572_16 vss 2.92378e-17
C6715 n4572_15 vss 2.92378e-17
C6716 n4572_17 vss 2.92378e-17
C6717 n4572_16 vss 2.92378e-17
C6718 n4572_18 vss 2.92378e-17
C6719 n4572_17 vss 2.92378e-17
C6720 n4572_19 vss 2.92378e-17
C6721 n4572_18 vss 2.92378e-17
C6722 n4572_20 vss 2.92378e-17
C6723 n4572_19 vss 2.92378e-17
C6724 n4572_21 vss 2.92378e-17
C6725 n4572_20 vss 2.92378e-17
C6726 n4572_22 vss 2.92378e-17
C6727 n4572_21 vss 2.92378e-17
C6728 n4572_23 vss 2.92378e-17
C6729 n4572_22 vss 2.92378e-17
C6730 n4572_24 vss 2.92378e-17
C6731 n4572_23 vss 2.92378e-17
C6732 n4572_25 vss 2.92378e-17
C6733 n4572_24 vss 2.92378e-17
C6734 n4572_26 vss 2.92378e-17
C6735 n4572_25 vss 2.92378e-17
C6736 n4572_27 vss 2.92378e-17
C6737 n4572_26 vss 2.92378e-17
C6738 n4572_28 vss 2.92378e-17
C6739 n4572_27 vss 2.92378e-17
C6740 n4572_29 vss 2.92378e-17
C6741 n4572_28 vss 2.92378e-17
C6742 n4572_30 vss 8.77133e-17
C6743 n4572_29 vss 8.77133e-17
C6744 n4572_31 vss 9.50227e-17
C6745 n4572_30 vss 9.50227e-17
C6746 n4572_32 vss 2.92378e-17
C6747 n4572_31 vss 2.92378e-17
C6748 n4572_33 vss 2.92378e-17
C6749 n4572_32 vss 2.92378e-17
C6750 n4572_34 vss 2.92378e-17
C6751 n4572_33 vss 2.92378e-17
C6752 n4572_35 vss 2.92378e-17
C6753 n4572_34 vss 2.92378e-17
C6754 n4572_36 vss 2.92378e-17
C6755 n4572_35 vss 2.92378e-17
C6756 n4572_37 vss 2.92378e-17
C6757 n4572_36 vss 2.92378e-17

R152_1 s_3_1 s_3_379 0.001
R152_2 s_3_1 s_3_380 0.001
R152_3 s_3_1 s_3_378 0.001
R152_4 s_3_1 s_3_377 0.001
R152_5 s_3_1 s_3_375 0.001
R152_6 s_3_1 s_3_376 0.001
R152_7 s_3_1 s_3_374 0.001
R152_8 s_3_1 s_3_372 0.001
R152_9 s_3_1 s_3_373 0.001
R152_10 s_3_1 s_3_371 0.001
R152_11 s_3_1 s_3_370 0.001
R152_12 s_3_1 s_3_369 0.001
R152_13 s_3_1 s_3_368 0.001
R152_14 s_3_1 s_3_367 0.001
R152_15 s_3_1 s_3_366 0.001
R152_16 s_3_1 s_3_365 0.001
R152_17 s_3_1 s_3_364 0.001
R152_18 s_3_1 s_3_363 0.001
R152_19 s_3_1 s_3_362 0.001
R152_20 s_3_1 s_3_361 0.001
R152_21 s_3_360 s_3_2 0.001
R152_22 s_3_359 s_3_2 0.001
R152_23 s_3_358 s_3_2 0.001
R152_24 s_3_357 s_3_2 0.001
R152_25 s_3_356 s_3_2 0.001
R152_26 s_3_355 s_3_2 0.001
R152_27 s_3_354 s_3_2 0.001
R152_28 s_3_353 s_3_2 0.001
R152_29 s_3_112 s_3_3 0.001
R152_30 s_3_111 s_3_3 0.001
R152_31 s_3_110 s_3_3 0.001
R152_32 s_3_109 s_3_3 0.001
R152_33 s_3_107 s_3_3 0.001
R152_34 s_3_108 s_3_3 0.001
R152_35 s_3_106 s_3_3 0.001
R152_36 s_3_104 s_3_3 0.001
R152_37 s_3_105 s_3_3 0.001
R152_38 s_3_103 s_3_3 0.001
R152_39 s_3_102 s_3_3 0.001
R152_40 s_3_101 s_3_3 0.001
R152_41 s_3_100 s_3_3 0.001
R152_42 s_3_99 s_3_3 0.001
R152_43 s_3_98 s_3_3 0.001
R152_44 s_3_97 s_3_3 0.001
R152_45 s_3_96 s_3_3 0.001
R152_46 s_3_95 s_3_3 0.001
R152_47 s_3_94 s_3_3 0.001
R152_48 s_3_93 s_3_3 0.001
R152_49 s_3_91 s_3_4 0.001
R152_50 s_3_92 s_3_4 0.001
R152_51 s_3_90 s_3_4 0.001
R152_52 s_3_89 s_3_4 0.001
R152_53 s_3_88 s_3_4 0.001
R152_54 s_3_87 s_3_4 0.001
R152_55 s_3_86 s_3_4 0.001
R152_56 s_3_85 s_3_4 0.001
R152_57 s_3_82 s_3_5 0.001
R152_58 s_3_83 s_3_5 0.001
R152_59 s_3_81 s_3_5 0.001
R152_60 s_3_80 s_3_5 0.001
R152_61 s_3_78 s_3_5 0.001
R152_62 s_3_79 s_3_5 0.001
R152_63 s_3_77 s_3_5 0.001
R152_64 s_3_75 s_3_5 0.001
R152_65 s_3_76 s_3_5 0.001
R152_66 s_3_74 s_3_5 0.001
R152_67 s_3_73 s_3_5 0.001
R152_68 s_3_72 s_3_5 0.001
R152_69 s_3_71 s_3_5 0.001
R152_70 s_3_70 s_3_5 0.001
R152_71 s_3_69 s_3_5 0.001
R152_72 s_3_68 s_3_5 0.001
R152_73 s_3_67 s_3_5 0.001
R152_74 s_3_66 s_3_5 0.001
R152_75 s_3_64 s_3_5 0.001
R152_76 s_3_65 s_3_5 0.001
R152_77 s_3_63 s_3_6 0.001
R152_78 s_3_62 s_3_6 0.001
R152_79 s_3_61 s_3_6 0.001
R152_80 s_3_60 s_3_6 0.001
R152_81 s_3_59 s_3_6 0.001
R152_82 s_3_58 s_3_6 0.001
R152_83 s_3_57 s_3_6 0.001
R152_84 s_3_56 s_3_6 0.001
R152_85 s_3_54 s_3_7 0.001
R152_86 s_3_53 s_3_7 0.001
R152_87 s_3_52 s_3_7 0.001
R152_88 s_3_51 s_3_7 0.001
R152_89 s_3_49 s_3_7 0.001
R152_90 s_3_50 s_3_7 0.001
R152_91 s_3_48 s_3_7 0.001
R152_92 s_3_46 s_3_7 0.001
R152_93 s_3_47 s_3_7 0.001
R152_94 s_3_45 s_3_7 0.001
R152_95 s_3_44 s_3_7 0.001
R152_96 s_3_43 s_3_7 0.001
R152_97 s_3_42 s_3_7 0.001
R152_98 s_3_41 s_3_7 0.001
R152_99 s_3_40 s_3_7 0.001
R152_100 s_3_39 s_3_7 0.001
R152_101 s_3_38 s_3_7 0.001
R152_102 s_3_37 s_3_7 0.001
R152_103 s_3_35 s_3_7 0.001
R152_104 s_3_36 s_3_7 0.001
R152_105 s_3_34 s_3_8 0.001
R152_106 s_3_33 s_3_8 0.001
R152_107 s_3_32 s_3_8 0.001
R152_108 s_3_31 s_3_8 0.001
R152_109 s_3_30 s_3_8 0.001
R152_110 s_3_29 s_3_8 0.001
R152_111 s_3_28 s_3_8 0.001
R152_112 s_3_27 s_3_8 0.001
R152_113 s_3_199 s_3_9 0.001
R152_114 s_3_198 s_3_9 0.001
R152_115 s_3_197 s_3_9 0.001
R152_116 s_3_196 s_3_9 0.001
R152_117 s_3_194 s_3_9 0.001
R152_118 s_3_195 s_3_9 0.001
R152_119 s_3_193 s_3_9 0.001
R152_120 s_3_191 s_3_9 0.001
R152_121 s_3_192 s_3_9 0.001
R152_122 s_3_190 s_3_9 0.001
R152_123 s_3_189 s_3_9 0.001
R152_124 s_3_188 s_3_9 0.001
R152_125 s_3_187 s_3_9 0.001
R152_126 s_3_186 s_3_9 0.001
R152_127 s_3_185 s_3_9 0.001
R152_128 s_3_184 s_3_9 0.001
R152_129 s_3_183 s_3_9 0.001
R152_130 s_3_182 s_3_9 0.001
R152_131 s_3_180 s_3_9 0.001
R152_132 s_3_181 s_3_9 0.001
R152_133 s_3_179 s_3_10 0.001
R152_134 s_3_178 s_3_10 0.001
R152_135 s_3_177 s_3_10 0.001
R152_136 s_3_176 s_3_10 0.001
R152_137 s_3_175 s_3_10 0.001
R152_138 s_3_174 s_3_10 0.001
R152_139 s_3_173 s_3_10 0.001
R152_140 s_3_172 s_3_10 0.001
R152_141 s_3_170 s_3_11 0.001
R152_142 s_3_169 s_3_11 0.001
R152_143 s_3_168 s_3_11 0.001
R152_144 s_3_167 s_3_11 0.001
R152_145 s_3_165 s_3_11 0.001
R152_146 s_3_166 s_3_11 0.001
R152_147 s_3_164 s_3_11 0.001
R152_148 s_3_162 s_3_11 0.001
R152_149 s_3_163 s_3_11 0.001
R152_150 s_3_161 s_3_11 0.001
R152_151 s_3_160 s_3_11 0.001
R152_152 s_3_159 s_3_11 0.001
R152_153 s_3_158 s_3_11 0.001
R152_154 s_3_157 s_3_11 0.001
R152_155 s_3_156 s_3_11 0.001
R152_156 s_3_155 s_3_11 0.001
R152_157 s_3_154 s_3_11 0.001
R152_158 s_3_153 s_3_11 0.001
R152_159 s_3_152 s_3_11 0.001
R152_160 s_3_151 s_3_11 0.001
R152_161 s_3_149 s_3_12 0.001
R152_162 s_3_150 s_3_12 0.001
R152_163 s_3_148 s_3_12 0.001
R152_164 s_3_147 s_3_12 0.001
R152_165 s_3_146 s_3_12 0.001
R152_166 s_3_145 s_3_12 0.001
R152_167 s_3_144 s_3_12 0.001
R152_168 s_3_143 s_3_12 0.001
R152_169 s_3_140 s_3_13 0.001
R152_170 s_3_141 s_3_13 0.001
R152_171 s_3_139 s_3_13 0.001
R152_172 s_3_138 s_3_13 0.001
R152_173 s_3_136 s_3_13 0.001
R152_174 s_3_137 s_3_13 0.001
R152_175 s_3_135 s_3_13 0.001
R152_176 s_3_133 s_3_13 0.001
R152_177 s_3_134 s_3_13 0.001
R152_178 s_3_132 s_3_13 0.001
R152_179 s_3_131 s_3_13 0.001
R152_180 s_3_130 s_3_13 0.001
R152_181 s_3_129 s_3_13 0.001
R152_182 s_3_128 s_3_13 0.001
R152_183 s_3_127 s_3_13 0.001
R152_184 s_3_126 s_3_13 0.001
R152_185 s_3_125 s_3_13 0.001
R152_186 s_3_124 s_3_13 0.001
R152_187 s_3_122 s_3_13 0.001
R152_188 s_3_123 s_3_13 0.001
R152_189 s_3_121 s_3_14 0.001
R152_190 s_3_120 s_3_14 0.001
R152_191 s_3_119 s_3_14 0.001
R152_192 s_3_118 s_3_14 0.001
R152_193 s_3_117 s_3_14 0.001
R152_194 s_3_116 s_3_14 0.001
R152_195 s_3_115 s_3_14 0.001
R152_196 s_3_114 s_3_14 0.001
R152_197 s_3_257 s_3_15 0.001
R152_198 s_3_256 s_3_15 0.001
R152_199 s_3_255 s_3_15 0.001
R152_200 s_3_254 s_3_15 0.001
R152_201 s_3_252 s_3_15 0.001
R152_202 s_3_253 s_3_15 0.001
R152_203 s_3_251 s_3_15 0.001
R152_204 s_3_249 s_3_15 0.001
R152_205 s_3_250 s_3_15 0.001
R152_206 s_3_248 s_3_15 0.001
R152_207 s_3_247 s_3_15 0.001
R152_208 s_3_246 s_3_15 0.001
R152_209 s_3_245 s_3_15 0.001
R152_210 s_3_244 s_3_15 0.001
R152_211 s_3_243 s_3_15 0.001
R152_212 s_3_242 s_3_15 0.001
R152_213 s_3_241 s_3_15 0.001
R152_214 s_3_240 s_3_15 0.001
R152_215 s_3_238 s_3_15 0.001
R152_216 s_3_239 s_3_15 0.001
R152_217 s_3_236 s_3_16 0.001
R152_218 s_3_237 s_3_16 0.001
R152_219 s_3_235 s_3_16 0.001
R152_220 s_3_234 s_3_16 0.001
R152_221 s_3_233 s_3_16 0.001
R152_222 s_3_232 s_3_16 0.001
R152_223 s_3_231 s_3_16 0.001
R152_224 s_3_230 s_3_16 0.001
R152_225 s_3_228 s_3_17 0.001
R152_226 s_3_227 s_3_17 0.001
R152_227 s_3_226 s_3_17 0.001
R152_228 s_3_225 s_3_17 0.001
R152_229 s_3_223 s_3_17 0.001
R152_230 s_3_224 s_3_17 0.001
R152_231 s_3_222 s_3_17 0.001
R152_232 s_3_221 s_3_17 0.001
R152_233 s_3_220 s_3_17 0.001
R152_234 s_3_219 s_3_17 0.001
R152_235 s_3_218 s_3_17 0.001
R152_236 s_3_217 s_3_17 0.001
R152_237 s_3_216 s_3_17 0.001
R152_238 s_3_215 s_3_17 0.001
R152_239 s_3_214 s_3_17 0.001
R152_240 s_3_213 s_3_17 0.001
R152_241 s_3_212 s_3_17 0.001
R152_242 s_3_211 s_3_17 0.001
R152_243 s_3_210 s_3_17 0.001
R152_244 s_3_209 s_3_17 0.001
R152_245 s_3_208 s_3_18 0.001
R152_246 s_3_207 s_3_18 0.001
R152_247 s_3_206 s_3_18 0.001
R152_248 s_3_205 s_3_18 0.001
R152_249 s_3_204 s_3_18 0.001
R152_250 s_3_203 s_3_18 0.001
R152_251 s_3_202 s_3_18 0.001
R152_252 s_3_201 s_3_18 0.001
R152_253 s_3_344 s_3_19 0.001
R152_254 s_3_343 s_3_19 0.001
R152_255 s_3_342 s_3_19 0.001
R152_256 s_3_341 s_3_19 0.001
R152_257 s_3_339 s_3_19 0.001
R152_258 s_3_340 s_3_19 0.001
R152_259 s_3_338 s_3_19 0.001
R152_260 s_3_336 s_3_19 0.001
R152_261 s_3_337 s_3_19 0.001
R152_262 s_3_335 s_3_19 0.001
R152_263 s_3_334 s_3_19 0.001
R152_264 s_3_333 s_3_19 0.001
R152_265 s_3_332 s_3_19 0.001
R152_266 s_3_331 s_3_19 0.001
R152_267 s_3_330 s_3_19 0.001
R152_268 s_3_329 s_3_19 0.001
R152_269 s_3_328 s_3_19 0.001
R152_270 s_3_327 s_3_19 0.001
R152_271 s_3_326 s_3_19 0.001
R152_272 s_3_325 s_3_19 0.001
R152_273 s_3_323 s_3_20 0.001
R152_274 s_3_324 s_3_20 0.001
R152_275 s_3_322 s_3_20 0.001
R152_276 s_3_321 s_3_20 0.001
R152_277 s_3_320 s_3_20 0.001
R152_278 s_3_319 s_3_20 0.001
R152_279 s_3_318 s_3_20 0.001
R152_280 s_3_317 s_3_20 0.001
R152_281 s_3_314 s_3_21 0.001
R152_282 s_3_315 s_3_21 0.001
R152_283 s_3_313 s_3_21 0.001
R152_284 s_3_312 s_3_21 0.001
R152_285 s_3_310 s_3_21 0.001
R152_286 s_3_311 s_3_21 0.001
R152_287 s_3_309 s_3_21 0.001
R152_288 s_3_307 s_3_21 0.001
R152_289 s_3_308 s_3_21 0.001
R152_290 s_3_306 s_3_21 0.001
R152_291 s_3_305 s_3_21 0.001
R152_292 s_3_304 s_3_21 0.001
R152_293 s_3_303 s_3_21 0.001
R152_294 s_3_302 s_3_21 0.001
R152_295 s_3_301 s_3_21 0.001
R152_296 s_3_300 s_3_21 0.001
R152_297 s_3_299 s_3_21 0.001
R152_298 s_3_298 s_3_21 0.001
R152_299 s_3_296 s_3_21 0.001
R152_300 s_3_297 s_3_21 0.001
R152_301 s_3_295 s_3_22 0.001
R152_302 s_3_294 s_3_22 0.001
R152_303 s_3_293 s_3_22 0.001
R152_304 s_3_292 s_3_22 0.001
R152_305 s_3_291 s_3_22 0.001
R152_306 s_3_290 s_3_22 0.001
R152_307 s_3_289 s_3_22 0.001
R152_308 s_3_288 s_3_22 0.001
R152_309 s_3 s_3_23 0.001
R152_310 s_3_286 s_3_24 0.001
R152_311 s_3_285 s_3_24 0.001
R152_312 s_3_284 s_3_24 0.001
R152_313 s_3_283 s_3_24 0.001
R152_314 s_3_281 s_3_24 0.001
R152_315 s_3_282 s_3_24 0.001
R152_316 s_3_280 s_3_24 0.001
R152_317 s_3_278 s_3_24 0.001
R152_318 s_3_279 s_3_24 0.001
R152_319 s_3_277 s_3_24 0.001
R152_320 s_3_276 s_3_24 0.001
R152_321 s_3_275 s_3_24 0.001
R152_322 s_3_274 s_3_24 0.001
R152_323 s_3_273 s_3_24 0.001
R152_324 s_3_272 s_3_24 0.001
R152_325 s_3_271 s_3_24 0.001
R152_326 s_3_270 s_3_24 0.001
R152_327 s_3_269 s_3_24 0.001
R152_328 s_3_267 s_3_24 0.001
R152_329 s_3_268 s_3_24 0.001
R152_330 s_3_266 s_3_25 0.001
R152_331 s_3_265 s_3_25 0.001
R152_332 s_3_264 s_3_25 0.001
R152_333 s_3_263 s_3_25 0.001
R152_334 s_3_262 s_3_25 0.001
R152_335 s_3_261 s_3_25 0.001
R152_336 s_3_260 s_3_25 0.001
R152_337 s_3_259 s_3_25 0.001
R152_338 s_3_349 s_3 0.108
R152_339 s_3_27 s_3_349 1.296
R152_340 s_3_28 s_3_27 0.108
R152_341 s_3_29 s_3_28 0.108
R152_342 s_3_30 s_3_29 0.108
R152_343 s_3_31 s_3_30 0.108
R152_344 s_3_32 s_3_31 0.108
R152_345 s_3_33 s_3_32 0.108
R152_346 s_3_34 s_3_33 0.108
R152_347 s_3_35 s_3_34 0.864
R152_348 s_3_36 s_3_35 0.108
R152_349 s_3_37 s_3_36 0.108
R152_350 s_3_38 s_3_37 0.108
R152_351 s_3_39 s_3_38 0.108
R152_352 s_3_40 s_3_39 0.108
R152_353 s_3_41 s_3_40 0.108
R152_354 s_3_42 s_3_41 0.108
R152_355 s_3_43 s_3_42 0.108
R152_356 s_3_44 s_3_43 0.108
R152_357 s_3_45 s_3_44 0.108
R152_358 s_3_46 s_3_45 0.108
R152_359 s_3_47 s_3_46 0.108
R152_360 s_3_48 s_3_47 0.108
R152_361 s_3_49 s_3_48 0.108
R152_362 s_3_50 s_3_49 0.108
R152_363 s_3_51 s_3_50 0.108
R152_364 s_3_52 s_3_51 0.108
R152_365 s_3_53 s_3_52 0.108
R152_366 s_3_54 s_3_53 0.108
R152_367 s_3_55 s_3_54 0.001
R152_368 s_3_56 s_3_349 1.296
R152_369 s_3_57 s_3_56 0.108
R152_370 s_3_58 s_3_57 0.108
R152_371 s_3_59 s_3_58 0.108
R152_372 s_3_60 s_3_59 0.108
R152_373 s_3_61 s_3_60 0.108
R152_374 s_3_62 s_3_61 0.108
R152_375 s_3_63 s_3_62 0.108
R152_376 s_3_64 s_3_63 0.864
R152_377 s_3_65 s_3_64 0.108
R152_378 s_3_66 s_3_65 0.108
R152_379 s_3_67 s_3_66 0.108
R152_380 s_3_68 s_3_67 0.108
R152_381 s_3_69 s_3_68 0.108
R152_382 s_3_70 s_3_69 0.108
R152_383 s_3_71 s_3_70 0.108
R152_384 s_3_72 s_3_71 0.108
R152_385 s_3_73 s_3_72 0.108
R152_386 s_3_74 s_3_73 0.108
R152_387 s_3_75 s_3_74 0.108
R152_388 s_3_76 s_3_75 0.108
R152_389 s_3_77 s_3_76 0.108
R152_390 s_3_78 s_3_77 0.108
R152_391 s_3_79 s_3_78 0.108
R152_392 s_3_80 s_3_79 0.108
R152_393 s_3_81 s_3_80 0.108
R152_394 s_3_82 s_3_81 0.108
R152_395 s_3_83 s_3_82 0.108
R152_396 s_3_84 s_3_83 0.001
R152_397 s_3_85 s_3_350 0.54
R152_398 s_3_86 s_3_85 0.108
R152_399 s_3_87 s_3_86 0.108
R152_400 s_3_88 s_3_87 0.108
R152_401 s_3_89 s_3_88 0.108
R152_402 s_3_90 s_3_89 0.108
R152_403 s_3_91 s_3_90 0.108
R152_404 s_3_92 s_3_91 0.108
R152_405 s_3_93 s_3_92 0.864
R152_406 s_3_94 s_3_93 0.108
R152_407 s_3_95 s_3_94 0.108
R152_408 s_3_96 s_3_95 0.108
R152_409 s_3_97 s_3_96 0.108
R152_410 s_3_98 s_3_97 0.108
R152_411 s_3_99 s_3_98 0.108
R152_412 s_3_100 s_3_99 0.108
R152_413 s_3_101 s_3_100 0.108
R152_414 s_3_102 s_3_101 0.108
R152_415 s_3_103 s_3_102 0.108
R152_416 s_3_104 s_3_103 0.108
R152_417 s_3_105 s_3_104 0.108
R152_418 s_3_106 s_3_105 0.108
R152_419 s_3_107 s_3_106 0.108
R152_420 s_3_108 s_3_107 0.108
R152_421 s_3_109 s_3_108 0.108
R152_422 s_3_110 s_3_109 0.108
R152_423 s_3_111 s_3_110 0.108
R152_424 s_3_112 s_3_111 0.108
R152_425 s_3_113 s_3_112 0.001
R152_426 s_3_114 s_3_349 1.296
R152_427 s_3_115 s_3_114 0.108
R152_428 s_3_116 s_3_115 0.108
R152_429 s_3_117 s_3_116 0.108
R152_430 s_3_118 s_3_117 0.108
R152_431 s_3_119 s_3_118 0.108
R152_432 s_3_120 s_3_119 0.108
R152_433 s_3_121 s_3_120 0.108
R152_434 s_3_122 s_3_121 0.864
R152_435 s_3_123 s_3_122 0.108
R152_436 s_3_124 s_3_123 0.108
R152_437 s_3_125 s_3_124 0.108
R152_438 s_3_126 s_3_125 0.108
R152_439 s_3_127 s_3_126 0.108
R152_440 s_3_128 s_3_127 0.108
R152_441 s_3_129 s_3_128 0.108
R152_442 s_3_130 s_3_129 0.108
R152_443 s_3_131 s_3_130 0.108
R152_444 s_3_132 s_3_131 0.108
R152_445 s_3_133 s_3_132 0.108
R152_446 s_3_134 s_3_133 0.108
R152_447 s_3_135 s_3_134 0.108
R152_448 s_3_136 s_3_135 0.108
R152_449 s_3_137 s_3_136 0.108
R152_450 s_3_138 s_3_137 0.108
R152_451 s_3_139 s_3_138 0.108
R152_452 s_3_140 s_3_139 0.108
R152_453 s_3_141 s_3_140 0.108
R152_454 s_3_142 s_3_141 0.001
R152_455 s_3_143 s_3_349 1.296
R152_456 s_3_144 s_3_143 0.108
R152_457 s_3_145 s_3_144 0.108
R152_458 s_3_146 s_3_145 0.108
R152_459 s_3_147 s_3_146 0.108
R152_460 s_3_148 s_3_147 0.108
R152_461 s_3_149 s_3_148 0.108
R152_462 s_3_150 s_3_149 0.108
R152_463 s_3_151 s_3_150 0.864
R152_464 s_3_152 s_3_151 0.108
R152_465 s_3_153 s_3_152 0.108
R152_466 s_3_154 s_3_153 0.108
R152_467 s_3_155 s_3_154 0.108
R152_468 s_3_156 s_3_155 0.108
R152_469 s_3_157 s_3_156 0.108
R152_470 s_3_158 s_3_157 0.108
R152_471 s_3_159 s_3_158 0.108
R152_472 s_3_160 s_3_159 0.108
R152_473 s_3_161 s_3_160 0.108
R152_474 s_3_162 s_3_161 0.108
R152_475 s_3_163 s_3_162 0.108
R152_476 s_3_164 s_3_163 0.108
R152_477 s_3_165 s_3_164 0.108
R152_478 s_3_166 s_3_165 0.108
R152_479 s_3_167 s_3_166 0.108
R152_480 s_3_168 s_3_167 0.108
R152_481 s_3_169 s_3_168 0.108
R152_482 s_3_170 s_3_169 0.108
R152_483 s_3_171 s_3_170 0.001
R152_484 s_3_172 s_3_349 1.296
R152_485 s_3_173 s_3_172 0.108
R152_486 s_3_174 s_3_173 0.108
R152_487 s_3_175 s_3_174 0.108
R152_488 s_3_176 s_3_175 0.108
R152_489 s_3_177 s_3_176 0.108
R152_490 s_3_178 s_3_177 0.108
R152_491 s_3_179 s_3_178 0.108
R152_492 s_3_180 s_3_179 0.864
R152_493 s_3_181 s_3_180 0.108
R152_494 s_3_182 s_3_181 0.108
R152_495 s_3_183 s_3_182 0.108
R152_496 s_3_184 s_3_183 0.108
R152_497 s_3_185 s_3_184 0.108
R152_498 s_3_186 s_3_185 0.108
R152_499 s_3_187 s_3_186 0.108
R152_500 s_3_188 s_3_187 0.108
R152_501 s_3_189 s_3_188 0.108
R152_502 s_3_190 s_3_189 0.108
R152_503 s_3_191 s_3_190 0.108
R152_504 s_3_192 s_3_191 0.108
R152_505 s_3_193 s_3_192 0.108
R152_506 s_3_194 s_3_193 0.108
R152_507 s_3_195 s_3_194 0.108
R152_508 s_3_196 s_3_195 0.108
R152_509 s_3_197 s_3_196 0.108
R152_510 s_3_198 s_3_197 0.108
R152_511 s_3_199 s_3_198 0.108
R152_512 s_3_200 s_3_199 0.001
R152_513 s_3_201 s_3_349 1.296
R152_514 s_3_202 s_3_201 0.108
R152_515 s_3_203 s_3_202 0.108
R152_516 s_3_204 s_3_203 0.108
R152_517 s_3_205 s_3_204 0.108
R152_518 s_3_206 s_3_205 0.108
R152_519 s_3_207 s_3_206 0.108
R152_520 s_3_208 s_3_207 0.108
R152_521 s_3_209 s_3_208 0.864
R152_522 s_3_210 s_3_209 0.108
R152_523 s_3_211 s_3_210 0.108
R152_524 s_3_212 s_3_211 0.108
R152_525 s_3_213 s_3_212 0.108
R152_526 s_3_214 s_3_213 0.108
R152_527 s_3_215 s_3_214 0.108
R152_528 s_3_216 s_3_215 0.108
R152_529 s_3_217 s_3_216 0.108
R152_530 s_3_218 s_3_217 0.108
R152_531 s_3_219 s_3_218 0.108
R152_532 s_3_220 s_3_219 0.108
R152_533 s_3_221 s_3_220 0.108
R152_534 s_3_222 s_3_221 0.108
R152_535 s_3_223 s_3_222 0.108
R152_536 s_3_224 s_3_223 0.108
R152_537 s_3_225 s_3_224 0.108
R152_538 s_3_226 s_3_225 0.108
R152_539 s_3_227 s_3_226 0.108
R152_540 s_3_228 s_3_227 0.108
R152_541 s_3_229 s_3_228 0.001
R152_542 s_3_230 s_3_349 1.296
R152_543 s_3_231 s_3_230 0.108
R152_544 s_3_232 s_3_231 0.108
R152_545 s_3_233 s_3_232 0.108
R152_546 s_3_234 s_3_233 0.108
R152_547 s_3_235 s_3_234 0.108
R152_548 s_3_236 s_3_235 0.108
R152_549 s_3_237 s_3_236 0.108
R152_550 s_3_238 s_3_237 0.864
R152_551 s_3_239 s_3_238 0.108
R152_552 s_3_240 s_3_239 0.108
R152_553 s_3_241 s_3_240 0.108
R152_554 s_3_242 s_3_241 0.108
R152_555 s_3_243 s_3_242 0.108
R152_556 s_3_244 s_3_243 0.108
R152_557 s_3_245 s_3_244 0.108
R152_558 s_3_246 s_3_245 0.108
R152_559 s_3_247 s_3_246 0.108
R152_560 s_3_248 s_3_247 0.108
R152_561 s_3_249 s_3_248 0.108
R152_562 s_3_250 s_3_249 0.108
R152_563 s_3_251 s_3_250 0.108
R152_564 s_3_252 s_3_251 0.108
R152_565 s_3_253 s_3_252 0.108
R152_566 s_3_254 s_3_253 0.108
R152_567 s_3_255 s_3_254 0.108
R152_568 s_3_256 s_3_255 0.108
R152_569 s_3_257 s_3_256 0.108
R152_570 s_3_258 s_3_257 0.001
R152_571 s_3_259 s_3_346 0.54
R152_572 s_3_260 s_3_259 0.108
R152_573 s_3_261 s_3_260 0.108
R152_574 s_3_262 s_3_261 0.108
R152_575 s_3_263 s_3_262 0.108
R152_576 s_3_264 s_3_263 0.108
R152_577 s_3_265 s_3_264 0.108
R152_578 s_3_266 s_3_265 0.108
R152_579 s_3_267 s_3_266 0.864
R152_580 s_3_268 s_3_267 0.108
R152_581 s_3_269 s_3_268 0.108
R152_582 s_3_270 s_3_269 0.108
R152_583 s_3_271 s_3_270 0.108
R152_584 s_3_272 s_3_271 0.108
R152_585 s_3_273 s_3_272 0.108
R152_586 s_3_274 s_3_273 0.108
R152_587 s_3_275 s_3_274 0.108
R152_588 s_3_276 s_3_275 0.108
R152_589 s_3_277 s_3_276 0.108
R152_590 s_3_278 s_3_277 0.108
R152_591 s_3_279 s_3_278 0.108
R152_592 s_3_280 s_3_279 0.108
R152_593 s_3_281 s_3_280 0.108
R152_594 s_3_282 s_3_281 0.108
R152_595 s_3_283 s_3_282 0.108
R152_596 s_3_284 s_3_283 0.108
R152_597 s_3_285 s_3_284 0.108
R152_598 s_3_286 s_3_285 0.108
R152_599 s_3_287 s_3_286 0.001
R152_600 s_3_288 s_3_348 0.54
R152_601 s_3_289 s_3_288 0.108
R152_602 s_3_290 s_3_289 0.108
R152_603 s_3_291 s_3_290 0.108
R152_604 s_3_292 s_3_291 0.108
R152_605 s_3_293 s_3_292 0.108
R152_606 s_3_294 s_3_293 0.108
R152_607 s_3_295 s_3_294 0.108
R152_608 s_3_296 s_3_295 0.864
R152_609 s_3_297 s_3_296 0.108
R152_610 s_3_298 s_3_297 0.108
R152_611 s_3_299 s_3_298 0.108
R152_612 s_3_300 s_3_299 0.108
R152_613 s_3_301 s_3_300 0.108
R152_614 s_3_302 s_3_301 0.108
R152_615 s_3_303 s_3_302 0.108
R152_616 s_3_304 s_3_303 0.108
R152_617 s_3_305 s_3_304 0.108
R152_618 s_3_306 s_3_305 0.108
R152_619 s_3_307 s_3_306 0.108
R152_620 s_3_308 s_3_307 0.108
R152_621 s_3_309 s_3_308 0.108
R152_622 s_3_310 s_3_309 0.108
R152_623 s_3_311 s_3_310 0.108
R152_624 s_3_312 s_3_311 0.108
R152_625 s_3_313 s_3_312 0.108
R152_626 s_3_314 s_3_313 0.108
R152_627 s_3_315 s_3_314 0.108
R152_628 s_3_316 s_3_315 0.001
R152_629 s_3_317 s_3_349 1.296
R152_630 s_3_318 s_3_317 0.108
R152_631 s_3_319 s_3_318 0.108
R152_632 s_3_320 s_3_319 0.108
R152_633 s_3_321 s_3_320 0.108
R152_634 s_3_322 s_3_321 0.108
R152_635 s_3_323 s_3_322 0.108
R152_636 s_3_324 s_3_323 0.108
R152_637 s_3_325 s_3_324 0.864
R152_638 s_3_326 s_3_325 0.108
R152_639 s_3_327 s_3_326 0.108
R152_640 s_3_328 s_3_327 0.108
R152_641 s_3_329 s_3_328 0.108
R152_642 s_3_330 s_3_329 0.108
R152_643 s_3_331 s_3_330 0.108
R152_644 s_3_332 s_3_331 0.108
R152_645 s_3_333 s_3_332 0.108
R152_646 s_3_334 s_3_333 0.108
R152_647 s_3_335 s_3_334 0.108
R152_648 s_3_336 s_3_335 0.108
R152_649 s_3_337 s_3_336 0.108
R152_650 s_3_338 s_3_337 0.108
R152_651 s_3_339 s_3_338 0.108
R152_652 s_3_340 s_3_339 0.108
R152_653 s_3_341 s_3_340 0.108
R152_654 s_3_342 s_3_341 0.108
R152_655 s_3_343 s_3_342 0.108
R152_656 s_3_344 s_3_343 0.108
R152_657 s_3_345 s_3_344 0.001
R152_658 s_3_347 s_3_346 0.001
R152_659 s_3_348 s_3_347 0.001
R152_660 s_3_349 s_3_348 0.001
R152_661 s_3_350 s_3_349 0.001
R152_662 s_3_351 s_3_350 0.001
R152_663 s_3_352 s_3_351 0.001
R152_664 s_3_353 s_3_352 0.54
R152_665 s_3_354 s_3_353 0.108
R152_666 s_3_355 s_3_354 0.108
R152_667 s_3_356 s_3_355 0.108
R152_668 s_3_357 s_3_356 0.108
R152_669 s_3_358 s_3_357 0.108
R152_670 s_3_359 s_3_358 0.108
R152_671 s_3_360 s_3_359 0.108
R152_672 s_3_361 s_3_360 0.864
R152_673 s_3_362 s_3_361 0.108
R152_674 s_3_363 s_3_362 0.108
R152_675 s_3_364 s_3_363 0.108
R152_676 s_3_365 s_3_364 0.108
R152_677 s_3_366 s_3_365 0.108
R152_678 s_3_367 s_3_366 0.108
R152_679 s_3_368 s_3_367 0.108
R152_680 s_3_369 s_3_368 0.108
R152_681 s_3_370 s_3_369 0.108
R152_682 s_3_371 s_3_370 0.108
R152_683 s_3_372 s_3_371 0.108
R152_684 s_3_373 s_3_372 0.108
R152_685 s_3_374 s_3_373 0.108
R152_686 s_3_375 s_3_374 0.108
R152_687 s_3_376 s_3_375 0.108
R152_688 s_3_377 s_3_376 0.108
R152_689 s_3_378 s_3_377 0.108
R152_690 s_3_379 s_3_378 0.108
R152_691 s_3_380 s_3_379 0.108
R152_692 s_3_381 s_3_380 0.001

C6758 s_3_349 vss 6.29069e-15
C6759 s_3 vss 6.29069e-15
C6760 s_3_27 vss 3.60081e-16
C6761 s_3_349 vss 3.60081e-16
C6762 s_3_28 vss 3.13114e-17
C6763 s_3_27 vss 3.13114e-17
C6764 s_3_29 vss 3.13114e-17
C6765 s_3_28 vss 3.13114e-17
C6766 s_3_30 vss 3.13114e-17
C6767 s_3_29 vss 3.13114e-17
C6768 s_3_31 vss 3.13114e-17
C6769 s_3_30 vss 3.13114e-17
C6770 s_3_32 vss 3.13114e-17
C6771 s_3_31 vss 3.13114e-17
C6772 s_3_33 vss 3.13114e-17
C6773 s_3_32 vss 3.13114e-17
C6774 s_3_34 vss 3.13114e-17
C6775 s_3_33 vss 3.13114e-17
C6776 s_3_35 vss 2.42663e-16
C6777 s_3_34 vss 2.42663e-16
C6778 s_3_36 vss 3.13114e-17
C6779 s_3_35 vss 3.13114e-17
C6780 s_3_37 vss 3.13114e-17
C6781 s_3_36 vss 3.13114e-17
C6782 s_3_38 vss 3.13114e-17
C6783 s_3_37 vss 3.13114e-17
C6784 s_3_39 vss 3.13114e-17
C6785 s_3_38 vss 3.13114e-17
C6786 s_3_40 vss 3.13114e-17
C6787 s_3_39 vss 3.13114e-17
C6788 s_3_41 vss 3.13114e-17
C6789 s_3_40 vss 3.13114e-17
C6790 s_3_42 vss 3.13114e-17
C6791 s_3_41 vss 3.13114e-17
C6792 s_3_43 vss 3.13114e-17
C6793 s_3_42 vss 3.13114e-17
C6794 s_3_44 vss 3.13114e-17
C6795 s_3_43 vss 3.13114e-17
C6796 s_3_45 vss 3.13114e-17
C6797 s_3_44 vss 3.13114e-17
C6798 s_3_46 vss 3.13114e-17
C6799 s_3_45 vss 3.13114e-17
C6800 s_3_47 vss 3.13114e-17
C6801 s_3_46 vss 3.13114e-17
C6802 s_3_48 vss 3.13114e-17
C6803 s_3_47 vss 3.13114e-17
C6804 s_3_49 vss 3.13114e-17
C6805 s_3_48 vss 3.13114e-17
C6806 s_3_50 vss 3.13114e-17
C6807 s_3_49 vss 3.13114e-17
C6808 s_3_51 vss 3.13114e-17
C6809 s_3_50 vss 3.13114e-17
C6810 s_3_52 vss 3.13114e-17
C6811 s_3_51 vss 3.13114e-17
C6812 s_3_53 vss 3.13114e-17
C6813 s_3_52 vss 3.13114e-17
C6814 s_3_54 vss 3.13114e-17
C6815 s_3_53 vss 3.13114e-17
C6816 s_3_55 vss 1.40901e-17
C6817 s_3_54 vss 1.40901e-17
C6818 s_3_56 vss 3.60081e-16
C6819 s_3_349 vss 3.60081e-16
C6820 s_3_57 vss 3.13114e-17
C6821 s_3_56 vss 3.13114e-17
C6822 s_3_58 vss 3.13114e-17
C6823 s_3_57 vss 3.13114e-17
C6824 s_3_59 vss 3.13114e-17
C6825 s_3_58 vss 3.13114e-17
C6826 s_3_60 vss 3.13114e-17
C6827 s_3_59 vss 3.13114e-17
C6828 s_3_61 vss 3.13114e-17
C6829 s_3_60 vss 3.13114e-17
C6830 s_3_62 vss 3.13114e-17
C6831 s_3_61 vss 3.13114e-17
C6832 s_3_63 vss 3.13114e-17
C6833 s_3_62 vss 3.13114e-17
C6834 s_3_64 vss 2.42663e-16
C6835 s_3_63 vss 2.42663e-16
C6836 s_3_65 vss 3.13114e-17
C6837 s_3_64 vss 3.13114e-17
C6838 s_3_66 vss 3.13114e-17
C6839 s_3_65 vss 3.13114e-17
C6840 s_3_67 vss 3.13114e-17
C6841 s_3_66 vss 3.13114e-17
C6842 s_3_68 vss 3.13114e-17
C6843 s_3_67 vss 3.13114e-17
C6844 s_3_69 vss 3.13114e-17
C6845 s_3_68 vss 3.13114e-17
C6846 s_3_70 vss 3.13114e-17
C6847 s_3_69 vss 3.13114e-17
C6848 s_3_71 vss 3.13114e-17
C6849 s_3_70 vss 3.13114e-17
C6850 s_3_72 vss 3.13114e-17
C6851 s_3_71 vss 3.13114e-17
C6852 s_3_73 vss 3.13114e-17
C6853 s_3_72 vss 3.13114e-17
C6854 s_3_74 vss 3.13114e-17
C6855 s_3_73 vss 3.13114e-17
C6856 s_3_75 vss 3.13114e-17
C6857 s_3_74 vss 3.13114e-17
C6858 s_3_76 vss 3.13114e-17
C6859 s_3_75 vss 3.13114e-17
C6860 s_3_77 vss 3.13114e-17
C6861 s_3_76 vss 3.13114e-17
C6862 s_3_78 vss 3.13114e-17
C6863 s_3_77 vss 3.13114e-17
C6864 s_3_79 vss 3.13114e-17
C6865 s_3_78 vss 3.13114e-17
C6866 s_3_80 vss 3.13114e-17
C6867 s_3_79 vss 3.13114e-17
C6868 s_3_81 vss 3.13114e-17
C6869 s_3_80 vss 3.13114e-17
C6870 s_3_82 vss 3.13114e-17
C6871 s_3_81 vss 3.13114e-17
C6872 s_3_83 vss 3.13114e-17
C6873 s_3_82 vss 3.13114e-17
C6874 s_3_84 vss 1.40901e-17
C6875 s_3_83 vss 1.40901e-17
C6876 s_3_85 vss 1.40901e-16
C6877 s_3_350 vss 1.40901e-16
C6878 s_3_86 vss 3.13114e-17
C6879 s_3_85 vss 3.13114e-17
C6880 s_3_87 vss 3.13114e-17
C6881 s_3_86 vss 3.13114e-17
C6882 s_3_88 vss 3.13114e-17
C6883 s_3_87 vss 3.13114e-17
C6884 s_3_89 vss 3.13114e-17
C6885 s_3_88 vss 3.13114e-17
C6886 s_3_90 vss 3.13114e-17
C6887 s_3_89 vss 3.13114e-17
C6888 s_3_91 vss 3.13114e-17
C6889 s_3_90 vss 3.13114e-17
C6890 s_3_92 vss 3.13114e-17
C6891 s_3_91 vss 3.13114e-17
C6892 s_3_93 vss 2.42663e-16
C6893 s_3_92 vss 2.42663e-16
C6894 s_3_94 vss 3.13114e-17
C6895 s_3_93 vss 3.13114e-17
C6896 s_3_95 vss 3.13114e-17
C6897 s_3_94 vss 3.13114e-17
C6898 s_3_96 vss 3.13114e-17
C6899 s_3_95 vss 3.13114e-17
C6900 s_3_97 vss 3.13114e-17
C6901 s_3_96 vss 3.13114e-17
C6902 s_3_98 vss 3.13114e-17
C6903 s_3_97 vss 3.13114e-17
C6904 s_3_99 vss 3.13114e-17
C6905 s_3_98 vss 3.13114e-17
C6906 s_3_100 vss 3.13114e-17
C6907 s_3_99 vss 3.13114e-17
C6908 s_3_101 vss 3.13114e-17
C6909 s_3_100 vss 3.13114e-17
C6910 s_3_102 vss 3.13114e-17
C6911 s_3_101 vss 3.13114e-17
C6912 s_3_103 vss 3.13114e-17
C6913 s_3_102 vss 3.13114e-17
C6914 s_3_104 vss 3.13114e-17
C6915 s_3_103 vss 3.13114e-17
C6916 s_3_105 vss 3.13114e-17
C6917 s_3_104 vss 3.13114e-17
C6918 s_3_106 vss 3.13114e-17
C6919 s_3_105 vss 3.13114e-17
C6920 s_3_107 vss 3.13114e-17
C6921 s_3_106 vss 3.13114e-17
C6922 s_3_108 vss 3.13114e-17
C6923 s_3_107 vss 3.13114e-17
C6924 s_3_109 vss 3.13114e-17
C6925 s_3_108 vss 3.13114e-17
C6926 s_3_110 vss 3.13114e-17
C6927 s_3_109 vss 3.13114e-17
C6928 s_3_111 vss 3.13114e-17
C6929 s_3_110 vss 3.13114e-17
C6930 s_3_112 vss 3.13114e-17
C6931 s_3_111 vss 3.13114e-17
C6932 s_3_113 vss 1.40901e-17
C6933 s_3_112 vss 1.40901e-17
C6934 s_3_114 vss 3.60081e-16
C6935 s_3_349 vss 3.60081e-16
C6936 s_3_115 vss 3.13114e-17
C6937 s_3_114 vss 3.13114e-17
C6938 s_3_116 vss 3.13114e-17
C6939 s_3_115 vss 3.13114e-17
C6940 s_3_117 vss 3.13114e-17
C6941 s_3_116 vss 3.13114e-17
C6942 s_3_118 vss 3.13114e-17
C6943 s_3_117 vss 3.13114e-17
C6944 s_3_119 vss 3.13114e-17
C6945 s_3_118 vss 3.13114e-17
C6946 s_3_120 vss 3.13114e-17
C6947 s_3_119 vss 3.13114e-17
C6948 s_3_121 vss 3.13114e-17
C6949 s_3_120 vss 3.13114e-17
C6950 s_3_122 vss 2.42663e-16
C6951 s_3_121 vss 2.42663e-16
C6952 s_3_123 vss 3.13114e-17
C6953 s_3_122 vss 3.13114e-17
C6954 s_3_124 vss 3.13114e-17
C6955 s_3_123 vss 3.13114e-17
C6956 s_3_125 vss 3.13114e-17
C6957 s_3_124 vss 3.13114e-17
C6958 s_3_126 vss 3.13114e-17
C6959 s_3_125 vss 3.13114e-17
C6960 s_3_127 vss 3.13114e-17
C6961 s_3_126 vss 3.13114e-17
C6962 s_3_128 vss 3.13114e-17
C6963 s_3_127 vss 3.13114e-17
C6964 s_3_129 vss 3.13114e-17
C6965 s_3_128 vss 3.13114e-17
C6966 s_3_130 vss 3.13114e-17
C6967 s_3_129 vss 3.13114e-17
C6968 s_3_131 vss 3.13114e-17
C6969 s_3_130 vss 3.13114e-17
C6970 s_3_132 vss 3.13114e-17
C6971 s_3_131 vss 3.13114e-17
C6972 s_3_133 vss 3.13114e-17
C6973 s_3_132 vss 3.13114e-17
C6974 s_3_134 vss 3.13114e-17
C6975 s_3_133 vss 3.13114e-17
C6976 s_3_135 vss 3.13114e-17
C6977 s_3_134 vss 3.13114e-17
C6978 s_3_136 vss 3.13114e-17
C6979 s_3_135 vss 3.13114e-17
C6980 s_3_137 vss 3.13114e-17
C6981 s_3_136 vss 3.13114e-17
C6982 s_3_138 vss 3.13114e-17
C6983 s_3_137 vss 3.13114e-17
C6984 s_3_139 vss 3.13114e-17
C6985 s_3_138 vss 3.13114e-17
C6986 s_3_140 vss 3.13114e-17
C6987 s_3_139 vss 3.13114e-17
C6988 s_3_141 vss 3.13114e-17
C6989 s_3_140 vss 3.13114e-17
C6990 s_3_142 vss 1.40901e-17
C6991 s_3_141 vss 1.40901e-17
C6992 s_3_143 vss 3.60081e-16
C6993 s_3_349 vss 3.60081e-16
C6994 s_3_144 vss 3.13114e-17
C6995 s_3_143 vss 3.13114e-17
C6996 s_3_145 vss 3.13114e-17
C6997 s_3_144 vss 3.13114e-17
C6998 s_3_146 vss 3.13114e-17
C6999 s_3_145 vss 3.13114e-17
C7000 s_3_147 vss 3.13114e-17
C7001 s_3_146 vss 3.13114e-17
C7002 s_3_148 vss 3.13114e-17
C7003 s_3_147 vss 3.13114e-17
C7004 s_3_149 vss 3.13114e-17
C7005 s_3_148 vss 3.13114e-17
C7006 s_3_150 vss 3.13114e-17
C7007 s_3_149 vss 3.13114e-17
C7008 s_3_151 vss 2.42663e-16
C7009 s_3_150 vss 2.42663e-16
C7010 s_3_152 vss 3.13114e-17
C7011 s_3_151 vss 3.13114e-17
C7012 s_3_153 vss 3.13114e-17
C7013 s_3_152 vss 3.13114e-17
C7014 s_3_154 vss 3.13114e-17
C7015 s_3_153 vss 3.13114e-17
C7016 s_3_155 vss 3.13114e-17
C7017 s_3_154 vss 3.13114e-17
C7018 s_3_156 vss 3.13114e-17
C7019 s_3_155 vss 3.13114e-17
C7020 s_3_157 vss 3.13114e-17
C7021 s_3_156 vss 3.13114e-17
C7022 s_3_158 vss 3.13114e-17
C7023 s_3_157 vss 3.13114e-17
C7024 s_3_159 vss 3.13114e-17
C7025 s_3_158 vss 3.13114e-17
C7026 s_3_160 vss 3.13114e-17
C7027 s_3_159 vss 3.13114e-17
C7028 s_3_161 vss 3.13114e-17
C7029 s_3_160 vss 3.13114e-17
C7030 s_3_162 vss 3.13114e-17
C7031 s_3_161 vss 3.13114e-17
C7032 s_3_163 vss 3.13114e-17
C7033 s_3_162 vss 3.13114e-17
C7034 s_3_164 vss 3.13114e-17
C7035 s_3_163 vss 3.13114e-17
C7036 s_3_165 vss 3.13114e-17
C7037 s_3_164 vss 3.13114e-17
C7038 s_3_166 vss 3.13114e-17
C7039 s_3_165 vss 3.13114e-17
C7040 s_3_167 vss 3.13114e-17
C7041 s_3_166 vss 3.13114e-17
C7042 s_3_168 vss 3.13114e-17
C7043 s_3_167 vss 3.13114e-17
C7044 s_3_169 vss 3.13114e-17
C7045 s_3_168 vss 3.13114e-17
C7046 s_3_170 vss 3.13114e-17
C7047 s_3_169 vss 3.13114e-17
C7048 s_3_171 vss 1.40901e-17
C7049 s_3_170 vss 1.40901e-17
C7050 s_3_172 vss 3.60081e-16
C7051 s_3_349 vss 3.60081e-16
C7052 s_3_173 vss 3.13114e-17
C7053 s_3_172 vss 3.13114e-17
C7054 s_3_174 vss 3.13114e-17
C7055 s_3_173 vss 3.13114e-17
C7056 s_3_175 vss 3.13114e-17
C7057 s_3_174 vss 3.13114e-17
C7058 s_3_176 vss 3.13114e-17
C7059 s_3_175 vss 3.13114e-17
C7060 s_3_177 vss 3.13114e-17
C7061 s_3_176 vss 3.13114e-17
C7062 s_3_178 vss 3.13114e-17
C7063 s_3_177 vss 3.13114e-17
C7064 s_3_179 vss 3.13114e-17
C7065 s_3_178 vss 3.13114e-17
C7066 s_3_180 vss 2.42663e-16
C7067 s_3_179 vss 2.42663e-16
C7068 s_3_181 vss 3.13114e-17
C7069 s_3_180 vss 3.13114e-17
C7070 s_3_182 vss 3.13114e-17
C7071 s_3_181 vss 3.13114e-17
C7072 s_3_183 vss 3.13114e-17
C7073 s_3_182 vss 3.13114e-17
C7074 s_3_184 vss 3.13114e-17
C7075 s_3_183 vss 3.13114e-17
C7076 s_3_185 vss 3.13114e-17
C7077 s_3_184 vss 3.13114e-17
C7078 s_3_186 vss 3.13114e-17
C7079 s_3_185 vss 3.13114e-17
C7080 s_3_187 vss 3.13114e-17
C7081 s_3_186 vss 3.13114e-17
C7082 s_3_188 vss 3.13114e-17
C7083 s_3_187 vss 3.13114e-17
C7084 s_3_189 vss 3.13114e-17
C7085 s_3_188 vss 3.13114e-17
C7086 s_3_190 vss 3.13114e-17
C7087 s_3_189 vss 3.13114e-17
C7088 s_3_191 vss 3.13114e-17
C7089 s_3_190 vss 3.13114e-17
C7090 s_3_192 vss 3.13114e-17
C7091 s_3_191 vss 3.13114e-17
C7092 s_3_193 vss 3.13114e-17
C7093 s_3_192 vss 3.13114e-17
C7094 s_3_194 vss 3.13114e-17
C7095 s_3_193 vss 3.13114e-17
C7096 s_3_195 vss 3.13114e-17
C7097 s_3_194 vss 3.13114e-17
C7098 s_3_196 vss 3.13114e-17
C7099 s_3_195 vss 3.13114e-17
C7100 s_3_197 vss 3.13114e-17
C7101 s_3_196 vss 3.13114e-17
C7102 s_3_198 vss 3.13114e-17
C7103 s_3_197 vss 3.13114e-17
C7104 s_3_199 vss 3.13114e-17
C7105 s_3_198 vss 3.13114e-17
C7106 s_3_200 vss 1.40901e-17
C7107 s_3_199 vss 1.40901e-17
C7108 s_3_201 vss 3.60081e-16
C7109 s_3_349 vss 3.60081e-16
C7110 s_3_202 vss 3.13114e-17
C7111 s_3_201 vss 3.13114e-17
C7112 s_3_203 vss 3.13114e-17
C7113 s_3_202 vss 3.13114e-17
C7114 s_3_204 vss 3.13114e-17
C7115 s_3_203 vss 3.13114e-17
C7116 s_3_205 vss 3.13114e-17
C7117 s_3_204 vss 3.13114e-17
C7118 s_3_206 vss 3.13114e-17
C7119 s_3_205 vss 3.13114e-17
C7120 s_3_207 vss 3.13114e-17
C7121 s_3_206 vss 3.13114e-17
C7122 s_3_208 vss 3.13114e-17
C7123 s_3_207 vss 3.13114e-17
C7124 s_3_209 vss 2.42663e-16
C7125 s_3_208 vss 2.42663e-16
C7126 s_3_210 vss 3.13114e-17
C7127 s_3_209 vss 3.13114e-17
C7128 s_3_211 vss 3.13114e-17
C7129 s_3_210 vss 3.13114e-17
C7130 s_3_212 vss 3.13114e-17
C7131 s_3_211 vss 3.13114e-17
C7132 s_3_213 vss 3.13114e-17
C7133 s_3_212 vss 3.13114e-17
C7134 s_3_214 vss 3.13114e-17
C7135 s_3_213 vss 3.13114e-17
C7136 s_3_215 vss 3.13114e-17
C7137 s_3_214 vss 3.13114e-17
C7138 s_3_216 vss 3.13114e-17
C7139 s_3_215 vss 3.13114e-17
C7140 s_3_217 vss 3.13114e-17
C7141 s_3_216 vss 3.13114e-17
C7142 s_3_218 vss 3.13114e-17
C7143 s_3_217 vss 3.13114e-17
C7144 s_3_219 vss 3.13114e-17
C7145 s_3_218 vss 3.13114e-17
C7146 s_3_220 vss 3.13114e-17
C7147 s_3_219 vss 3.13114e-17
C7148 s_3_221 vss 3.13114e-17
C7149 s_3_220 vss 3.13114e-17
C7150 s_3_222 vss 3.13114e-17
C7151 s_3_221 vss 3.13114e-17
C7152 s_3_223 vss 3.13114e-17
C7153 s_3_222 vss 3.13114e-17
C7154 s_3_224 vss 3.13114e-17
C7155 s_3_223 vss 3.13114e-17
C7156 s_3_225 vss 3.13114e-17
C7157 s_3_224 vss 3.13114e-17
C7158 s_3_226 vss 3.13114e-17
C7159 s_3_225 vss 3.13114e-17
C7160 s_3_227 vss 3.13114e-17
C7161 s_3_226 vss 3.13114e-17
C7162 s_3_228 vss 3.13114e-17
C7163 s_3_227 vss 3.13114e-17
C7164 s_3_229 vss 1.40901e-17
C7165 s_3_228 vss 1.40901e-17
C7166 s_3_230 vss 3.60081e-16
C7167 s_3_349 vss 3.60081e-16
C7168 s_3_231 vss 3.13114e-17
C7169 s_3_230 vss 3.13114e-17
C7170 s_3_232 vss 3.13114e-17
C7171 s_3_231 vss 3.13114e-17
C7172 s_3_233 vss 3.13114e-17
C7173 s_3_232 vss 3.13114e-17
C7174 s_3_234 vss 3.13114e-17
C7175 s_3_233 vss 3.13114e-17
C7176 s_3_235 vss 3.13114e-17
C7177 s_3_234 vss 3.13114e-17
C7178 s_3_236 vss 3.13114e-17
C7179 s_3_235 vss 3.13114e-17
C7180 s_3_237 vss 3.13114e-17
C7181 s_3_236 vss 3.13114e-17
C7182 s_3_238 vss 2.42663e-16
C7183 s_3_237 vss 2.42663e-16
C7184 s_3_239 vss 3.13114e-17
C7185 s_3_238 vss 3.13114e-17
C7186 s_3_240 vss 3.13114e-17
C7187 s_3_239 vss 3.13114e-17
C7188 s_3_241 vss 3.13114e-17
C7189 s_3_240 vss 3.13114e-17
C7190 s_3_242 vss 3.13114e-17
C7191 s_3_241 vss 3.13114e-17
C7192 s_3_243 vss 3.13114e-17
C7193 s_3_242 vss 3.13114e-17
C7194 s_3_244 vss 3.13114e-17
C7195 s_3_243 vss 3.13114e-17
C7196 s_3_245 vss 3.13114e-17
C7197 s_3_244 vss 3.13114e-17
C7198 s_3_246 vss 3.13114e-17
C7199 s_3_245 vss 3.13114e-17
C7200 s_3_247 vss 3.13114e-17
C7201 s_3_246 vss 3.13114e-17
C7202 s_3_248 vss 3.13114e-17
C7203 s_3_247 vss 3.13114e-17
C7204 s_3_249 vss 3.13114e-17
C7205 s_3_248 vss 3.13114e-17
C7206 s_3_250 vss 3.13114e-17
C7207 s_3_249 vss 3.13114e-17
C7208 s_3_251 vss 3.13114e-17
C7209 s_3_250 vss 3.13114e-17
C7210 s_3_252 vss 3.13114e-17
C7211 s_3_251 vss 3.13114e-17
C7212 s_3_253 vss 3.13114e-17
C7213 s_3_252 vss 3.13114e-17
C7214 s_3_254 vss 3.13114e-17
C7215 s_3_253 vss 3.13114e-17
C7216 s_3_255 vss 3.13114e-17
C7217 s_3_254 vss 3.13114e-17
C7218 s_3_256 vss 3.13114e-17
C7219 s_3_255 vss 3.13114e-17
C7220 s_3_257 vss 3.13114e-17
C7221 s_3_256 vss 3.13114e-17
C7222 s_3_258 vss 1.40901e-17
C7223 s_3_257 vss 1.40901e-17
C7224 s_3_259 vss 1.40901e-16
C7225 s_3_346 vss 1.40901e-16
C7226 s_3_260 vss 3.13114e-17
C7227 s_3_259 vss 3.13114e-17
C7228 s_3_261 vss 3.13114e-17
C7229 s_3_260 vss 3.13114e-17
C7230 s_3_262 vss 3.13114e-17
C7231 s_3_261 vss 3.13114e-17
C7232 s_3_263 vss 3.13114e-17
C7233 s_3_262 vss 3.13114e-17
C7234 s_3_264 vss 3.13114e-17
C7235 s_3_263 vss 3.13114e-17
C7236 s_3_265 vss 3.13114e-17
C7237 s_3_264 vss 3.13114e-17
C7238 s_3_266 vss 3.13114e-17
C7239 s_3_265 vss 3.13114e-17
C7240 s_3_267 vss 2.42663e-16
C7241 s_3_266 vss 2.42663e-16
C7242 s_3_268 vss 3.13114e-17
C7243 s_3_267 vss 3.13114e-17
C7244 s_3_269 vss 3.13114e-17
C7245 s_3_268 vss 3.13114e-17
C7246 s_3_270 vss 3.13114e-17
C7247 s_3_269 vss 3.13114e-17
C7248 s_3_271 vss 3.13114e-17
C7249 s_3_270 vss 3.13114e-17
C7250 s_3_272 vss 3.13114e-17
C7251 s_3_271 vss 3.13114e-17
C7252 s_3_273 vss 3.13114e-17
C7253 s_3_272 vss 3.13114e-17
C7254 s_3_274 vss 3.13114e-17
C7255 s_3_273 vss 3.13114e-17
C7256 s_3_275 vss 3.13114e-17
C7257 s_3_274 vss 3.13114e-17
C7258 s_3_276 vss 3.13114e-17
C7259 s_3_275 vss 3.13114e-17
C7260 s_3_277 vss 3.13114e-17
C7261 s_3_276 vss 3.13114e-17
C7262 s_3_278 vss 3.13114e-17
C7263 s_3_277 vss 3.13114e-17
C7264 s_3_279 vss 3.13114e-17
C7265 s_3_278 vss 3.13114e-17
C7266 s_3_280 vss 3.13114e-17
C7267 s_3_279 vss 3.13114e-17
C7268 s_3_281 vss 3.13114e-17
C7269 s_3_280 vss 3.13114e-17
C7270 s_3_282 vss 3.13114e-17
C7271 s_3_281 vss 3.13114e-17
C7272 s_3_283 vss 3.13114e-17
C7273 s_3_282 vss 3.13114e-17
C7274 s_3_284 vss 3.13114e-17
C7275 s_3_283 vss 3.13114e-17
C7276 s_3_285 vss 3.13114e-17
C7277 s_3_284 vss 3.13114e-17
C7278 s_3_286 vss 3.13114e-17
C7279 s_3_285 vss 3.13114e-17
C7280 s_3_287 vss 1.40901e-17
C7281 s_3_286 vss 1.40901e-17
C7282 s_3_288 vss 1.40901e-16
C7283 s_3_348 vss 1.40901e-16
C7284 s_3_289 vss 3.13114e-17
C7285 s_3_288 vss 3.13114e-17
C7286 s_3_290 vss 3.13114e-17
C7287 s_3_289 vss 3.13114e-17
C7288 s_3_291 vss 3.13114e-17
C7289 s_3_290 vss 3.13114e-17
C7290 s_3_292 vss 3.13114e-17
C7291 s_3_291 vss 3.13114e-17
C7292 s_3_293 vss 3.13114e-17
C7293 s_3_292 vss 3.13114e-17
C7294 s_3_294 vss 3.13114e-17
C7295 s_3_293 vss 3.13114e-17
C7296 s_3_295 vss 3.13114e-17
C7297 s_3_294 vss 3.13114e-17
C7298 s_3_296 vss 2.42663e-16
C7299 s_3_295 vss 2.42663e-16
C7300 s_3_297 vss 3.13114e-17
C7301 s_3_296 vss 3.13114e-17
C7302 s_3_298 vss 3.13114e-17
C7303 s_3_297 vss 3.13114e-17
C7304 s_3_299 vss 3.13114e-17
C7305 s_3_298 vss 3.13114e-17
C7306 s_3_300 vss 3.13114e-17
C7307 s_3_299 vss 3.13114e-17
C7308 s_3_301 vss 3.13114e-17
C7309 s_3_300 vss 3.13114e-17
C7310 s_3_302 vss 3.13114e-17
C7311 s_3_301 vss 3.13114e-17
C7312 s_3_303 vss 3.13114e-17
C7313 s_3_302 vss 3.13114e-17
C7314 s_3_304 vss 3.13114e-17
C7315 s_3_303 vss 3.13114e-17
C7316 s_3_305 vss 3.13114e-17
C7317 s_3_304 vss 3.13114e-17
C7318 s_3_306 vss 3.13114e-17
C7319 s_3_305 vss 3.13114e-17
C7320 s_3_307 vss 3.13114e-17
C7321 s_3_306 vss 3.13114e-17
C7322 s_3_308 vss 3.13114e-17
C7323 s_3_307 vss 3.13114e-17
C7324 s_3_309 vss 3.13114e-17
C7325 s_3_308 vss 3.13114e-17
C7326 s_3_310 vss 3.13114e-17
C7327 s_3_309 vss 3.13114e-17
C7328 s_3_311 vss 3.13114e-17
C7329 s_3_310 vss 3.13114e-17
C7330 s_3_312 vss 3.13114e-17
C7331 s_3_311 vss 3.13114e-17
C7332 s_3_313 vss 3.13114e-17
C7333 s_3_312 vss 3.13114e-17
C7334 s_3_314 vss 3.13114e-17
C7335 s_3_313 vss 3.13114e-17
C7336 s_3_315 vss 3.13114e-17
C7337 s_3_314 vss 3.13114e-17
C7338 s_3_316 vss 1.40901e-17
C7339 s_3_315 vss 1.40901e-17
C7340 s_3_317 vss 3.60081e-16
C7341 s_3_349 vss 3.60081e-16
C7342 s_3_318 vss 3.13114e-17
C7343 s_3_317 vss 3.13114e-17
C7344 s_3_319 vss 3.13114e-17
C7345 s_3_318 vss 3.13114e-17
C7346 s_3_320 vss 3.13114e-17
C7347 s_3_319 vss 3.13114e-17
C7348 s_3_321 vss 3.13114e-17
C7349 s_3_320 vss 3.13114e-17
C7350 s_3_322 vss 3.13114e-17
C7351 s_3_321 vss 3.13114e-17
C7352 s_3_323 vss 3.13114e-17
C7353 s_3_322 vss 3.13114e-17
C7354 s_3_324 vss 3.13114e-17
C7355 s_3_323 vss 3.13114e-17
C7356 s_3_325 vss 2.42663e-16
C7357 s_3_324 vss 2.42663e-16
C7358 s_3_326 vss 3.13114e-17
C7359 s_3_325 vss 3.13114e-17
C7360 s_3_327 vss 3.13114e-17
C7361 s_3_326 vss 3.13114e-17
C7362 s_3_328 vss 3.13114e-17
C7363 s_3_327 vss 3.13114e-17
C7364 s_3_329 vss 3.13114e-17
C7365 s_3_328 vss 3.13114e-17
C7366 s_3_330 vss 3.13114e-17
C7367 s_3_329 vss 3.13114e-17
C7368 s_3_331 vss 3.13114e-17
C7369 s_3_330 vss 3.13114e-17
C7370 s_3_332 vss 3.13114e-17
C7371 s_3_331 vss 3.13114e-17
C7372 s_3_333 vss 3.13114e-17
C7373 s_3_332 vss 3.13114e-17
C7374 s_3_334 vss 3.13114e-17
C7375 s_3_333 vss 3.13114e-17
C7376 s_3_335 vss 3.13114e-17
C7377 s_3_334 vss 3.13114e-17
C7378 s_3_336 vss 3.13114e-17
C7379 s_3_335 vss 3.13114e-17
C7380 s_3_337 vss 3.13114e-17
C7381 s_3_336 vss 3.13114e-17
C7382 s_3_338 vss 3.13114e-17
C7383 s_3_337 vss 3.13114e-17
C7384 s_3_339 vss 3.13114e-17
C7385 s_3_338 vss 3.13114e-17
C7386 s_3_340 vss 3.13114e-17
C7387 s_3_339 vss 3.13114e-17
C7388 s_3_341 vss 3.13114e-17
C7389 s_3_340 vss 3.13114e-17
C7390 s_3_342 vss 3.13114e-17
C7391 s_3_341 vss 3.13114e-17
C7392 s_3_343 vss 3.13114e-17
C7393 s_3_342 vss 3.13114e-17
C7394 s_3_344 vss 3.13114e-17
C7395 s_3_343 vss 3.13114e-17
C7396 s_3_345 vss 1.40901e-17
C7397 s_3_344 vss 1.40901e-17
C7398 s_3_347 vss 2.95333e-17
C7399 s_3_346 vss 2.95333e-17
C7400 s_3_348 vss 3.71708e-16
C7401 s_3_347 vss 3.71708e-16
C7402 s_3_349 vss 2.15831e-15
C7403 s_3_348 vss 2.15831e-15
C7404 s_3_350 vss 2.15831e-15
C7405 s_3_349 vss 2.15831e-15
C7406 s_3_351 vss 3.71708e-16
C7407 s_3_350 vss 3.71708e-16
C7408 s_3_352 vss 2.95333e-17
C7409 s_3_351 vss 2.95333e-17
C7410 s_3_353 vss 1.40901e-16
C7411 s_3_352 vss 1.40901e-16
C7412 s_3_354 vss 3.13114e-17
C7413 s_3_353 vss 3.13114e-17
C7414 s_3_355 vss 3.13114e-17
C7415 s_3_354 vss 3.13114e-17
C7416 s_3_356 vss 3.13114e-17
C7417 s_3_355 vss 3.13114e-17
C7418 s_3_357 vss 3.13114e-17
C7419 s_3_356 vss 3.13114e-17
C7420 s_3_358 vss 3.13114e-17
C7421 s_3_357 vss 3.13114e-17
C7422 s_3_359 vss 3.13114e-17
C7423 s_3_358 vss 3.13114e-17
C7424 s_3_360 vss 3.13114e-17
C7425 s_3_359 vss 3.13114e-17
C7426 s_3_361 vss 2.42663e-16
C7427 s_3_360 vss 2.42663e-16
C7428 s_3_362 vss 3.13114e-17
C7429 s_3_361 vss 3.13114e-17
C7430 s_3_363 vss 3.13114e-17
C7431 s_3_362 vss 3.13114e-17
C7432 s_3_364 vss 3.13114e-17
C7433 s_3_363 vss 3.13114e-17
C7434 s_3_365 vss 3.13114e-17
C7435 s_3_364 vss 3.13114e-17
C7436 s_3_366 vss 3.13114e-17
C7437 s_3_365 vss 3.13114e-17
C7438 s_3_367 vss 3.13114e-17
C7439 s_3_366 vss 3.13114e-17
C7440 s_3_368 vss 3.13114e-17
C7441 s_3_367 vss 3.13114e-17
C7442 s_3_369 vss 3.13114e-17
C7443 s_3_368 vss 3.13114e-17
C7444 s_3_370 vss 3.13114e-17
C7445 s_3_369 vss 3.13114e-17
C7446 s_3_371 vss 3.13114e-17
C7447 s_3_370 vss 3.13114e-17
C7448 s_3_372 vss 3.13114e-17
C7449 s_3_371 vss 3.13114e-17
C7450 s_3_373 vss 3.13114e-17
C7451 s_3_372 vss 3.13114e-17
C7452 s_3_374 vss 3.13114e-17
C7453 s_3_373 vss 3.13114e-17
C7454 s_3_375 vss 3.13114e-17
C7455 s_3_374 vss 3.13114e-17
C7456 s_3_376 vss 3.13114e-17
C7457 s_3_375 vss 3.13114e-17
C7458 s_3_377 vss 3.13114e-17
C7459 s_3_376 vss 3.13114e-17
C7460 s_3_378 vss 3.13114e-17
C7461 s_3_377 vss 3.13114e-17
C7462 s_3_379 vss 3.13114e-17
C7463 s_3_378 vss 3.13114e-17
C7464 s_3_380 vss 3.13114e-17
C7465 s_3_379 vss 3.13114e-17
C7466 s_3_381 vss 1.40901e-17
C7467 s_3_380 vss 1.40901e-17

R153_1 n5111_3 n5111_153 0.001
R153_2 n5111_123 n5111_8 0.001
R153_3 n5111_7 n5111_11 0.001
R153_4 n5111_152 n5111_18 0.001
R153_5 n5111_115 n5111_27 0.001
R153_6 n5111_26 n5111 0.001
R153_7 n5111_29 n5111 0.001
R153_8 n5111_28 n5111 0.001
R153_9 n5111_24 n5111 0.001
R153_10 n5111_23 n5111 0.001
R153_11 n5111_25 n5111 0.001
R153_12 n5111_166 n5111_31 0.001
R153_13 n5111_168 n5111_31 0.001
R153_14 n5111_167 n5111_31 0.001
R153_15 n5111_169 n5111_31 0.001
R153_16 n5111_164 n5111_31 0.001
R153_17 n5111_165 n5111_31 0.001
R153_18 n5111_162 n5111_31 0.001
R153_19 n5111_163 n5111_31 0.001
R153_20 n5111_158 n5111_31 0.001
R153_21 n5111_161 n5111_31 0.001
R153_22 n5111_159 n5111_31 0.001
R153_23 n5111_160 n5111_31 0.001
R153_24 n5111_155 n5111_31 0.001
R153_25 n5111_156 n5111_31 0.001
R153_26 n5111_157 n5111_31 0.001
R153_27 n5111_122 n5111_33 0.001
R153_28 n5111_32 n5111_36 0.001
R153_29 n5111_114 n5111_46 0.001
R153_30 n5111_45 n5111_41 0.001
R153_31 n5111_47 n5111_41 0.001
R153_32 n5111_48 n5111_41 0.001
R153_33 n5111_44 n5111_41 0.001
R153_34 n5111_43 n5111_41 0.001
R153_35 n5111_42 n5111_41 0.001
R153_36 n5111_140 n5111_50 0.001
R153_37 n5111_141 n5111_50 0.001
R153_38 n5111_142 n5111_50 0.001
R153_39 n5111_143 n5111_50 0.001
R153_40 n5111_138 n5111_50 0.001
R153_41 n5111_139 n5111_50 0.001
R153_42 n5111_136 n5111_50 0.001
R153_43 n5111_137 n5111_50 0.001
R153_44 n5111_132 n5111_50 0.001
R153_45 n5111_135 n5111_50 0.001
R153_46 n5111_133 n5111_50 0.001
R153_47 n5111_134 n5111_50 0.001
R153_48 n5111_129 n5111_50 0.001
R153_49 n5111_130 n5111_50 0.001
R153_50 n5111_131 n5111_50 0.001
R153_51 n5111_150 n5111_53 0.001
R153_52 n5111_121 n5111_58 0.001
R153_53 n5111_57 n5111_61 0.001
R153_54 n5111_149 n5111_68 0.001
R153_55 n5111_120 n5111_73 0.001
R153_56 n5111_72 n5111_76 0.001
R153_57 n5111_148 n5111_83 0.001
R153_58 n5111_119 n5111_88 0.001
R153_59 n5111_87 n5111_91 0.001
R153_60 n5111_147 n5111_98 0.001
R153_61 n5111_118 n5111_103 0.001
R153_62 n5111_102 n5111_106 0.001
R153_63 n5111_145 n5111_111 0.001
R153_64 n5111_124 n5111_112 0.001
R153_65 n5111_125 n5111_113 0.001
R153_66 n5111_144 n5111_116 0.001
R153_67 n5111_127 n5111_117 0.001
R153_68 n5111_35 n5111_34 21.6
R153_69 n5111_38 n5111_35 21.6
R153_70 n5111_39 n5111_38 43.2
R153_71 n5111_40 n5111_39 43.2
R153_72 n5111_10 n5111_9 21.6
R153_73 n5111_13 n5111_10 21.6
R153_74 n5111_14 n5111_13 43.2
R153_75 n5111_15 n5111_14 43.2
R153_76 n5111_60 n5111_59 21.6
R153_77 n5111_63 n5111_60 21.6
R153_78 n5111_64 n5111_63 43.2
R153_79 n5111_65 n5111_64 43.2
R153_80 n5111_75 n5111_74 21.6
R153_81 n5111_78 n5111_75 21.6
R153_82 n5111_79 n5111_78 43.2
R153_83 n5111_80 n5111_79 43.2
R153_84 n5111_90 n5111_89 21.6
R153_85 n5111_93 n5111_90 21.6
R153_86 n5111_94 n5111_93 43.2
R153_87 n5111_95 n5111_94 43.2
R153_88 n5111_105 n5111_104 21.6
R153_89 n5111_108 n5111_105 21.6
R153_90 n5111_109 n5111_108 43.2
R153_91 n5111_110 n5111_109 43.2
R153_92 n5111_37 n5111_35 28.8
R153_93 n5111_12 n5111_10 28.8
R153_94 n5111_62 n5111_60 28.8
R153_95 n5111_77 n5111_75 28.8
R153_96 n5111_92 n5111_90 28.8
R153_97 n5111_107 n5111_105 28.8
R153_98 n5111_37 n5111_36 7.2
R153_99 n5111_12 n5111_11 7.2
R153_100 n5111_62 n5111_61 7.2
R153_101 n5111_77 n5111_76 7.2
R153_102 n5111_92 n5111_91 7.2
R153_103 n5111_107 n5111_106 7.2
R153_104 n5111_43 n5111_42 0.108
R153_105 n5111_44 n5111_43 0.108
R153_106 n5111_45 n5111_44 0.108
R153_107 n5111_46 n5111_45 0.108
R153_108 n5111_47 n5111_46 0.108
R153_109 n5111_48 n5111_47 0.108
R153_110 n5111_49 n5111_48 0.001
R153_111 n5111_24 n5111_23 0.108
R153_112 n5111_25 n5111_24 0.108
R153_113 n5111_26 n5111_25 0.108
R153_114 n5111_27 n5111_26 0.108
R153_115 n5111_28 n5111_27 0.108
R153_116 n5111_29 n5111_28 0.108
R153_117 n5111_30 n5111_29 0.001
R153_118 n5111_33 n5111_32 0.216
R153_119 n5111_8 n5111_7 0.216
R153_120 n5111_58 n5111_57 0.216
R153_121 n5111_73 n5111_72 0.216
R153_122 n5111_88 n5111_87 0.216
R153_123 n5111_103 n5111_102 0.216
R153_124 n5111_17 n5111_16 21.6
R153_125 n5111_19 n5111_17 21.6
R153_126 n5111_20 n5111_19 43.2
R153_127 n5111_21 n5111_20 43.2
R153_128 n5111_52 n5111_51 21.6
R153_129 n5111_54 n5111_52 21.6
R153_130 n5111_55 n5111_54 43.2
R153_131 n5111_56 n5111_55 43.2
R153_132 n5111_67 n5111_66 21.6
R153_133 n5111_69 n5111_67 21.6
R153_134 n5111_70 n5111_69 43.2
R153_135 n5111_71 n5111_70 43.2
R153_136 n5111_97 n5111_96 21.6
R153_137 n5111_99 n5111_97 21.6
R153_138 n5111_100 n5111_99 43.2
R153_139 n5111_101 n5111_100 43.2
R153_140 n5111_82 n5111_81 21.6
R153_141 n5111_84 n5111_82 21.6
R153_142 n5111_85 n5111_84 43.2
R153_143 n5111_86 n5111_85 43.2
R153_144 n5111_18 n5111_17 28.8
R153_145 n5111_53 n5111_52 28.8
R153_146 n5111_68 n5111_67 28.8
R153_147 n5111_98 n5111_97 28.8
R153_148 n5111_83 n5111_82 28.8
R153_149 n5111_112 n5111_111 0.054
R153_150 n5111_113 n5111_112 0.054
R153_151 n5111_114 n5111_113 1.458
R153_152 n5111_115 n5111_114 0.216
R153_153 n5111_117 n5111_116 0.054
R153_154 n5111_118 n5111_117 0.108
R153_155 n5111_119 n5111_118 0.432
R153_156 n5111_120 n5111_119 0.432
R153_157 n5111_121 n5111_120 0.432
R153_158 n5111_122 n5111_121 0.432
R153_159 n5111_123 n5111_122 0.432
R153_160 n5111_124 n5111_145 0.108
R153_161 n5111_125 n5111_124 0.108
R153_162 n5111_126 n5111_125 0.001
R153_163 n5111_127 n5111_144 0.108
R153_164 n5111_128 n5111_127 0.001
R153_165 n5111_129 n5111_150 0.648
R153_166 n5111_130 n5111_129 0.108
R153_167 n5111_131 n5111_130 0.108
R153_168 n5111_132 n5111_131 0.108
R153_169 n5111_133 n5111_132 0.108
R153_170 n5111_134 n5111_133 0.108
R153_171 n5111_135 n5111_134 0.108
R153_172 n5111_136 n5111_135 0.108
R153_173 n5111_137 n5111_136 0.108
R153_174 n5111_138 n5111_137 0.108
R153_175 n5111_139 n5111_138 0.108
R153_176 n5111_140 n5111_139 0.108
R153_177 n5111_141 n5111_140 0.108
R153_178 n5111_142 n5111_141 0.108
R153_179 n5111_143 n5111_142 0.108
R153_180 n5111_155 n5111_151 0.648
R153_181 n5111_156 n5111_155 0.108
R153_182 n5111_157 n5111_156 0.108
R153_183 n5111_158 n5111_157 0.108
R153_184 n5111_159 n5111_158 0.108
R153_185 n5111_160 n5111_159 0.108
R153_186 n5111_161 n5111_160 0.108
R153_187 n5111_162 n5111_161 0.108
R153_188 n5111_163 n5111_162 0.108
R153_189 n5111_164 n5111_163 0.108
R153_190 n5111_165 n5111_164 0.108
R153_191 n5111_166 n5111_165 0.108
R153_192 n5111_167 n5111_166 0.108
R153_193 n5111_168 n5111_167 0.108
R153_194 n5111_169 n5111_168 0.108
R153_195 n5111_146 n5111_144 3.024
R153_196 n5111_145 n5111_146 3.348
R153_197 n5111_147 n5111_146 0.432
R153_198 n5111_148 n5111_147 0.648
R153_199 n5111_149 n5111_148 0.648
R153_200 n5111_150 n5111_149 0.648
R153_201 n5111_151 n5111_150 0.324
R153_202 n5111_152 n5111_151 0.216
R153_203 n5111_153 n5111_152 0.648
R153_204 n5111_154 n5111_153 0.001
R153_205 n5111_2 n5111_1 21.6
R153_206 n5111_4 n5111_2 21.6
R153_207 n5111_5 n5111_4 43.2
R153_208 n5111_6 n5111_5 43.2
R153_209 n5111_3 n5111_2 28.8

C7468 n5111_35 vss 2.34738e-17
C7469 n5111_34 vss 2.34738e-17
C7470 n5111_38 vss 2.34738e-17
C7471 n5111_35 vss 2.34738e-17
C7472 n5111_39 vss 4.69476e-17
C7473 n5111_38 vss 4.69476e-17
C7474 n5111_40 vss 4.69476e-17
C7475 n5111_39 vss 4.69476e-17
C7476 n5111_10 vss 2.34738e-17
C7477 n5111_9 vss 2.34738e-17
C7478 n5111_13 vss 2.34738e-17
C7479 n5111_10 vss 2.34738e-17
C7480 n5111_14 vss 4.69476e-17
C7481 n5111_13 vss 4.69476e-17
C7482 n5111_15 vss 4.69476e-17
C7483 n5111_14 vss 4.69476e-17
C7484 n5111_60 vss 2.34738e-17
C7485 n5111_59 vss 2.34738e-17
C7486 n5111_63 vss 2.34738e-17
C7487 n5111_60 vss 2.34738e-17
C7488 n5111_64 vss 4.69476e-17
C7489 n5111_63 vss 4.69476e-17
C7490 n5111_65 vss 4.69476e-17
C7491 n5111_64 vss 4.69476e-17
C7492 n5111_75 vss 2.34738e-17
C7493 n5111_74 vss 2.34738e-17
C7494 n5111_78 vss 2.34738e-17
C7495 n5111_75 vss 2.34738e-17
C7496 n5111_79 vss 4.69476e-17
C7497 n5111_78 vss 4.69476e-17
C7498 n5111_80 vss 4.69476e-17
C7499 n5111_79 vss 4.69476e-17
C7500 n5111_90 vss 2.34738e-17
C7501 n5111_89 vss 2.34738e-17
C7502 n5111_93 vss 2.34738e-17
C7503 n5111_90 vss 2.34738e-17
C7504 n5111_94 vss 4.69476e-17
C7505 n5111_93 vss 4.69476e-17
C7506 n5111_95 vss 4.69476e-17
C7507 n5111_94 vss 4.69476e-17
C7508 n5111_105 vss 2.34738e-17
C7509 n5111_104 vss 2.34738e-17
C7510 n5111_108 vss 2.34738e-17
C7511 n5111_105 vss 2.34738e-17
C7512 n5111_109 vss 4.69476e-17
C7513 n5111_108 vss 4.69476e-17
C7514 n5111_110 vss 4.69476e-17
C7515 n5111_109 vss 4.69476e-17
C7516 n5111_37 vss 7.33536e-17
C7517 n5111_35 vss 7.33536e-17
C7518 n5111_12 vss 7.33536e-17
C7519 n5111_10 vss 7.33536e-17
C7520 n5111_62 vss 7.33536e-17
C7521 n5111_60 vss 7.33536e-17
C7522 n5111_77 vss 7.33536e-17
C7523 n5111_75 vss 7.33536e-17
C7524 n5111_92 vss 7.33536e-17
C7525 n5111_90 vss 7.33536e-17
C7526 n5111_107 vss 7.33536e-17
C7527 n5111_105 vss 7.33536e-17
C7528 n5111_37 vss 5.2569e-17
C7529 n5111_36 vss 5.2569e-17
C7530 n5111_12 vss 5.2569e-17
C7531 n5111_11 vss 5.2569e-17
C7532 n5111_62 vss 5.2569e-17
C7533 n5111_61 vss 5.2569e-17
C7534 n5111_77 vss 5.2569e-17
C7535 n5111_76 vss 5.2569e-17
C7536 n5111_92 vss 5.2569e-17
C7537 n5111_91 vss 5.2569e-17
C7538 n5111_107 vss 5.2569e-17
C7539 n5111_106 vss 5.2569e-17
C7540 n5111_43 vss 2.92378e-17
C7541 n5111_42 vss 2.92378e-17
C7542 n5111_44 vss 2.92378e-17
C7543 n5111_43 vss 2.92378e-17
C7544 n5111_45 vss 2.92378e-17
C7545 n5111_44 vss 2.92378e-17
C7546 n5111_46 vss 3.65472e-17
C7547 n5111_45 vss 3.65472e-17
C7548 n5111_47 vss 2.92378e-17
C7549 n5111_46 vss 2.92378e-17
C7550 n5111_48 vss 3.65472e-17
C7551 n5111_47 vss 3.65472e-17
C7552 n5111_49 vss 1.3157e-17
C7553 n5111_48 vss 1.3157e-17
C7554 n5111_24 vss 2.92378e-17
C7555 n5111_23 vss 2.92378e-17
C7556 n5111_25 vss 2.92378e-17
C7557 n5111_24 vss 2.92378e-17
C7558 n5111_26 vss 2.92378e-17
C7559 n5111_25 vss 2.92378e-17
C7560 n5111_27 vss 3.65472e-17
C7561 n5111_26 vss 3.65472e-17
C7562 n5111_28 vss 2.92378e-17
C7563 n5111_27 vss 2.92378e-17
C7564 n5111_29 vss 3.65472e-17
C7565 n5111_28 vss 3.65472e-17
C7566 n5111_30 vss 1.3157e-17
C7567 n5111_29 vss 1.3157e-17
C7568 n5111_33 vss 4.38566e-17
C7569 n5111_32 vss 4.38566e-17
C7570 n5111_8 vss 4.38566e-17
C7571 n5111_7 vss 4.38566e-17
C7572 n5111_58 vss 4.38566e-17
C7573 n5111_57 vss 4.38566e-17
C7574 n5111_73 vss 4.38566e-17
C7575 n5111_72 vss 4.38566e-17
C7576 n5111_88 vss 4.38566e-17
C7577 n5111_87 vss 4.38566e-17
C7578 n5111_103 vss 4.38566e-17
C7579 n5111_102 vss 4.38566e-17
C7580 n5111_17 vss 2.34738e-17
C7581 n5111_16 vss 2.34738e-17
C7582 n5111_19 vss 2.34738e-17
C7583 n5111_17 vss 2.34738e-17
C7584 n5111_20 vss 4.69476e-17
C7585 n5111_19 vss 4.69476e-17
C7586 n5111_21 vss 4.69476e-17
C7587 n5111_20 vss 4.69476e-17
C7588 n5111_52 vss 2.34738e-17
C7589 n5111_51 vss 2.34738e-17
C7590 n5111_54 vss 2.34738e-17
C7591 n5111_52 vss 2.34738e-17
C7592 n5111_55 vss 4.69476e-17
C7593 n5111_54 vss 4.69476e-17
C7594 n5111_56 vss 4.69476e-17
C7595 n5111_55 vss 4.69476e-17
C7596 n5111_67 vss 2.34738e-17
C7597 n5111_66 vss 2.34738e-17
C7598 n5111_69 vss 2.34738e-17
C7599 n5111_67 vss 2.34738e-17
C7600 n5111_70 vss 4.69476e-17
C7601 n5111_69 vss 4.69476e-17
C7602 n5111_71 vss 4.69476e-17
C7603 n5111_70 vss 4.69476e-17
C7604 n5111_97 vss 2.34738e-17
C7605 n5111_96 vss 2.34738e-17
C7606 n5111_99 vss 2.34738e-17
C7607 n5111_97 vss 2.34738e-17
C7608 n5111_100 vss 4.69476e-17
C7609 n5111_99 vss 4.69476e-17
C7610 n5111_101 vss 4.69476e-17
C7611 n5111_100 vss 4.69476e-17
C7612 n5111_82 vss 2.34738e-17
C7613 n5111_81 vss 2.34738e-17
C7614 n5111_84 vss 2.34738e-17
C7615 n5111_82 vss 2.34738e-17
C7616 n5111_85 vss 4.69476e-17
C7617 n5111_84 vss 4.69476e-17
C7618 n5111_86 vss 4.69476e-17
C7619 n5111_85 vss 4.69476e-17
C7620 n5111_18 vss 7.33536e-17
C7621 n5111_17 vss 7.33536e-17
C7622 n5111_53 vss 7.33536e-17
C7623 n5111_52 vss 7.33536e-17
C7624 n5111_68 vss 7.33536e-17
C7625 n5111_67 vss 7.33536e-17
C7626 n5111_98 vss 7.33536e-17
C7627 n5111_97 vss 7.33536e-17
C7628 n5111_83 vss 7.33536e-17
C7629 n5111_82 vss 7.33536e-17
C7630 n5111_112 vss 2.60496e-17
C7631 n5111_111 vss 2.60496e-17
C7632 n5111_113 vss 2.60496e-17
C7633 n5111_112 vss 2.60496e-17
C7634 n5111_114 vss 5.40529e-16
C7635 n5111_113 vss 5.40529e-16
C7636 n5111_115 vss 7.81488e-17
C7637 n5111_114 vss 7.81488e-17
C7638 n5111_117 vss 3.2562e-17
C7639 n5111_116 vss 3.2562e-17
C7640 n5111_118 vss 4.55868e-17
C7641 n5111_117 vss 4.55868e-17
C7642 n5111_119 vss 1.56298e-16
C7643 n5111_118 vss 1.56298e-16
C7644 n5111_120 vss 1.56298e-16
C7645 n5111_119 vss 1.56298e-16
C7646 n5111_121 vss 1.56298e-16
C7647 n5111_120 vss 1.56298e-16
C7648 n5111_122 vss 1.56298e-16
C7649 n5111_121 vss 1.56298e-16
C7650 n5111_123 vss 1.56298e-16
C7651 n5111_122 vss 1.56298e-16
C7652 n5111_124 vss 3.13114e-17
C7653 n5111_145 vss 3.13114e-17
C7654 n5111_125 vss 3.13114e-17
C7655 n5111_124 vss 3.13114e-17
C7656 n5111_126 vss 1.40901e-17
C7657 n5111_125 vss 1.40901e-17
C7658 n5111_127 vss 3.91392e-17
C7659 n5111_144 vss 3.91392e-17
C7660 n5111_128 vss 1.40901e-17
C7661 n5111_127 vss 1.40901e-17
C7662 n5111_129 vss 1.20606e-16
C7663 n5111_150 vss 1.20606e-16
C7664 n5111_130 vss 2.92378e-17
C7665 n5111_129 vss 2.92378e-17
C7666 n5111_131 vss 2.92378e-17
C7667 n5111_130 vss 2.92378e-17
C7668 n5111_132 vss 2.92378e-17
C7669 n5111_131 vss 2.92378e-17
C7670 n5111_133 vss 2.92378e-17
C7671 n5111_132 vss 2.92378e-17
C7672 n5111_134 vss 2.92378e-17
C7673 n5111_133 vss 2.92378e-17
C7674 n5111_135 vss 2.92378e-17
C7675 n5111_134 vss 2.92378e-17
C7676 n5111_136 vss 2.92378e-17
C7677 n5111_135 vss 2.92378e-17
C7678 n5111_137 vss 2.92378e-17
C7679 n5111_136 vss 2.92378e-17
C7680 n5111_138 vss 2.92378e-17
C7681 n5111_137 vss 2.92378e-17
C7682 n5111_139 vss 2.92378e-17
C7683 n5111_138 vss 2.92378e-17
C7684 n5111_140 vss 2.92378e-17
C7685 n5111_139 vss 2.92378e-17
C7686 n5111_141 vss 2.92378e-17
C7687 n5111_140 vss 2.92378e-17
C7688 n5111_142 vss 2.92378e-17
C7689 n5111_141 vss 2.92378e-17
C7690 n5111_143 vss 2.92378e-17
C7691 n5111_142 vss 2.92378e-17
C7692 n5111_155 vss 1.20606e-16
C7693 n5111_151 vss 1.20606e-16
C7694 n5111_156 vss 2.92378e-17
C7695 n5111_155 vss 2.92378e-17
C7696 n5111_157 vss 2.92378e-17
C7697 n5111_156 vss 2.92378e-17
C7698 n5111_158 vss 2.92378e-17
C7699 n5111_157 vss 2.92378e-17
C7700 n5111_159 vss 2.92378e-17
C7701 n5111_158 vss 2.92378e-17
C7702 n5111_160 vss 2.92378e-17
C7703 n5111_159 vss 2.92378e-17
C7704 n5111_161 vss 2.92378e-17
C7705 n5111_160 vss 2.92378e-17
C7706 n5111_162 vss 2.92378e-17
C7707 n5111_161 vss 2.92378e-17
C7708 n5111_163 vss 2.92378e-17
C7709 n5111_162 vss 2.92378e-17
C7710 n5111_164 vss 2.92378e-17
C7711 n5111_163 vss 2.92378e-17
C7712 n5111_165 vss 2.92378e-17
C7713 n5111_164 vss 2.92378e-17
C7714 n5111_166 vss 2.92378e-17
C7715 n5111_165 vss 2.92378e-17
C7716 n5111_167 vss 2.92378e-17
C7717 n5111_166 vss 2.92378e-17
C7718 n5111_168 vss 2.92378e-17
C7719 n5111_167 vss 2.92378e-17
C7720 n5111_169 vss 2.92378e-17
C7721 n5111_168 vss 2.92378e-17
C7722 n5111_146 vss 7.94526e-16
C7723 n5111_144 vss 7.94526e-16
C7724 n5111_145 vss 8.96288e-16
C7725 n5111_146 vss 8.96288e-16
C7726 n5111_147 vss 1.33073e-16
C7727 n5111_146 vss 1.33073e-16
C7728 n5111_148 vss 1.87868e-16
C7729 n5111_147 vss 1.87868e-16
C7730 n5111_149 vss 1.87868e-16
C7731 n5111_148 vss 1.87868e-16
C7732 n5111_150 vss 1.95696e-16
C7733 n5111_149 vss 1.95696e-16
C7734 n5111_151 vss 1.01762e-16
C7735 n5111_150 vss 1.01762e-16
C7736 n5111_152 vss 7.82784e-17
C7737 n5111_151 vss 7.82784e-17
C7738 n5111_153 vss 1.87868e-16
C7739 n5111_152 vss 1.87868e-16
C7740 n5111_154 vss 1.40901e-17
C7741 n5111_153 vss 1.40901e-17
C7742 n5111_2 vss 2.34738e-17
C7743 n5111_1 vss 2.34738e-17
C7744 n5111_4 vss 2.34738e-17
C7745 n5111_2 vss 2.34738e-17
C7746 n5111_5 vss 4.69476e-17
C7747 n5111_4 vss 4.69476e-17
C7748 n5111_6 vss 4.69476e-17
C7749 n5111_5 vss 4.69476e-17
C7750 n5111_3 vss 7.33536e-17
C7751 n5111_2 vss 7.33536e-17

R154_1 n5139_2 n5139_33 0.001
R154_2 n5139_20 n5139_6 0.001
R154_3 n5139_1 n5139_32 0.001
R154_4 n5139_29 n5139_5 0.001
R154_5 n5139_38 n5139_9 0.001
R154_6 n5139_39 n5139_9 0.001
R154_7 n5139_36 n5139_9 0.001
R154_8 n5139_37 n5139_9 0.001
R154_9 n5139_35 n5139_9 0.001
R154_10 n5139_27 n5139_10 0.001
R154_11 n5139_28 n5139_10 0.001
R154_12 n5139_26 n5139_10 0.001
R154_13 n5139_24 n5139_10 0.001
R154_14 n5139_25 n5139_12 0.001
R154_15 n5139_18 n5139_13 0.001
R154_16 n5139_17 n5139_13 0.001
R154_17 n5139_16 n5139_13 0.001
R154_18 n5139_11 n5139_15 0.001
R154_19 n5139_14 n5139_13 0.001
R154_20 n5139_6 n5139_5 7.2
R154_21 n5139_7 n5139_6 21.6
R154_22 n5139 n5139_7 0.001
R154_23 n5139_14 n5139_22 0.324
R154_24 n5139_15 n5139_14 0.108
R154_25 n5139_16 n5139_15 0.108
R154_26 n5139_17 n5139_16 0.108
R154_27 n5139_18 n5139_17 0.108
R154_28 n5139_19 n5139_18 0.001
R154_29 n5139_12 n5139_11 0.216
R154_30 n5139_20 n5139_29 0.108
R154_31 n5139_21 n5139_20 0.001
R154_32 n5139_23 n5139_22 0.324
R154_33 n5139_24 n5139_23 0.324
R154_34 n5139_25 n5139_24 0.108
R154_35 n5139_26 n5139_25 0.108
R154_36 n5139_27 n5139_26 0.108
R154_37 n5139_28 n5139_27 0.108
R154_38 n5139_29 n5139_28 0.108
R154_39 n5139_30 n5139_29 0.216
R154_40 n5139_31 n5139_30 0.108
R154_41 n5139_32 n5139_31 0.216
R154_42 n5139_35 n5139_32 0.108
R154_43 n5139_36 n5139_35 0.108
R154_44 n5139_37 n5139_36 0.108
R154_45 n5139_38 n5139_37 0.108
R154_46 n5139_39 n5139_38 0.108
R154_47 n5139_40 n5139_39 0.001
R154_48 n5139_33 n5139_32 0.108
R154_49 n5139_34 n5139_33 0.001
R154_50 n5139_2 n5139_1 7.2
R154_51 n5139_3 n5139_2 21.6
R154_52 n5139_4 n5139_3 0.001

C7752 n5139_6 vss 4.20552e-17
C7753 n5139_5 vss 4.20552e-17
C7754 n5139_7 vss 9.46242e-17
C7755 n5139_6 vss 9.46242e-17
C7756 n5139 vss 3.05111e-16
C7757 n5139_7 vss 3.05111e-16
C7758 n5139_14 vss 1.0959e-16
C7759 n5139_22 vss 1.0959e-16
C7760 n5139_15 vss 3.91392e-17
C7761 n5139_14 vss 3.91392e-17
C7762 n5139_16 vss 3.91392e-17
C7763 n5139_15 vss 3.91392e-17
C7764 n5139_17 vss 3.91392e-17
C7765 n5139_16 vss 3.91392e-17
C7766 n5139_18 vss 3.91392e-17
C7767 n5139_17 vss 3.91392e-17
C7768 n5139_19 vss 1.40901e-17
C7769 n5139_18 vss 1.40901e-17
C7770 n5139_12 vss 7.81488e-17
C7771 n5139_11 vss 7.81488e-17
C7772 n5139_20 vss 3.71822e-17
C7773 n5139_29 vss 3.71822e-17
C7774 n5139_21 vss 1.40901e-17
C7775 n5139_20 vss 1.40901e-17
C7776 n5139_23 vss 9.39341e-17
C7777 n5139_22 vss 9.39341e-17
C7778 n5139_24 vss 1.0959e-16
C7779 n5139_23 vss 1.0959e-16
C7780 n5139_25 vss 3.91392e-17
C7781 n5139_24 vss 3.91392e-17
C7782 n5139_26 vss 3.91392e-17
C7783 n5139_25 vss 3.91392e-17
C7784 n5139_27 vss 3.91392e-17
C7785 n5139_26 vss 3.91392e-17
C7786 n5139_28 vss 3.91392e-17
C7787 n5139_27 vss 3.91392e-17
C7788 n5139_29 vss 4.6967e-17
C7789 n5139_28 vss 4.6967e-17
C7790 n5139_30 vss 5.63604e-17
C7791 n5139_29 vss 5.63604e-17
C7792 n5139_31 vss 2.81802e-17
C7793 n5139_30 vss 2.81802e-17
C7794 n5139_32 vss 6.41883e-17
C7795 n5139_31 vss 6.41883e-17
C7796 n5139_35 vss 4.6967e-17
C7797 n5139_32 vss 4.6967e-17
C7798 n5139_36 vss 3.91392e-17
C7799 n5139_35 vss 3.91392e-17
C7800 n5139_37 vss 4.6967e-17
C7801 n5139_36 vss 4.6967e-17
C7802 n5139_38 vss 3.91392e-17
C7803 n5139_37 vss 3.91392e-17
C7804 n5139_39 vss 3.91392e-17
C7805 n5139_38 vss 3.91392e-17
C7806 n5139_40 vss 1.40901e-17
C7807 n5139_39 vss 1.40901e-17
C7808 n5139_33 vss 3.71822e-17
C7809 n5139_32 vss 3.71822e-17
C7810 n5139_34 vss 1.40901e-17
C7811 n5139_33 vss 1.40901e-17
C7812 n5139_2 vss 4.20552e-17
C7813 n5139_1 vss 4.20552e-17
C7814 n5139_3 vss 9.46242e-17
C7815 n5139_2 vss 9.46242e-17
C7816 n5139_4 vss 5.47139e-16
C7817 n5139_3 vss 5.47139e-16

R155_1 aa_1_1 aa_1_34 0.001
R155_2 aa_1_1 aa_1_33 0.001
R155_3 aa_1_1 aa_1_38 0.001
R155_4 aa_1_1 aa_1_37 0.001
R155_5 aa_1_1 aa_1_35 0.001
R155_6 aa_1_1 aa_1_36 0.001
R155_7 aa_1_1 aa_1_39 0.001
R155_8 aa_1_1 aa_1_40 0.001
R155_9 aa_1_1 aa_1_41 0.001
R155_10 aa_1_1 aa_1_46 0.001
R155_11 aa_1_1 aa_1_45 0.001
R155_12 aa_1_1 aa_1_44 0.001
R155_13 aa_1_1 aa_1_43 0.001
R155_14 aa_1_1 aa_1_42 0.001
R155_15 aa_1_29 aa_1_2 0.001
R155_16 aa_1_32 aa_1_2 0.001
R155_17 aa_1_30 aa_1_2 0.001
R155_18 aa_1_31 aa_1_2 0.001
R155_19 aa_1_28 aa_1_4 0.001
R155_20 aa_1_26 aa_1_7 0.001
R155_21 aa_1_9 aa_1_13 0.001
R155_22 aa_1_12 aa_1_25 0.001
R155_23 aa_1_6 aa_1_11 0.001
R155_24 aa_1_10 aa_1_8 0.001
R155_25 aa_1_20 aa_1_15 0.001
R155_26 aa_1_14 aa_1_17 0.001
R155_27 aa_1_17 aa_1_16 72
R155_28 aa_1 aa_1_17 43.2
R155_29 aa_1_15 aa_1_14 0.108
R155_30 aa_1_20 aa_1_19 0.756
R155_31 aa_1_21 aa_1_20 0.324
R155_32 aa_1_22 aa_1_21 0.054
R155_33 aa_1_23 aa_1_22 0.648
R155_34 aa_1_24 aa_1_23 0.054
R155_35 aa_1_25 aa_1_24 0.486
R155_36 aa_1_13 aa_1_12 12.42
R155_37 aa_1_9 aa_1_8 0.81
R155_38 aa_1_11 aa_1_10 9.072
R155_39 aa_1_7 aa_1_6 2.7
R155_40 aa_1_4 aa_1_3 0.054
R155_41 aa_1_5 aa_1_4 0.001
R155_42 aa_1_27 aa_1_26 0.864
R155_43 aa_1_28 aa_1_27 0.001
R155_44 aa_1_29 aa_1_28 0.54
R155_45 aa_1_30 aa_1_29 0.108
R155_46 aa_1_31 aa_1_30 0.108
R155_47 aa_1_32 aa_1_31 0.108
R155_48 aa_1_33 aa_1_32 0.864
R155_49 aa_1_34 aa_1_33 0.108
R155_50 aa_1_35 aa_1_34 0.108
R155_51 aa_1_36 aa_1_35 0.108
R155_52 aa_1_37 aa_1_36 0.108
R155_53 aa_1_38 aa_1_37 0.108
R155_54 aa_1_39 aa_1_38 0.108
R155_55 aa_1_40 aa_1_39 0.108
R155_56 aa_1_41 aa_1_40 0.108
R155_57 aa_1_42 aa_1_41 0.108
R155_58 aa_1_43 aa_1_42 0.108
R155_59 aa_1_44 aa_1_43 0.108
R155_60 aa_1_45 aa_1_44 0.108
R155_61 aa_1_46 aa_1_45 0.108
R155_62 aa_1_47 aa_1_46 0.001

C7818 aa_1_17 vss 8.21582e-17
C7819 aa_1_16 vss 8.21582e-17
C7820 aa_1 vss 5.086e-17
C7821 aa_1_17 vss 5.086e-17
C7822 aa_1_15 vss 3.65472e-17
C7823 aa_1_14 vss 3.65472e-17
C7824 aa_1_20 vss 1.78524e-16
C7825 aa_1_19 vss 1.78524e-16
C7826 aa_1_21 vss 8.0028e-17
C7827 aa_1_20 vss 8.0028e-17
C7828 aa_1_22 vss 1.2312e-17
C7829 aa_1_21 vss 1.2312e-17
C7830 aa_1_23 vss 1.539e-16
C7831 aa_1_22 vss 1.539e-16
C7832 aa_1_24 vss 1.2312e-17
C7833 aa_1_23 vss 1.2312e-17
C7834 aa_1_25 vss 1.16964e-16
C7835 aa_1_24 vss 1.16964e-16
C7836 aa_1_13 vss 1.25634e-15
C7837 aa_1_12 vss 1.25634e-15
C7838 aa_1_9 vss 1.8468e-16
C7839 aa_1_8 vss 1.8468e-16
C7840 aa_1_11 vss 9.1679e-16
C7841 aa_1_10 vss 9.1679e-16
C7842 aa_1_7 vss 6.21756e-16
C7843 aa_1_6 vss 6.21756e-16
C7844 aa_1_4 vss 1.95372e-17
C7845 aa_1_3 vss 1.95372e-17
C7846 aa_1_5 vss 1.30248e-17
C7847 aa_1_4 vss 1.30248e-17
C7848 aa_1_27 vss 9.64328e-17
C7849 aa_1_26 vss 9.64328e-17
C7850 aa_1_28 vss 2.1918e-17
C7851 aa_1_27 vss 2.1918e-17
C7852 aa_1_29 vss 1.64385e-16
C7853 aa_1_28 vss 1.64385e-16
C7854 aa_1_30 vss 3.91392e-17
C7855 aa_1_29 vss 3.91392e-17
C7856 aa_1_31 vss 3.91392e-17
C7857 aa_1_30 vss 3.91392e-17
C7858 aa_1_32 vss 3.91392e-17
C7859 aa_1_31 vss 3.91392e-17
C7860 aa_1_33 vss 2.42663e-16
C7861 aa_1_32 vss 2.42663e-16
C7862 aa_1_34 vss 3.13114e-17
C7863 aa_1_33 vss 3.13114e-17
C7864 aa_1_35 vss 3.13114e-17
C7865 aa_1_34 vss 3.13114e-17
C7866 aa_1_36 vss 3.13114e-17
C7867 aa_1_35 vss 3.13114e-17
C7868 aa_1_37 vss 3.13114e-17
C7869 aa_1_36 vss 3.13114e-17
C7870 aa_1_38 vss 3.13114e-17
C7871 aa_1_37 vss 3.13114e-17
C7872 aa_1_39 vss 3.13114e-17
C7873 aa_1_38 vss 3.13114e-17
C7874 aa_1_40 vss 3.13114e-17
C7875 aa_1_39 vss 3.13114e-17
C7876 aa_1_41 vss 3.13114e-17
C7877 aa_1_40 vss 3.13114e-17
C7878 aa_1_42 vss 3.13114e-17
C7879 aa_1_41 vss 3.13114e-17
C7880 aa_1_43 vss 3.13114e-17
C7881 aa_1_42 vss 3.13114e-17
C7882 aa_1_44 vss 3.13114e-17
C7883 aa_1_43 vss 3.13114e-17
C7884 aa_1_45 vss 3.13114e-17
C7885 aa_1_44 vss 3.13114e-17
C7886 aa_1_46 vss 3.13114e-17
C7887 aa_1_45 vss 3.13114e-17
C7888 aa_1_47 vss 1.40901e-17
C7889 aa_1_46 vss 1.40901e-17

R4_1 a_1_50 a_1_1 0.001
R4_2 a_1_48 a_1_1 0.001
R4_3 a_1_49 a_1_1 0.001
R4_4 a_1_47 a_1_1 0.001
R4_5 a_1_46 a_1_1 0.001
R4_6 a_1_45 a_1_1 0.001
R4_7 a_1_44 a_1_1 0.001
R4_8 a_1_43 a_1_1 0.001
R4_9 a_1_42 a_1_2 0.001
R4_10 a_1_41 a_1_2 0.001
R4_11 a_1_39 a_1_2 0.001
R4_12 a_1_40 a_1_2 0.001
R4_13 a_1_36 a_1_2 0.001
R4_14 a_1_38 a_1_2 0.001
R4_15 a_1_37 a_1_2 0.001
R4_16 a_1_34 a_1_2 0.001
R4_17 a_1_35 a_1_2 0.001
R4_18 a_1_33 a_1_2 0.001
R4_19 a_1_32 a_1_2 0.001
R4_20 a_1_30 a_1_2 0.001
R4_21 a_1_31 a_1_2 0.001
R4_22 a_1_29 a_1_2 0.001
R4_23 a_1_28 a_1_2 0.001
R4_24 a_1_27 a_1_2 0.001
R4_25 a_1_26 a_1_2 0.001
R4_26 a_1_25 a_1_2 0.001
R4_27 a_1_24 a_1_2 0.001
R4_28 a_1_23 a_1_2 0.001
R4_29 a_1_79 a_1_3 0.001
R4_30 a_1_77 a_1_3 0.001
R4_31 a_1_78 a_1_3 0.001
R4_32 a_1_75 a_1_3 0.001
R4_33 a_1_76 a_1_3 0.001
R4_34 a_1_73 a_1_3 0.001
R4_35 a_1_74 a_1_3 0.001
R4_36 a_1_72 a_1_3 0.001
R4_37 a_1_70 a_1_4 0.001
R4_38 a_1_71 a_1_4 0.001
R4_39 a_1_68 a_1_4 0.001
R4_40 a_1_69 a_1_4 0.001
R4_41 a_1_65 a_1_4 0.001
R4_42 a_1_67 a_1_4 0.001
R4_43 a_1_66 a_1_4 0.001
R4_44 a_1_64 a_1_4 0.001
R4_45 a_1_63 a_1_4 0.001
R4_46 a_1_62 a_1_4 0.001
R4_47 a_1_61 a_1_4 0.001
R4_48 a_1_59 a_1_4 0.001
R4_49 a_1_60 a_1_4 0.001
R4_50 a_1_58 a_1_4 0.001
R4_51 a_1_57 a_1_4 0.001
R4_52 a_1_55 a_1_4 0.001
R4_53 a_1_56 a_1_4 0.001
R4_54 a_1_54 a_1_4 0.001
R4_55 a_1_53 a_1_4 0.001
R4_56 a_1_52 a_1_4 0.001
R4_57 a_1_14 a_1_5 0.001
R4_58 a_1_13 a_1_8 0.001
R4_59 a_1 a_1_11 0.001
R4_60 a_1_6 a_1_5 21.6
R4_61 a_1_8 a_1_7 7.2
R4_62 a_1_9 a_1_8 7.2
R4_63 a_1_10 a_1_9 14.4
R4_64 a_1_13 a_1_12 0.001
R4_65 a_1_16 a_1_13 0.216
R4_66 a_1_14 a_1_16 0.216
R4_67 a_1_15 a_1_14 0.001
R4_68 a_1_16 a_1_17 0.324
R4_69 a_1_18 a_1_17 2.268
R4_70 a_1_19 a_1_18 1.08
R4_71 a_1_20 a_1_19 0.001
R4_72 a_1_21 a_1_20 0.001
R4_73 a_1_51 a_1_21 0.216
R4_74 a_1_23 a_1_22 0.001
R4_75 a_1_24 a_1_23 0.108
R4_76 a_1_25 a_1_24 0.108
R4_77 a_1_26 a_1_25 0.108
R4_78 a_1_27 a_1_26 0.108
R4_79 a_1_28 a_1_27 0.108
R4_80 a_1_29 a_1_28 0.108
R4_81 a_1_30 a_1_29 0.108
R4_82 a_1_31 a_1_30 0.108
R4_83 a_1_32 a_1_31 0.108
R4_84 a_1_33 a_1_32 0.108
R4_85 a_1_34 a_1_33 0.108
R4_86 a_1_35 a_1_34 0.108
R4_87 a_1_36 a_1_35 0.108
R4_88 a_1_37 a_1_36 0.108
R4_89 a_1_38 a_1_37 0.108
R4_90 a_1_39 a_1_38 0.108
R4_91 a_1_40 a_1_39 0.108
R4_92 a_1_41 a_1_40 0.108
R4_93 a_1_42 a_1_41 0.108
R4_94 a_1_43 a_1_42 0.864
R4_95 a_1_44 a_1_43 0.108
R4_96 a_1_45 a_1_44 0.108
R4_97 a_1_46 a_1_45 0.108
R4_98 a_1_47 a_1_46 0.108
R4_99 a_1_48 a_1_47 0.108
R4_100 a_1_49 a_1_48 0.108
R4_101 a_1_50 a_1_49 0.108
R4_102 a_1_81 a_1_50 0.54
R4_103 a_1_52 a_1_51 0.001
R4_104 a_1_53 a_1_52 0.108
R4_105 a_1_54 a_1_53 0.108
R4_106 a_1_55 a_1_54 0.108
R4_107 a_1_56 a_1_55 0.108
R4_108 a_1_57 a_1_56 0.108
R4_109 a_1_58 a_1_57 0.108
R4_110 a_1_59 a_1_58 0.108
R4_111 a_1_60 a_1_59 0.108
R4_112 a_1_61 a_1_60 0.108
R4_113 a_1_62 a_1_61 0.108
R4_114 a_1_63 a_1_62 0.108
R4_115 a_1_64 a_1_63 0.108
R4_116 a_1_65 a_1_64 0.108
R4_117 a_1_66 a_1_65 0.108
R4_118 a_1_67 a_1_66 0.108
R4_119 a_1_68 a_1_67 0.108
R4_120 a_1_69 a_1_68 0.108
R4_121 a_1_70 a_1_69 0.108
R4_122 a_1_71 a_1_70 0.108
R4_123 a_1_72 a_1_71 0.864
R4_124 a_1_73 a_1_72 0.108
R4_125 a_1_74 a_1_73 0.108
R4_126 a_1_75 a_1_74 0.108
R4_127 a_1_76 a_1_75 0.108
R4_128 a_1_77 a_1_76 0.108
R4_129 a_1_78 a_1_77 0.108
R4_130 a_1_79 a_1_78 0.108
R4_131 a_1_82 a_1_79 0.54
R4_132 a_1_82 a_1_80 0.001
R4_133 a_1_81 a_1_82 0.108
R4_134 a_1_83 a_1_82 0.54
R4_135 a_1_84 a_1_83 0.001
R4_136 a_1 a_1_84 0.001

C7890 a_1_6 vss 9.46242e-17
C7891 a_1_5 vss 9.46242e-17
C7892 a_1_8 vss 3.15414e-17
C7893 a_1_7 vss 3.15414e-17
C7894 a_1_9 vss 3.15414e-17
C7895 a_1_8 vss 3.15414e-17
C7896 a_1_10 vss 6.30828e-17
C7897 a_1_9 vss 6.30828e-17
C7898 a_1_13 vss 1.40901e-17
C7899 a_1_12 vss 1.40901e-17
C7900 a_1_16 vss 7.82784e-17
C7901 a_1_13 vss 7.82784e-17
C7902 a_1_14 vss 7.04506e-17
C7903 a_1_16 vss 7.04506e-17
C7904 a_1_15 vss 1.40901e-17
C7905 a_1_14 vss 1.40901e-17
C7906 a_1_16 vss 9.39341e-17
C7907 a_1_17 vss 9.39341e-17
C7908 a_1_18 vss 6.18399e-16
C7909 a_1_17 vss 6.18399e-16
C7910 a_1_19 vss 2.97458e-16
C7911 a_1_18 vss 2.97458e-16
C7912 a_1_20 vss 2.50491e-17
C7913 a_1_19 vss 2.50491e-17
C7914 a_1_21 vss 1.25245e-17
C7915 a_1_20 vss 1.25245e-17
C7916 a_1_51 vss 8.14095e-17
C7917 a_1_21 vss 8.14095e-17
C7918 a_1_23 vss 1.40901e-17
C7919 a_1_22 vss 1.40901e-17
C7920 a_1_24 vss 3.13114e-17
C7921 a_1_23 vss 3.13114e-17
C7922 a_1_25 vss 3.13114e-17
C7923 a_1_24 vss 3.13114e-17
C7924 a_1_26 vss 3.13114e-17
C7925 a_1_25 vss 3.13114e-17
C7926 a_1_27 vss 3.13114e-17
C7927 a_1_26 vss 3.13114e-17
C7928 a_1_28 vss 3.13114e-17
C7929 a_1_27 vss 3.13114e-17
C7930 a_1_29 vss 3.13114e-17
C7931 a_1_28 vss 3.13114e-17
C7932 a_1_30 vss 3.13114e-17
C7933 a_1_29 vss 3.13114e-17
C7934 a_1_31 vss 3.13114e-17
C7935 a_1_30 vss 3.13114e-17
C7936 a_1_32 vss 3.13114e-17
C7937 a_1_31 vss 3.13114e-17
C7938 a_1_33 vss 3.13114e-17
C7939 a_1_32 vss 3.13114e-17
C7940 a_1_34 vss 3.13114e-17
C7941 a_1_33 vss 3.13114e-17
C7942 a_1_35 vss 3.13114e-17
C7943 a_1_34 vss 3.13114e-17
C7944 a_1_36 vss 3.13114e-17
C7945 a_1_35 vss 3.13114e-17
C7946 a_1_37 vss 3.13114e-17
C7947 a_1_36 vss 3.13114e-17
C7948 a_1_38 vss 3.13114e-17
C7949 a_1_37 vss 3.13114e-17
C7950 a_1_39 vss 3.13114e-17
C7951 a_1_38 vss 3.13114e-17
C7952 a_1_40 vss 3.13114e-17
C7953 a_1_39 vss 3.13114e-17
C7954 a_1_41 vss 3.13114e-17
C7955 a_1_40 vss 3.13114e-17
C7956 a_1_42 vss 3.13114e-17
C7957 a_1_41 vss 3.13114e-17
C7958 a_1_43 vss 2.42663e-16
C7959 a_1_42 vss 2.42663e-16
C7960 a_1_44 vss 3.13114e-17
C7961 a_1_43 vss 3.13114e-17
C7962 a_1_45 vss 3.13114e-17
C7963 a_1_44 vss 3.13114e-17
C7964 a_1_46 vss 3.13114e-17
C7965 a_1_45 vss 3.13114e-17
C7966 a_1_47 vss 3.13114e-17
C7967 a_1_46 vss 3.13114e-17
C7968 a_1_48 vss 3.13114e-17
C7969 a_1_47 vss 3.13114e-17
C7970 a_1_49 vss 3.13114e-17
C7971 a_1_48 vss 3.13114e-17
C7972 a_1_50 vss 3.13114e-17
C7973 a_1_49 vss 3.13114e-17
C7974 a_1_81 vss 1.40901e-16
C7975 a_1_50 vss 1.40901e-16
C7976 a_1_52 vss 1.40901e-17
C7977 a_1_51 vss 1.40901e-17
C7978 a_1_53 vss 3.13114e-17
C7979 a_1_52 vss 3.13114e-17
C7980 a_1_54 vss 3.13114e-17
C7981 a_1_53 vss 3.13114e-17
C7982 a_1_55 vss 3.13114e-17
C7983 a_1_54 vss 3.13114e-17
C7984 a_1_56 vss 3.13114e-17
C7985 a_1_55 vss 3.13114e-17
C7986 a_1_57 vss 3.13114e-17
C7987 a_1_56 vss 3.13114e-17
C7988 a_1_58 vss 3.13114e-17
C7989 a_1_57 vss 3.13114e-17
C7990 a_1_59 vss 3.13114e-17
C7991 a_1_58 vss 3.13114e-17
C7992 a_1_60 vss 3.13114e-17
C7993 a_1_59 vss 3.13114e-17
C7994 a_1_61 vss 3.13114e-17
C7995 a_1_60 vss 3.13114e-17
C7996 a_1_62 vss 3.13114e-17
C7997 a_1_61 vss 3.13114e-17
C7998 a_1_63 vss 3.13114e-17
C7999 a_1_62 vss 3.13114e-17
C8000 a_1_64 vss 3.13114e-17
C8001 a_1_63 vss 3.13114e-17
C8002 a_1_65 vss 3.13114e-17
C8003 a_1_64 vss 3.13114e-17
C8004 a_1_66 vss 3.13114e-17
C8005 a_1_65 vss 3.13114e-17
C8006 a_1_67 vss 3.13114e-17
C8007 a_1_66 vss 3.13114e-17
C8008 a_1_68 vss 3.13114e-17
C8009 a_1_67 vss 3.13114e-17
C8010 a_1_69 vss 3.13114e-17
C8011 a_1_68 vss 3.13114e-17
C8012 a_1_70 vss 3.13114e-17
C8013 a_1_69 vss 3.13114e-17
C8014 a_1_71 vss 3.13114e-17
C8015 a_1_70 vss 3.13114e-17
C8016 a_1_72 vss 2.42663e-16
C8017 a_1_71 vss 2.42663e-16
C8018 a_1_73 vss 3.13114e-17
C8019 a_1_72 vss 3.13114e-17
C8020 a_1_74 vss 3.13114e-17
C8021 a_1_73 vss 3.13114e-17
C8022 a_1_75 vss 3.13114e-17
C8023 a_1_74 vss 3.13114e-17
C8024 a_1_76 vss 3.13114e-17
C8025 a_1_75 vss 3.13114e-17
C8026 a_1_77 vss 3.13114e-17
C8027 a_1_76 vss 3.13114e-17
C8028 a_1_78 vss 3.13114e-17
C8029 a_1_77 vss 3.13114e-17
C8030 a_1_79 vss 3.13114e-17
C8031 a_1_78 vss 3.13114e-17
C8032 a_1_82 vss 1.40901e-16
C8033 a_1_79 vss 1.40901e-16
C8034 a_1_82 vss 6.34418e-17
C8035 a_1_80 vss 6.34418e-17
C8036 a_1_81 vss 1.42197e-16
C8037 a_1_82 vss 1.42197e-16
C8038 a_1_83 vss 6.8969e-16
C8039 a_1_82 vss 6.8969e-16
C8040 a_1_84 vss 3.48676e-17
C8041 a_1_83 vss 3.48676e-17
C8042 a_1 vss 4.3846e-15
C8043 a_1_84 vss 4.3846e-15

R156_1 n5334 n5334_26 0.001
R156_2 n5334 n5334_27 0.001
R156_3 n5334 n5334_28 0.001
R156_4 n5334 n5334_25 0.001
R156_5 n5334 n5334_23 0.001
R156_6 n5334 n5334_22 0.001
R156_7 n5334 n5334_24 0.001
R156_8 n5334_20 n5334_2 0.001
R156_9 n5334_16 n5334_2 0.001
R156_10 n5334_17 n5334_2 0.001
R156_11 n5334_18 n5334_2 0.001
R156_12 n5334_19 n5334_2 0.001
R156_13 n5334_14 n5334_2 0.001
R156_14 n5334_13 n5334_2 0.001
R156_15 n5334_15 n5334_2 0.001
R156_16 n5334_11 n5334_2 0.001
R156_17 n5334_10 n5334_2 0.001
R156_18 n5334_12 n5334_2 0.001
R156_19 n5334_9 n5334_2 0.001
R156_20 n5334_7 n5334_2 0.001
R156_21 n5334_8 n5334_2 0.001
R156_22 n5334_6 n5334_2 0.001
R156_23 n5334_21 n5334_5 0.001
R156_24 n5334_3 n5334_4 453.6
R156_25 n5334_5 n5334_4 14.4
R156_26 n5334_7 n5334_6 0.108
R156_27 n5334_8 n5334_7 0.108
R156_28 n5334_9 n5334_8 0.108
R156_29 n5334_10 n5334_9 0.108
R156_30 n5334_11 n5334_10 0.108
R156_31 n5334_12 n5334_11 0.108
R156_32 n5334_13 n5334_12 0.108
R156_33 n5334_14 n5334_13 0.108
R156_34 n5334_15 n5334_14 0.108
R156_35 n5334_16 n5334_15 0.108
R156_36 n5334_17 n5334_16 0.108
R156_37 n5334_18 n5334_17 0.108
R156_38 n5334_19 n5334_18 0.108
R156_39 n5334_20 n5334_19 0.108
R156_40 n5334_21 n5334_20 0.108
R156_41 n5334_22 n5334_21 0.756
R156_42 n5334_23 n5334_22 0.108
R156_43 n5334_24 n5334_23 0.108
R156_44 n5334_25 n5334_24 0.108
R156_45 n5334_26 n5334_25 0.108
R156_46 n5334_27 n5334_26 0.108
R156_47 n5334_28 n5334_27 0.108

C8044 n5334_3 vss 4.98819e-16
C8045 n5334_4 vss 4.98819e-16
C8046 n5334_5 vss 8.41104e-17
C8047 n5334_4 vss 8.41104e-17
C8048 n5334_7 vss 2.92378e-17
C8049 n5334_6 vss 2.92378e-17
C8050 n5334_8 vss 2.92378e-17
C8051 n5334_7 vss 2.92378e-17
C8052 n5334_9 vss 2.92378e-17
C8053 n5334_8 vss 2.92378e-17
C8054 n5334_10 vss 2.92378e-17
C8055 n5334_9 vss 2.92378e-17
C8056 n5334_11 vss 2.92378e-17
C8057 n5334_10 vss 2.92378e-17
C8058 n5334_12 vss 2.92378e-17
C8059 n5334_11 vss 2.92378e-17
C8060 n5334_13 vss 2.92378e-17
C8061 n5334_12 vss 2.92378e-17
C8062 n5334_14 vss 2.92378e-17
C8063 n5334_13 vss 2.92378e-17
C8064 n5334_15 vss 2.92378e-17
C8065 n5334_14 vss 2.92378e-17
C8066 n5334_16 vss 2.92378e-17
C8067 n5334_15 vss 2.92378e-17
C8068 n5334_17 vss 2.92378e-17
C8069 n5334_16 vss 2.92378e-17
C8070 n5334_18 vss 2.92378e-17
C8071 n5334_17 vss 2.92378e-17
C8072 n5334_19 vss 2.92378e-17
C8073 n5334_18 vss 2.92378e-17
C8074 n5334_20 vss 2.92378e-17
C8075 n5334_19 vss 2.92378e-17
C8076 n5334_21 vss 3.65472e-17
C8077 n5334_20 vss 3.65472e-17
C8078 n5334_22 vss 1.46189e-16
C8079 n5334_21 vss 1.46189e-16
C8080 n5334_23 vss 2.92378e-17
C8081 n5334_22 vss 2.92378e-17
C8082 n5334_24 vss 2.92378e-17
C8083 n5334_23 vss 2.92378e-17
C8084 n5334_25 vss 2.92378e-17
C8085 n5334_24 vss 2.92378e-17
C8086 n5334_26 vss 2.92378e-17
C8087 n5334_25 vss 2.92378e-17
C8088 n5334_27 vss 2.92378e-17
C8089 n5334_26 vss 2.92378e-17
C8090 n5334_28 vss 2.92378e-17
C8091 n5334_27 vss 2.92378e-17

R157_1 n5373 n5373_35 0.001
R157_2 n5373 n5373_36 0.001
R157_3 n5373 n5373_37 0.001
R157_4 n5373 n5373_33 0.001
R157_5 n5373 n5373_34 0.001
R157_6 n5373 n5373_32 0.001
R157_7 n5373 n5373_31 0.001
R157_8 n5373_29 n5373_2 0.001
R157_9 n5373_25 n5373_2 0.001
R157_10 n5373_26 n5373_2 0.001
R157_11 n5373_27 n5373_2 0.001
R157_12 n5373_28 n5373_2 0.001
R157_13 n5373_22 n5373_2 0.001
R157_14 n5373_23 n5373_2 0.001
R157_15 n5373_24 n5373_2 0.001
R157_16 n5373_21 n5373_2 0.001
R157_17 n5373_19 n5373_2 0.001
R157_18 n5373_20 n5373_2 0.001
R157_19 n5373_18 n5373_2 0.001
R157_20 n5373_17 n5373_2 0.001
R157_21 n5373_16 n5373_2 0.001
R157_22 n5373_15 n5373_2 0.001
R157_23 n5373_14 n5373_12 0.001
R157_24 n5373_4 n5373_3 43.2
R157_25 n5373_11 n5373_4 21.6
R157_26 n5373_5 n5373_11 21.6
R157_27 n5373_6 n5373_5 43.2
R157_28 n5373_8 n5373_7 43.2
R157_29 n5373_13 n5373_8 21.6
R157_30 n5373_9 n5373_13 21.6
R157_31 n5373_10 n5373_9 43.2
R157_32 n5373_12 n5373_11 28.8
R157_33 n5373_13 n5373_12 28.8
R157_34 n5373_30 n5373_14 0.648
R157_35 n5373_16 n5373_15 0.108
R157_36 n5373_17 n5373_16 0.108
R157_37 n5373_18 n5373_17 0.108
R157_38 n5373_19 n5373_18 0.108
R157_39 n5373_20 n5373_19 0.108
R157_40 n5373_21 n5373_20 0.108
R157_41 n5373_22 n5373_21 0.108
R157_42 n5373_23 n5373_22 0.108
R157_43 n5373_24 n5373_23 0.108
R157_44 n5373_25 n5373_24 0.108
R157_45 n5373_26 n5373_25 0.108
R157_46 n5373_27 n5373_26 0.108
R157_47 n5373_28 n5373_27 0.108
R157_48 n5373_29 n5373_28 0.108
R157_49 n5373_30 n5373_29 0.432
R157_50 n5373_31 n5373_30 0.54
R157_51 n5373_32 n5373_31 0.108
R157_52 n5373_33 n5373_32 0.108
R157_53 n5373_34 n5373_33 0.108
R157_54 n5373_35 n5373_34 0.108
R157_55 n5373_36 n5373_35 0.108
R157_56 n5373_37 n5373_36 0.108

C8092 n5373_4 vss 4.69476e-17
C8093 n5373_3 vss 4.69476e-17
C8094 n5373_11 vss 2.34738e-17
C8095 n5373_4 vss 2.34738e-17
C8096 n5373_5 vss 2.34738e-17
C8097 n5373_11 vss 2.34738e-17
C8098 n5373_6 vss 4.69476e-17
C8099 n5373_5 vss 4.69476e-17
C8100 n5373_8 vss 4.69476e-17
C8101 n5373_7 vss 4.69476e-17
C8102 n5373_13 vss 2.34738e-17
C8103 n5373_8 vss 2.34738e-17
C8104 n5373_9 vss 2.34738e-17
C8105 n5373_13 vss 2.34738e-17
C8106 n5373_10 vss 4.69476e-17
C8107 n5373_9 vss 4.69476e-17
C8108 n5373_12 vss 7.33536e-17
C8109 n5373_11 vss 7.33536e-17
C8110 n5373_13 vss 8.25228e-17
C8111 n5373_12 vss 8.25228e-17
C8112 n5373_30 vss 1.3157e-16
C8113 n5373_14 vss 1.3157e-16
C8114 n5373_16 vss 2.92378e-17
C8115 n5373_15 vss 2.92378e-17
C8116 n5373_17 vss 2.92378e-17
C8117 n5373_16 vss 2.92378e-17
C8118 n5373_18 vss 2.92378e-17
C8119 n5373_17 vss 2.92378e-17
C8120 n5373_19 vss 2.92378e-17
C8121 n5373_18 vss 2.92378e-17
C8122 n5373_20 vss 2.92378e-17
C8123 n5373_19 vss 2.92378e-17
C8124 n5373_21 vss 2.92378e-17
C8125 n5373_20 vss 2.92378e-17
C8126 n5373_22 vss 2.92378e-17
C8127 n5373_21 vss 2.92378e-17
C8128 n5373_23 vss 2.92378e-17
C8129 n5373_22 vss 2.92378e-17
C8130 n5373_24 vss 2.92378e-17
C8131 n5373_23 vss 2.92378e-17
C8132 n5373_25 vss 2.92378e-17
C8133 n5373_24 vss 2.92378e-17
C8134 n5373_26 vss 2.92378e-17
C8135 n5373_25 vss 2.92378e-17
C8136 n5373_27 vss 2.92378e-17
C8137 n5373_26 vss 2.92378e-17
C8138 n5373_28 vss 2.92378e-17
C8139 n5373_27 vss 2.92378e-17
C8140 n5373_29 vss 2.92378e-17
C8141 n5373_28 vss 2.92378e-17
C8142 n5373_30 vss 8.77133e-17
C8143 n5373_29 vss 8.77133e-17
C8144 n5373_31 vss 9.50227e-17
C8145 n5373_30 vss 9.50227e-17
C8146 n5373_32 vss 2.92378e-17
C8147 n5373_31 vss 2.92378e-17
C8148 n5373_33 vss 2.92378e-17
C8149 n5373_32 vss 2.92378e-17
C8150 n5373_34 vss 2.92378e-17
C8151 n5373_33 vss 2.92378e-17
C8152 n5373_35 vss 2.92378e-17
C8153 n5373_34 vss 2.92378e-17
C8154 n5373_36 vss 2.92378e-17
C8155 n5373_35 vss 2.92378e-17
C8156 n5373_37 vss 2.92378e-17
C8157 n5373_36 vss 2.92378e-17

R158_1 s_2_82 s_2_1 0.001
R158_2 s_2_83 s_2_1 0.001
R158_3 s_2_81 s_2_1 0.001
R158_4 s_2_80 s_2_1 0.001
R158_5 s_2_78 s_2_1 0.001
R158_6 s_2_79 s_2_1 0.001
R158_7 s_2_77 s_2_1 0.001
R158_8 s_2_75 s_2_1 0.001
R158_9 s_2_76 s_2_1 0.001
R158_10 s_2_74 s_2_1 0.001
R158_11 s_2_73 s_2_1 0.001
R158_12 s_2_72 s_2_1 0.001
R158_13 s_2_71 s_2_1 0.001
R158_14 s_2_70 s_2_1 0.001
R158_15 s_2_69 s_2_1 0.001
R158_16 s_2_68 s_2_1 0.001
R158_17 s_2_67 s_2_1 0.001
R158_18 s_2_66 s_2_1 0.001
R158_19 s_2_64 s_2_1 0.001
R158_20 s_2_65 s_2_1 0.001
R158_21 s_2_62 s_2_2 0.001
R158_22 s_2_63 s_2_2 0.001
R158_23 s_2_61 s_2_2 0.001
R158_24 s_2_60 s_2_2 0.001
R158_25 s_2_59 s_2_2 0.001
R158_26 s_2_58 s_2_2 0.001
R158_27 s_2_57 s_2_2 0.001
R158_28 s_2_56 s_2_2 0.001
R158_29 s_2_54 s_2_3 0.001
R158_30 s_2_53 s_2_3 0.001
R158_31 s_2_52 s_2_3 0.001
R158_32 s_2_51 s_2_3 0.001
R158_33 s_2_49 s_2_3 0.001
R158_34 s_2_50 s_2_3 0.001
R158_35 s_2_48 s_2_3 0.001
R158_36 s_2_46 s_2_3 0.001
R158_37 s_2_47 s_2_3 0.001
R158_38 s_2_45 s_2_3 0.001
R158_39 s_2_44 s_2_3 0.001
R158_40 s_2_43 s_2_3 0.001
R158_41 s_2_42 s_2_3 0.001
R158_42 s_2_41 s_2_3 0.001
R158_43 s_2_40 s_2_3 0.001
R158_44 s_2_39 s_2_3 0.001
R158_45 s_2_38 s_2_3 0.001
R158_46 s_2_37 s_2_3 0.001
R158_47 s_2_36 s_2_3 0.001
R158_48 s_2_35 s_2_3 0.001
R158_49 s_2_33 s_2_4 0.001
R158_50 s_2_34 s_2_4 0.001
R158_51 s_2_32 s_2_4 0.001
R158_52 s_2_31 s_2_4 0.001
R158_53 s_2_30 s_2_4 0.001
R158_54 s_2_29 s_2_4 0.001
R158_55 s_2_28 s_2_4 0.001
R158_56 s_2_27 s_2_4 0.001
R158_57 s_2_5 s_2_379 0.001
R158_58 s_2_5 s_2_380 0.001
R158_59 s_2_5 s_2_378 0.001
R158_60 s_2_5 s_2_377 0.001
R158_61 s_2_5 s_2_375 0.001
R158_62 s_2_5 s_2_376 0.001
R158_63 s_2_5 s_2_374 0.001
R158_64 s_2_5 s_2_372 0.001
R158_65 s_2_5 s_2_373 0.001
R158_66 s_2_5 s_2_371 0.001
R158_67 s_2_5 s_2_370 0.001
R158_68 s_2_5 s_2_369 0.001
R158_69 s_2_5 s_2_368 0.001
R158_70 s_2_5 s_2_367 0.001
R158_71 s_2_5 s_2_366 0.001
R158_72 s_2_5 s_2_365 0.001
R158_73 s_2_5 s_2_364 0.001
R158_74 s_2_5 s_2_363 0.001
R158_75 s_2_5 s_2_361 0.001
R158_76 s_2_5 s_2_362 0.001
R158_77 s_2_360 s_2_6 0.001
R158_78 s_2_359 s_2_6 0.001
R158_79 s_2_358 s_2_6 0.001
R158_80 s_2_357 s_2_6 0.001
R158_81 s_2_356 s_2_6 0.001
R158_82 s_2_355 s_2_6 0.001
R158_83 s_2_354 s_2_6 0.001
R158_84 s_2_353 s_2_6 0.001
R158_85 s_2_141 s_2_7 0.001
R158_86 s_2_140 s_2_7 0.001
R158_87 s_2_139 s_2_7 0.001
R158_88 s_2_138 s_2_7 0.001
R158_89 s_2_136 s_2_7 0.001
R158_90 s_2_137 s_2_7 0.001
R158_91 s_2_135 s_2_7 0.001
R158_92 s_2_133 s_2_7 0.001
R158_93 s_2_134 s_2_7 0.001
R158_94 s_2_132 s_2_7 0.001
R158_95 s_2_131 s_2_7 0.001
R158_96 s_2_130 s_2_7 0.001
R158_97 s_2_129 s_2_7 0.001
R158_98 s_2_128 s_2_7 0.001
R158_99 s_2_127 s_2_7 0.001
R158_100 s_2_126 s_2_7 0.001
R158_101 s_2_125 s_2_7 0.001
R158_102 s_2_124 s_2_7 0.001
R158_103 s_2_122 s_2_7 0.001
R158_104 s_2_123 s_2_7 0.001
R158_105 s_2_120 s_2_8 0.001
R158_106 s_2_121 s_2_8 0.001
R158_107 s_2_119 s_2_8 0.001
R158_108 s_2_118 s_2_8 0.001
R158_109 s_2_117 s_2_8 0.001
R158_110 s_2_116 s_2_8 0.001
R158_111 s_2_115 s_2_8 0.001
R158_112 s_2_114 s_2_8 0.001
R158_113 s_2_112 s_2_9 0.001
R158_114 s_2_111 s_2_9 0.001
R158_115 s_2_110 s_2_9 0.001
R158_116 s_2_109 s_2_9 0.001
R158_117 s_2_107 s_2_9 0.001
R158_118 s_2_108 s_2_9 0.001
R158_119 s_2_106 s_2_9 0.001
R158_120 s_2_105 s_2_9 0.001
R158_121 s_2_104 s_2_9 0.001
R158_122 s_2_103 s_2_9 0.001
R158_123 s_2_102 s_2_9 0.001
R158_124 s_2_101 s_2_9 0.001
R158_125 s_2_100 s_2_9 0.001
R158_126 s_2_99 s_2_9 0.001
R158_127 s_2_98 s_2_9 0.001
R158_128 s_2_97 s_2_9 0.001
R158_129 s_2_96 s_2_9 0.001
R158_130 s_2_95 s_2_9 0.001
R158_131 s_2_94 s_2_9 0.001
R158_132 s_2_93 s_2_9 0.001
R158_133 s_2_92 s_2_10 0.001
R158_134 s_2_91 s_2_10 0.001
R158_135 s_2_90 s_2_10 0.001
R158_136 s_2_89 s_2_10 0.001
R158_137 s_2_88 s_2_10 0.001
R158_138 s_2_87 s_2_10 0.001
R158_139 s_2_86 s_2_10 0.001
R158_140 s_2_85 s_2_10 0.001
R158_141 s_2_228 s_2_11 0.001
R158_142 s_2_227 s_2_11 0.001
R158_143 s_2_226 s_2_11 0.001
R158_144 s_2_225 s_2_11 0.001
R158_145 s_2_223 s_2_11 0.001
R158_146 s_2_224 s_2_11 0.001
R158_147 s_2_222 s_2_11 0.001
R158_148 s_2_220 s_2_11 0.001
R158_149 s_2_221 s_2_11 0.001
R158_150 s_2_219 s_2_11 0.001
R158_151 s_2_218 s_2_11 0.001
R158_152 s_2_217 s_2_11 0.001
R158_153 s_2_216 s_2_11 0.001
R158_154 s_2_215 s_2_11 0.001
R158_155 s_2_214 s_2_11 0.001
R158_156 s_2_213 s_2_11 0.001
R158_157 s_2_212 s_2_11 0.001
R158_158 s_2_211 s_2_11 0.001
R158_159 s_2_210 s_2_11 0.001
R158_160 s_2_209 s_2_11 0.001
R158_161 s_2_207 s_2_12 0.001
R158_162 s_2_208 s_2_12 0.001
R158_163 s_2_206 s_2_12 0.001
R158_164 s_2_205 s_2_12 0.001
R158_165 s_2_204 s_2_12 0.001
R158_166 s_2_203 s_2_12 0.001
R158_167 s_2_202 s_2_12 0.001
R158_168 s_2_201 s_2_12 0.001
R158_169 s_2_198 s_2_13 0.001
R158_170 s_2_199 s_2_13 0.001
R158_171 s_2_197 s_2_13 0.001
R158_172 s_2_196 s_2_13 0.001
R158_173 s_2_194 s_2_13 0.001
R158_174 s_2_195 s_2_13 0.001
R158_175 s_2_193 s_2_13 0.001
R158_176 s_2_191 s_2_13 0.001
R158_177 s_2_192 s_2_13 0.001
R158_178 s_2_190 s_2_13 0.001
R158_179 s_2_189 s_2_13 0.001
R158_180 s_2_188 s_2_13 0.001
R158_181 s_2_187 s_2_13 0.001
R158_182 s_2_186 s_2_13 0.001
R158_183 s_2_185 s_2_13 0.001
R158_184 s_2_184 s_2_13 0.001
R158_185 s_2_183 s_2_13 0.001
R158_186 s_2_182 s_2_13 0.001
R158_187 s_2_180 s_2_13 0.001
R158_188 s_2_181 s_2_13 0.001
R158_189 s_2_179 s_2_14 0.001
R158_190 s_2_178 s_2_14 0.001
R158_191 s_2_177 s_2_14 0.001
R158_192 s_2_176 s_2_14 0.001
R158_193 s_2_175 s_2_14 0.001
R158_194 s_2_174 s_2_14 0.001
R158_195 s_2_173 s_2_14 0.001
R158_196 s_2_172 s_2_14 0.001
R158_197 s_2_170 s_2_15 0.001
R158_198 s_2_169 s_2_15 0.001
R158_199 s_2_168 s_2_15 0.001
R158_200 s_2_167 s_2_15 0.001
R158_201 s_2_165 s_2_15 0.001
R158_202 s_2_166 s_2_15 0.001
R158_203 s_2_164 s_2_15 0.001
R158_204 s_2_162 s_2_15 0.001
R158_205 s_2_163 s_2_15 0.001
R158_206 s_2_161 s_2_15 0.001
R158_207 s_2_160 s_2_15 0.001
R158_208 s_2_158 s_2_15 0.001
R158_209 s_2_159 s_2_15 0.001
R158_210 s_2_157 s_2_15 0.001
R158_211 s_2_156 s_2_15 0.001
R158_212 s_2_155 s_2_15 0.001
R158_213 s_2_154 s_2_15 0.001
R158_214 s_2_153 s_2_15 0.001
R158_215 s_2_152 s_2_15 0.001
R158_216 s_2_151 s_2_15 0.001
R158_217 s_2_149 s_2_16 0.001
R158_218 s_2_150 s_2_16 0.001
R158_219 s_2_148 s_2_16 0.001
R158_220 s_2_147 s_2_16 0.001
R158_221 s_2_146 s_2_16 0.001
R158_222 s_2_145 s_2_16 0.001
R158_223 s_2_144 s_2_16 0.001
R158_224 s_2_143 s_2_16 0.001
R158_225 s_2_285 s_2_17 0.001
R158_226 s_2_286 s_2_17 0.001
R158_227 s_2_284 s_2_17 0.001
R158_228 s_2_283 s_2_17 0.001
R158_229 s_2_281 s_2_17 0.001
R158_230 s_2_282 s_2_17 0.001
R158_231 s_2_280 s_2_17 0.001
R158_232 s_2_278 s_2_17 0.001
R158_233 s_2_279 s_2_17 0.001
R158_234 s_2_277 s_2_17 0.001
R158_235 s_2_276 s_2_17 0.001
R158_236 s_2_275 s_2_17 0.001
R158_237 s_2_274 s_2_17 0.001
R158_238 s_2_273 s_2_17 0.001
R158_239 s_2_272 s_2_17 0.001
R158_240 s_2_271 s_2_17 0.001
R158_241 s_2_270 s_2_17 0.001
R158_242 s_2_269 s_2_17 0.001
R158_243 s_2_267 s_2_17 0.001
R158_244 s_2_268 s_2_17 0.001
R158_245 s_2_266 s_2_18 0.001
R158_246 s_2_265 s_2_18 0.001
R158_247 s_2_264 s_2_18 0.001
R158_248 s_2_263 s_2_18 0.001
R158_249 s_2_262 s_2_18 0.001
R158_250 s_2_261 s_2_18 0.001
R158_251 s_2_260 s_2_18 0.001
R158_252 s_2_259 s_2_18 0.001
R158_253 s_2_256 s_2_19 0.001
R158_254 s_2_257 s_2_19 0.001
R158_255 s_2_255 s_2_19 0.001
R158_256 s_2_254 s_2_19 0.001
R158_257 s_2_252 s_2_19 0.001
R158_258 s_2_253 s_2_19 0.001
R158_259 s_2_251 s_2_19 0.001
R158_260 s_2_249 s_2_19 0.001
R158_261 s_2_250 s_2_19 0.001
R158_262 s_2_248 s_2_19 0.001
R158_263 s_2_247 s_2_19 0.001
R158_264 s_2_245 s_2_19 0.001
R158_265 s_2_246 s_2_19 0.001
R158_266 s_2_244 s_2_19 0.001
R158_267 s_2_243 s_2_19 0.001
R158_268 s_2_242 s_2_19 0.001
R158_269 s_2_241 s_2_19 0.001
R158_270 s_2_240 s_2_19 0.001
R158_271 s_2_239 s_2_19 0.001
R158_272 s_2_238 s_2_19 0.001
R158_273 s_2_236 s_2_20 0.001
R158_274 s_2_237 s_2_20 0.001
R158_275 s_2_235 s_2_20 0.001
R158_276 s_2_234 s_2_20 0.001
R158_277 s_2_233 s_2_20 0.001
R158_278 s_2_232 s_2_20 0.001
R158_279 s_2_231 s_2_20 0.001
R158_280 s_2_230 s_2_20 0.001
R158_281 s_2_344 s_2_21 0.001
R158_282 s_2_343 s_2_21 0.001
R158_283 s_2_342 s_2_21 0.001
R158_284 s_2_341 s_2_21 0.001
R158_285 s_2_339 s_2_21 0.001
R158_286 s_2_340 s_2_21 0.001
R158_287 s_2_338 s_2_21 0.001
R158_288 s_2_336 s_2_21 0.001
R158_289 s_2_337 s_2_21 0.001
R158_290 s_2_335 s_2_21 0.001
R158_291 s_2_334 s_2_21 0.001
R158_292 s_2_333 s_2_21 0.001
R158_293 s_2_332 s_2_21 0.001
R158_294 s_2_331 s_2_21 0.001
R158_295 s_2_330 s_2_21 0.001
R158_296 s_2_329 s_2_21 0.001
R158_297 s_2_328 s_2_21 0.001
R158_298 s_2_327 s_2_21 0.001
R158_299 s_2_325 s_2_21 0.001
R158_300 s_2_326 s_2_21 0.001
R158_301 s_2_324 s_2_22 0.001
R158_302 s_2_323 s_2_22 0.001
R158_303 s_2_322 s_2_22 0.001
R158_304 s_2_321 s_2_22 0.001
R158_305 s_2_320 s_2_22 0.001
R158_306 s_2_319 s_2_22 0.001
R158_307 s_2_318 s_2_22 0.001
R158_308 s_2_317 s_2_22 0.001
R158_309 s_2 s_2_23 0.001
R158_310 s_2_315 s_2_24 0.001
R158_311 s_2_314 s_2_24 0.001
R158_312 s_2_313 s_2_24 0.001
R158_313 s_2_312 s_2_24 0.001
R158_314 s_2_310 s_2_24 0.001
R158_315 s_2_311 s_2_24 0.001
R158_316 s_2_309 s_2_24 0.001
R158_317 s_2_307 s_2_24 0.001
R158_318 s_2_308 s_2_24 0.001
R158_319 s_2_306 s_2_24 0.001
R158_320 s_2_305 s_2_24 0.001
R158_321 s_2_304 s_2_24 0.001
R158_322 s_2_303 s_2_24 0.001
R158_323 s_2_302 s_2_24 0.001
R158_324 s_2_301 s_2_24 0.001
R158_325 s_2_300 s_2_24 0.001
R158_326 s_2_299 s_2_24 0.001
R158_327 s_2_298 s_2_24 0.001
R158_328 s_2_297 s_2_24 0.001
R158_329 s_2_296 s_2_24 0.001
R158_330 s_2_294 s_2_25 0.001
R158_331 s_2_295 s_2_25 0.001
R158_332 s_2_293 s_2_25 0.001
R158_333 s_2_292 s_2_25 0.001
R158_334 s_2_291 s_2_25 0.001
R158_335 s_2_290 s_2_25 0.001
R158_336 s_2_289 s_2_25 0.001
R158_337 s_2_288 s_2_25 0.001
R158_338 s_2_352 s_2 0.108
R158_339 s_2_27 s_2_349 0.54
R158_340 s_2_28 s_2_27 0.108
R158_341 s_2_29 s_2_28 0.108
R158_342 s_2_30 s_2_29 0.108
R158_343 s_2_31 s_2_30 0.108
R158_344 s_2_32 s_2_31 0.108
R158_345 s_2_33 s_2_32 0.108
R158_346 s_2_34 s_2_33 0.108
R158_347 s_2_35 s_2_34 0.864
R158_348 s_2_36 s_2_35 0.108
R158_349 s_2_37 s_2_36 0.108
R158_350 s_2_38 s_2_37 0.108
R158_351 s_2_39 s_2_38 0.108
R158_352 s_2_40 s_2_39 0.108
R158_353 s_2_41 s_2_40 0.108
R158_354 s_2_42 s_2_41 0.108
R158_355 s_2_43 s_2_42 0.108
R158_356 s_2_44 s_2_43 0.108
R158_357 s_2_45 s_2_44 0.108
R158_358 s_2_46 s_2_45 0.108
R158_359 s_2_47 s_2_46 0.108
R158_360 s_2_48 s_2_47 0.108
R158_361 s_2_49 s_2_48 0.108
R158_362 s_2_50 s_2_49 0.108
R158_363 s_2_51 s_2_50 0.108
R158_364 s_2_52 s_2_51 0.108
R158_365 s_2_53 s_2_52 0.108
R158_366 s_2_54 s_2_53 0.108
R158_367 s_2_55 s_2_54 0.001
R158_368 s_2_56 s_2_351 0.54
R158_369 s_2_57 s_2_56 0.108
R158_370 s_2_58 s_2_57 0.108
R158_371 s_2_59 s_2_58 0.108
R158_372 s_2_60 s_2_59 0.108
R158_373 s_2_61 s_2_60 0.108
R158_374 s_2_62 s_2_61 0.108
R158_375 s_2_63 s_2_62 0.108
R158_376 s_2_64 s_2_63 0.864
R158_377 s_2_65 s_2_64 0.108
R158_378 s_2_66 s_2_65 0.108
R158_379 s_2_67 s_2_66 0.108
R158_380 s_2_68 s_2_67 0.108
R158_381 s_2_69 s_2_68 0.108
R158_382 s_2_70 s_2_69 0.108
R158_383 s_2_71 s_2_70 0.108
R158_384 s_2_72 s_2_71 0.108
R158_385 s_2_73 s_2_72 0.108
R158_386 s_2_74 s_2_73 0.108
R158_387 s_2_75 s_2_74 0.108
R158_388 s_2_76 s_2_75 0.108
R158_389 s_2_77 s_2_76 0.108
R158_390 s_2_78 s_2_77 0.108
R158_391 s_2_79 s_2_78 0.108
R158_392 s_2_80 s_2_79 0.108
R158_393 s_2_81 s_2_80 0.108
R158_394 s_2_82 s_2_81 0.108
R158_395 s_2_83 s_2_82 0.108
R158_396 s_2_84 s_2_83 0.001
R158_397 s_2_85 s_2_352 1.296
R158_398 s_2_86 s_2_85 0.108
R158_399 s_2_87 s_2_86 0.108
R158_400 s_2_88 s_2_87 0.108
R158_401 s_2_89 s_2_88 0.108
R158_402 s_2_90 s_2_89 0.108
R158_403 s_2_91 s_2_90 0.108
R158_404 s_2_92 s_2_91 0.108
R158_405 s_2_93 s_2_92 0.864
R158_406 s_2_94 s_2_93 0.108
R158_407 s_2_95 s_2_94 0.108
R158_408 s_2_96 s_2_95 0.108
R158_409 s_2_97 s_2_96 0.108
R158_410 s_2_98 s_2_97 0.108
R158_411 s_2_99 s_2_98 0.108
R158_412 s_2_100 s_2_99 0.108
R158_413 s_2_101 s_2_100 0.108
R158_414 s_2_102 s_2_101 0.108
R158_415 s_2_103 s_2_102 0.108
R158_416 s_2_104 s_2_103 0.108
R158_417 s_2_105 s_2_104 0.108
R158_418 s_2_106 s_2_105 0.108
R158_419 s_2_107 s_2_106 0.108
R158_420 s_2_108 s_2_107 0.108
R158_421 s_2_109 s_2_108 0.108
R158_422 s_2_110 s_2_109 0.108
R158_423 s_2_111 s_2_110 0.108
R158_424 s_2_112 s_2_111 0.108
R158_425 s_2_113 s_2_112 0.001
R158_426 s_2_114 s_2_352 1.296
R158_427 s_2_115 s_2_114 0.108
R158_428 s_2_116 s_2_115 0.108
R158_429 s_2_117 s_2_116 0.108
R158_430 s_2_118 s_2_117 0.108
R158_431 s_2_119 s_2_118 0.108
R158_432 s_2_120 s_2_119 0.108
R158_433 s_2_121 s_2_120 0.108
R158_434 s_2_122 s_2_121 0.864
R158_435 s_2_123 s_2_122 0.108
R158_436 s_2_124 s_2_123 0.108
R158_437 s_2_125 s_2_124 0.108
R158_438 s_2_126 s_2_125 0.108
R158_439 s_2_127 s_2_126 0.108
R158_440 s_2_128 s_2_127 0.108
R158_441 s_2_129 s_2_128 0.108
R158_442 s_2_130 s_2_129 0.108
R158_443 s_2_131 s_2_130 0.108
R158_444 s_2_132 s_2_131 0.108
R158_445 s_2_133 s_2_132 0.108
R158_446 s_2_134 s_2_133 0.108
R158_447 s_2_135 s_2_134 0.108
R158_448 s_2_136 s_2_135 0.108
R158_449 s_2_137 s_2_136 0.108
R158_450 s_2_138 s_2_137 0.108
R158_451 s_2_139 s_2_138 0.108
R158_452 s_2_140 s_2_139 0.108
R158_453 s_2_141 s_2_140 0.108
R158_454 s_2_142 s_2_141 0.001
R158_455 s_2_143 s_2_352 1.296
R158_456 s_2_144 s_2_143 0.108
R158_457 s_2_145 s_2_144 0.108
R158_458 s_2_146 s_2_145 0.108
R158_459 s_2_147 s_2_146 0.108
R158_460 s_2_148 s_2_147 0.108
R158_461 s_2_149 s_2_148 0.108
R158_462 s_2_150 s_2_149 0.108
R158_463 s_2_151 s_2_150 0.864
R158_464 s_2_152 s_2_151 0.108
R158_465 s_2_153 s_2_152 0.108
R158_466 s_2_154 s_2_153 0.108
R158_467 s_2_155 s_2_154 0.108
R158_468 s_2_156 s_2_155 0.108
R158_469 s_2_157 s_2_156 0.108
R158_470 s_2_158 s_2_157 0.108
R158_471 s_2_159 s_2_158 0.108
R158_472 s_2_160 s_2_159 0.108
R158_473 s_2_161 s_2_160 0.108
R158_474 s_2_162 s_2_161 0.108
R158_475 s_2_163 s_2_162 0.108
R158_476 s_2_164 s_2_163 0.108
R158_477 s_2_165 s_2_164 0.108
R158_478 s_2_166 s_2_165 0.108
R158_479 s_2_167 s_2_166 0.108
R158_480 s_2_168 s_2_167 0.108
R158_481 s_2_169 s_2_168 0.108
R158_482 s_2_170 s_2_169 0.108
R158_483 s_2_171 s_2_170 0.001
R158_484 s_2_172 s_2_352 1.296
R158_485 s_2_173 s_2_172 0.108
R158_486 s_2_174 s_2_173 0.108
R158_487 s_2_175 s_2_174 0.108
R158_488 s_2_176 s_2_175 0.108
R158_489 s_2_177 s_2_176 0.108
R158_490 s_2_178 s_2_177 0.108
R158_491 s_2_179 s_2_178 0.108
R158_492 s_2_180 s_2_179 0.864
R158_493 s_2_181 s_2_180 0.108
R158_494 s_2_182 s_2_181 0.108
R158_495 s_2_183 s_2_182 0.108
R158_496 s_2_184 s_2_183 0.108
R158_497 s_2_185 s_2_184 0.108
R158_498 s_2_186 s_2_185 0.108
R158_499 s_2_187 s_2_186 0.108
R158_500 s_2_188 s_2_187 0.108
R158_501 s_2_189 s_2_188 0.108
R158_502 s_2_190 s_2_189 0.108
R158_503 s_2_191 s_2_190 0.108
R158_504 s_2_192 s_2_191 0.108
R158_505 s_2_193 s_2_192 0.108
R158_506 s_2_194 s_2_193 0.108
R158_507 s_2_195 s_2_194 0.108
R158_508 s_2_196 s_2_195 0.108
R158_509 s_2_197 s_2_196 0.108
R158_510 s_2_198 s_2_197 0.108
R158_511 s_2_199 s_2_198 0.108
R158_512 s_2_200 s_2_199 0.001
R158_513 s_2_201 s_2_352 1.296
R158_514 s_2_202 s_2_201 0.108
R158_515 s_2_203 s_2_202 0.108
R158_516 s_2_204 s_2_203 0.108
R158_517 s_2_205 s_2_204 0.108
R158_518 s_2_206 s_2_205 0.108
R158_519 s_2_207 s_2_206 0.108
R158_520 s_2_208 s_2_207 0.108
R158_521 s_2_209 s_2_208 0.864
R158_522 s_2_210 s_2_209 0.108
R158_523 s_2_211 s_2_210 0.108
R158_524 s_2_212 s_2_211 0.108
R158_525 s_2_213 s_2_212 0.108
R158_526 s_2_214 s_2_213 0.108
R158_527 s_2_215 s_2_214 0.108
R158_528 s_2_216 s_2_215 0.108
R158_529 s_2_217 s_2_216 0.108
R158_530 s_2_218 s_2_217 0.108
R158_531 s_2_219 s_2_218 0.108
R158_532 s_2_220 s_2_219 0.108
R158_533 s_2_221 s_2_220 0.108
R158_534 s_2_222 s_2_221 0.108
R158_535 s_2_223 s_2_222 0.108
R158_536 s_2_224 s_2_223 0.108
R158_537 s_2_225 s_2_224 0.108
R158_538 s_2_226 s_2_225 0.108
R158_539 s_2_227 s_2_226 0.108
R158_540 s_2_228 s_2_227 0.108
R158_541 s_2_229 s_2_228 0.001
R158_542 s_2_230 s_2_352 1.296
R158_543 s_2_231 s_2_230 0.108
R158_544 s_2_232 s_2_231 0.108
R158_545 s_2_233 s_2_232 0.108
R158_546 s_2_234 s_2_233 0.108
R158_547 s_2_235 s_2_234 0.108
R158_548 s_2_236 s_2_235 0.108
R158_549 s_2_237 s_2_236 0.108
R158_550 s_2_238 s_2_237 0.864
R158_551 s_2_239 s_2_238 0.108
R158_552 s_2_240 s_2_239 0.108
R158_553 s_2_241 s_2_240 0.108
R158_554 s_2_242 s_2_241 0.108
R158_555 s_2_243 s_2_242 0.108
R158_556 s_2_244 s_2_243 0.108
R158_557 s_2_245 s_2_244 0.108
R158_558 s_2_246 s_2_245 0.108
R158_559 s_2_247 s_2_246 0.108
R158_560 s_2_248 s_2_247 0.108
R158_561 s_2_249 s_2_248 0.108
R158_562 s_2_250 s_2_249 0.108
R158_563 s_2_251 s_2_250 0.108
R158_564 s_2_252 s_2_251 0.108
R158_565 s_2_253 s_2_252 0.108
R158_566 s_2_254 s_2_253 0.108
R158_567 s_2_255 s_2_254 0.108
R158_568 s_2_256 s_2_255 0.108
R158_569 s_2_257 s_2_256 0.108
R158_570 s_2_258 s_2_257 0.001
R158_571 s_2_259 s_2_352 1.296
R158_572 s_2_260 s_2_259 0.108
R158_573 s_2_261 s_2_260 0.108
R158_574 s_2_262 s_2_261 0.108
R158_575 s_2_263 s_2_262 0.108
R158_576 s_2_264 s_2_263 0.108
R158_577 s_2_265 s_2_264 0.108
R158_578 s_2_266 s_2_265 0.108
R158_579 s_2_267 s_2_266 0.864
R158_580 s_2_268 s_2_267 0.108
R158_581 s_2_269 s_2_268 0.108
R158_582 s_2_270 s_2_269 0.108
R158_583 s_2_271 s_2_270 0.108
R158_584 s_2_272 s_2_271 0.108
R158_585 s_2_273 s_2_272 0.108
R158_586 s_2_274 s_2_273 0.108
R158_587 s_2_275 s_2_274 0.108
R158_588 s_2_276 s_2_275 0.108
R158_589 s_2_277 s_2_276 0.108
R158_590 s_2_278 s_2_277 0.108
R158_591 s_2_279 s_2_278 0.108
R158_592 s_2_280 s_2_279 0.108
R158_593 s_2_281 s_2_280 0.108
R158_594 s_2_282 s_2_281 0.108
R158_595 s_2_283 s_2_282 0.108
R158_596 s_2_284 s_2_283 0.108
R158_597 s_2_285 s_2_284 0.108
R158_598 s_2_286 s_2_285 0.108
R158_599 s_2_287 s_2_286 0.001
R158_600 s_2_288 s_2_346 0.54
R158_601 s_2_289 s_2_288 0.108
R158_602 s_2_290 s_2_289 0.108
R158_603 s_2_291 s_2_290 0.108
R158_604 s_2_292 s_2_291 0.108
R158_605 s_2_293 s_2_292 0.108
R158_606 s_2_294 s_2_293 0.108
R158_607 s_2_295 s_2_294 0.108
R158_608 s_2_296 s_2_295 0.864
R158_609 s_2_297 s_2_296 0.108
R158_610 s_2_298 s_2_297 0.108
R158_611 s_2_299 s_2_298 0.108
R158_612 s_2_300 s_2_299 0.108
R158_613 s_2_301 s_2_300 0.108
R158_614 s_2_302 s_2_301 0.108
R158_615 s_2_303 s_2_302 0.108
R158_616 s_2_304 s_2_303 0.108
R158_617 s_2_305 s_2_304 0.108
R158_618 s_2_306 s_2_305 0.108
R158_619 s_2_307 s_2_306 0.108
R158_620 s_2_308 s_2_307 0.108
R158_621 s_2_309 s_2_308 0.108
R158_622 s_2_310 s_2_309 0.108
R158_623 s_2_311 s_2_310 0.108
R158_624 s_2_312 s_2_311 0.108
R158_625 s_2_313 s_2_312 0.108
R158_626 s_2_314 s_2_313 0.108
R158_627 s_2_315 s_2_314 0.108
R158_628 s_2_316 s_2_315 0.001
R158_629 s_2_317 s_2_348 0.54
R158_630 s_2_318 s_2_317 0.108
R158_631 s_2_319 s_2_318 0.108
R158_632 s_2_320 s_2_319 0.108
R158_633 s_2_321 s_2_320 0.108
R158_634 s_2_322 s_2_321 0.108
R158_635 s_2_323 s_2_322 0.108
R158_636 s_2_324 s_2_323 0.108
R158_637 s_2_325 s_2_324 0.864
R158_638 s_2_326 s_2_325 0.108
R158_639 s_2_327 s_2_326 0.108
R158_640 s_2_328 s_2_327 0.108
R158_641 s_2_329 s_2_328 0.108
R158_642 s_2_330 s_2_329 0.108
R158_643 s_2_331 s_2_330 0.108
R158_644 s_2_332 s_2_331 0.108
R158_645 s_2_333 s_2_332 0.108
R158_646 s_2_334 s_2_333 0.108
R158_647 s_2_335 s_2_334 0.108
R158_648 s_2_336 s_2_335 0.108
R158_649 s_2_337 s_2_336 0.108
R158_650 s_2_338 s_2_337 0.108
R158_651 s_2_339 s_2_338 0.108
R158_652 s_2_340 s_2_339 0.108
R158_653 s_2_341 s_2_340 0.108
R158_654 s_2_342 s_2_341 0.108
R158_655 s_2_343 s_2_342 0.108
R158_656 s_2_344 s_2_343 0.108
R158_657 s_2_345 s_2_344 0.001
R158_658 s_2_347 s_2_346 0.001
R158_659 s_2_348 s_2_347 0.001
R158_660 s_2_352 s_2_348 0.001
R158_661 s_2_349 s_2_352 0.001
R158_662 s_2_350 s_2_349 0.001
R158_663 s_2_351 s_2_350 0.001
R158_664 s_2_353 s_2_352 1.296
R158_665 s_2_354 s_2_353 0.108
R158_666 s_2_355 s_2_354 0.108
R158_667 s_2_356 s_2_355 0.108
R158_668 s_2_357 s_2_356 0.108
R158_669 s_2_358 s_2_357 0.108
R158_670 s_2_359 s_2_358 0.108
R158_671 s_2_360 s_2_359 0.108
R158_672 s_2_361 s_2_360 0.864
R158_673 s_2_362 s_2_361 0.108
R158_674 s_2_363 s_2_362 0.108
R158_675 s_2_364 s_2_363 0.108
R158_676 s_2_365 s_2_364 0.108
R158_677 s_2_366 s_2_365 0.108
R158_678 s_2_367 s_2_366 0.108
R158_679 s_2_368 s_2_367 0.108
R158_680 s_2_369 s_2_368 0.108
R158_681 s_2_370 s_2_369 0.108
R158_682 s_2_371 s_2_370 0.108
R158_683 s_2_372 s_2_371 0.108
R158_684 s_2_373 s_2_372 0.108
R158_685 s_2_374 s_2_373 0.108
R158_686 s_2_375 s_2_374 0.108
R158_687 s_2_376 s_2_375 0.108
R158_688 s_2_377 s_2_376 0.108
R158_689 s_2_378 s_2_377 0.108
R158_690 s_2_379 s_2_378 0.108
R158_691 s_2_380 s_2_379 0.108
R158_692 s_2_381 s_2_380 0.001

C8158 s_2_352 vss 6.29069e-15
C8159 s_2 vss 6.29069e-15
C8160 s_2_27 vss 1.40901e-16
C8161 s_2_349 vss 1.40901e-16
C8162 s_2_28 vss 3.13114e-17
C8163 s_2_27 vss 3.13114e-17
C8164 s_2_29 vss 3.13114e-17
C8165 s_2_28 vss 3.13114e-17
C8166 s_2_30 vss 3.13114e-17
C8167 s_2_29 vss 3.13114e-17
C8168 s_2_31 vss 3.13114e-17
C8169 s_2_30 vss 3.13114e-17
C8170 s_2_32 vss 3.13114e-17
C8171 s_2_31 vss 3.13114e-17
C8172 s_2_33 vss 3.13114e-17
C8173 s_2_32 vss 3.13114e-17
C8174 s_2_34 vss 3.13114e-17
C8175 s_2_33 vss 3.13114e-17
C8176 s_2_35 vss 2.42663e-16
C8177 s_2_34 vss 2.42663e-16
C8178 s_2_36 vss 3.13114e-17
C8179 s_2_35 vss 3.13114e-17
C8180 s_2_37 vss 3.13114e-17
C8181 s_2_36 vss 3.13114e-17
C8182 s_2_38 vss 3.13114e-17
C8183 s_2_37 vss 3.13114e-17
C8184 s_2_39 vss 3.13114e-17
C8185 s_2_38 vss 3.13114e-17
C8186 s_2_40 vss 3.13114e-17
C8187 s_2_39 vss 3.13114e-17
C8188 s_2_41 vss 3.13114e-17
C8189 s_2_40 vss 3.13114e-17
C8190 s_2_42 vss 3.13114e-17
C8191 s_2_41 vss 3.13114e-17
C8192 s_2_43 vss 3.13114e-17
C8193 s_2_42 vss 3.13114e-17
C8194 s_2_44 vss 3.13114e-17
C8195 s_2_43 vss 3.13114e-17
C8196 s_2_45 vss 3.13114e-17
C8197 s_2_44 vss 3.13114e-17
C8198 s_2_46 vss 3.13114e-17
C8199 s_2_45 vss 3.13114e-17
C8200 s_2_47 vss 3.13114e-17
C8201 s_2_46 vss 3.13114e-17
C8202 s_2_48 vss 3.13114e-17
C8203 s_2_47 vss 3.13114e-17
C8204 s_2_49 vss 3.13114e-17
C8205 s_2_48 vss 3.13114e-17
C8206 s_2_50 vss 3.13114e-17
C8207 s_2_49 vss 3.13114e-17
C8208 s_2_51 vss 3.13114e-17
C8209 s_2_50 vss 3.13114e-17
C8210 s_2_52 vss 3.13114e-17
C8211 s_2_51 vss 3.13114e-17
C8212 s_2_53 vss 3.13114e-17
C8213 s_2_52 vss 3.13114e-17
C8214 s_2_54 vss 3.13114e-17
C8215 s_2_53 vss 3.13114e-17
C8216 s_2_55 vss 1.40901e-17
C8217 s_2_54 vss 1.40901e-17
C8218 s_2_56 vss 1.40901e-16
C8219 s_2_351 vss 1.40901e-16
C8220 s_2_57 vss 3.13114e-17
C8221 s_2_56 vss 3.13114e-17
C8222 s_2_58 vss 3.13114e-17
C8223 s_2_57 vss 3.13114e-17
C8224 s_2_59 vss 3.13114e-17
C8225 s_2_58 vss 3.13114e-17
C8226 s_2_60 vss 3.13114e-17
C8227 s_2_59 vss 3.13114e-17
C8228 s_2_61 vss 3.13114e-17
C8229 s_2_60 vss 3.13114e-17
C8230 s_2_62 vss 3.13114e-17
C8231 s_2_61 vss 3.13114e-17
C8232 s_2_63 vss 3.13114e-17
C8233 s_2_62 vss 3.13114e-17
C8234 s_2_64 vss 2.42663e-16
C8235 s_2_63 vss 2.42663e-16
C8236 s_2_65 vss 3.13114e-17
C8237 s_2_64 vss 3.13114e-17
C8238 s_2_66 vss 3.13114e-17
C8239 s_2_65 vss 3.13114e-17
C8240 s_2_67 vss 3.13114e-17
C8241 s_2_66 vss 3.13114e-17
C8242 s_2_68 vss 3.13114e-17
C8243 s_2_67 vss 3.13114e-17
C8244 s_2_69 vss 3.13114e-17
C8245 s_2_68 vss 3.13114e-17
C8246 s_2_70 vss 3.13114e-17
C8247 s_2_69 vss 3.13114e-17
C8248 s_2_71 vss 3.13114e-17
C8249 s_2_70 vss 3.13114e-17
C8250 s_2_72 vss 3.13114e-17
C8251 s_2_71 vss 3.13114e-17
C8252 s_2_73 vss 3.13114e-17
C8253 s_2_72 vss 3.13114e-17
C8254 s_2_74 vss 3.13114e-17
C8255 s_2_73 vss 3.13114e-17
C8256 s_2_75 vss 3.13114e-17
C8257 s_2_74 vss 3.13114e-17
C8258 s_2_76 vss 3.13114e-17
C8259 s_2_75 vss 3.13114e-17
C8260 s_2_77 vss 3.13114e-17
C8261 s_2_76 vss 3.13114e-17
C8262 s_2_78 vss 3.13114e-17
C8263 s_2_77 vss 3.13114e-17
C8264 s_2_79 vss 3.13114e-17
C8265 s_2_78 vss 3.13114e-17
C8266 s_2_80 vss 3.13114e-17
C8267 s_2_79 vss 3.13114e-17
C8268 s_2_81 vss 3.13114e-17
C8269 s_2_80 vss 3.13114e-17
C8270 s_2_82 vss 3.13114e-17
C8271 s_2_81 vss 3.13114e-17
C8272 s_2_83 vss 3.13114e-17
C8273 s_2_82 vss 3.13114e-17
C8274 s_2_84 vss 1.40901e-17
C8275 s_2_83 vss 1.40901e-17
C8276 s_2_85 vss 3.60081e-16
C8277 s_2_352 vss 3.60081e-16
C8278 s_2_86 vss 3.13114e-17
C8279 s_2_85 vss 3.13114e-17
C8280 s_2_87 vss 3.13114e-17
C8281 s_2_86 vss 3.13114e-17
C8282 s_2_88 vss 3.13114e-17
C8283 s_2_87 vss 3.13114e-17
C8284 s_2_89 vss 3.13114e-17
C8285 s_2_88 vss 3.13114e-17
C8286 s_2_90 vss 3.13114e-17
C8287 s_2_89 vss 3.13114e-17
C8288 s_2_91 vss 3.13114e-17
C8289 s_2_90 vss 3.13114e-17
C8290 s_2_92 vss 3.13114e-17
C8291 s_2_91 vss 3.13114e-17
C8292 s_2_93 vss 2.42663e-16
C8293 s_2_92 vss 2.42663e-16
C8294 s_2_94 vss 3.13114e-17
C8295 s_2_93 vss 3.13114e-17
C8296 s_2_95 vss 3.13114e-17
C8297 s_2_94 vss 3.13114e-17
C8298 s_2_96 vss 3.13114e-17
C8299 s_2_95 vss 3.13114e-17
C8300 s_2_97 vss 3.13114e-17
C8301 s_2_96 vss 3.13114e-17
C8302 s_2_98 vss 3.13114e-17
C8303 s_2_97 vss 3.13114e-17
C8304 s_2_99 vss 3.13114e-17
C8305 s_2_98 vss 3.13114e-17
C8306 s_2_100 vss 3.13114e-17
C8307 s_2_99 vss 3.13114e-17
C8308 s_2_101 vss 3.13114e-17
C8309 s_2_100 vss 3.13114e-17
C8310 s_2_102 vss 3.13114e-17
C8311 s_2_101 vss 3.13114e-17
C8312 s_2_103 vss 3.13114e-17
C8313 s_2_102 vss 3.13114e-17
C8314 s_2_104 vss 3.13114e-17
C8315 s_2_103 vss 3.13114e-17
C8316 s_2_105 vss 3.13114e-17
C8317 s_2_104 vss 3.13114e-17
C8318 s_2_106 vss 3.13114e-17
C8319 s_2_105 vss 3.13114e-17
C8320 s_2_107 vss 3.13114e-17
C8321 s_2_106 vss 3.13114e-17
C8322 s_2_108 vss 3.13114e-17
C8323 s_2_107 vss 3.13114e-17
C8324 s_2_109 vss 3.13114e-17
C8325 s_2_108 vss 3.13114e-17
C8326 s_2_110 vss 3.13114e-17
C8327 s_2_109 vss 3.13114e-17
C8328 s_2_111 vss 3.13114e-17
C8329 s_2_110 vss 3.13114e-17
C8330 s_2_112 vss 3.13114e-17
C8331 s_2_111 vss 3.13114e-17
C8332 s_2_113 vss 1.40901e-17
C8333 s_2_112 vss 1.40901e-17
C8334 s_2_114 vss 3.60081e-16
C8335 s_2_352 vss 3.60081e-16
C8336 s_2_115 vss 3.13114e-17
C8337 s_2_114 vss 3.13114e-17
C8338 s_2_116 vss 3.13114e-17
C8339 s_2_115 vss 3.13114e-17
C8340 s_2_117 vss 3.13114e-17
C8341 s_2_116 vss 3.13114e-17
C8342 s_2_118 vss 3.13114e-17
C8343 s_2_117 vss 3.13114e-17
C8344 s_2_119 vss 3.13114e-17
C8345 s_2_118 vss 3.13114e-17
C8346 s_2_120 vss 3.13114e-17
C8347 s_2_119 vss 3.13114e-17
C8348 s_2_121 vss 3.13114e-17
C8349 s_2_120 vss 3.13114e-17
C8350 s_2_122 vss 2.42663e-16
C8351 s_2_121 vss 2.42663e-16
C8352 s_2_123 vss 3.13114e-17
C8353 s_2_122 vss 3.13114e-17
C8354 s_2_124 vss 3.13114e-17
C8355 s_2_123 vss 3.13114e-17
C8356 s_2_125 vss 3.13114e-17
C8357 s_2_124 vss 3.13114e-17
C8358 s_2_126 vss 3.13114e-17
C8359 s_2_125 vss 3.13114e-17
C8360 s_2_127 vss 3.13114e-17
C8361 s_2_126 vss 3.13114e-17
C8362 s_2_128 vss 3.13114e-17
C8363 s_2_127 vss 3.13114e-17
C8364 s_2_129 vss 3.13114e-17
C8365 s_2_128 vss 3.13114e-17
C8366 s_2_130 vss 3.13114e-17
C8367 s_2_129 vss 3.13114e-17
C8368 s_2_131 vss 3.13114e-17
C8369 s_2_130 vss 3.13114e-17
C8370 s_2_132 vss 3.13114e-17
C8371 s_2_131 vss 3.13114e-17
C8372 s_2_133 vss 3.13114e-17
C8373 s_2_132 vss 3.13114e-17
C8374 s_2_134 vss 3.13114e-17
C8375 s_2_133 vss 3.13114e-17
C8376 s_2_135 vss 3.13114e-17
C8377 s_2_134 vss 3.13114e-17
C8378 s_2_136 vss 3.13114e-17
C8379 s_2_135 vss 3.13114e-17
C8380 s_2_137 vss 3.13114e-17
C8381 s_2_136 vss 3.13114e-17
C8382 s_2_138 vss 3.13114e-17
C8383 s_2_137 vss 3.13114e-17
C8384 s_2_139 vss 3.13114e-17
C8385 s_2_138 vss 3.13114e-17
C8386 s_2_140 vss 3.13114e-17
C8387 s_2_139 vss 3.13114e-17
C8388 s_2_141 vss 3.13114e-17
C8389 s_2_140 vss 3.13114e-17
C8390 s_2_142 vss 1.40901e-17
C8391 s_2_141 vss 1.40901e-17
C8392 s_2_143 vss 3.60081e-16
C8393 s_2_352 vss 3.60081e-16
C8394 s_2_144 vss 3.13114e-17
C8395 s_2_143 vss 3.13114e-17
C8396 s_2_145 vss 3.13114e-17
C8397 s_2_144 vss 3.13114e-17
C8398 s_2_146 vss 3.13114e-17
C8399 s_2_145 vss 3.13114e-17
C8400 s_2_147 vss 3.13114e-17
C8401 s_2_146 vss 3.13114e-17
C8402 s_2_148 vss 3.13114e-17
C8403 s_2_147 vss 3.13114e-17
C8404 s_2_149 vss 3.13114e-17
C8405 s_2_148 vss 3.13114e-17
C8406 s_2_150 vss 3.13114e-17
C8407 s_2_149 vss 3.13114e-17
C8408 s_2_151 vss 2.42663e-16
C8409 s_2_150 vss 2.42663e-16
C8410 s_2_152 vss 3.13114e-17
C8411 s_2_151 vss 3.13114e-17
C8412 s_2_153 vss 3.13114e-17
C8413 s_2_152 vss 3.13114e-17
C8414 s_2_154 vss 3.13114e-17
C8415 s_2_153 vss 3.13114e-17
C8416 s_2_155 vss 3.13114e-17
C8417 s_2_154 vss 3.13114e-17
C8418 s_2_156 vss 3.13114e-17
C8419 s_2_155 vss 3.13114e-17
C8420 s_2_157 vss 3.13114e-17
C8421 s_2_156 vss 3.13114e-17
C8422 s_2_158 vss 3.13114e-17
C8423 s_2_157 vss 3.13114e-17
C8424 s_2_159 vss 3.13114e-17
C8425 s_2_158 vss 3.13114e-17
C8426 s_2_160 vss 3.13114e-17
C8427 s_2_159 vss 3.13114e-17
C8428 s_2_161 vss 3.13114e-17
C8429 s_2_160 vss 3.13114e-17
C8430 s_2_162 vss 3.13114e-17
C8431 s_2_161 vss 3.13114e-17
C8432 s_2_163 vss 3.13114e-17
C8433 s_2_162 vss 3.13114e-17
C8434 s_2_164 vss 3.13114e-17
C8435 s_2_163 vss 3.13114e-17
C8436 s_2_165 vss 3.13114e-17
C8437 s_2_164 vss 3.13114e-17
C8438 s_2_166 vss 3.13114e-17
C8439 s_2_165 vss 3.13114e-17
C8440 s_2_167 vss 3.13114e-17
C8441 s_2_166 vss 3.13114e-17
C8442 s_2_168 vss 3.13114e-17
C8443 s_2_167 vss 3.13114e-17
C8444 s_2_169 vss 3.13114e-17
C8445 s_2_168 vss 3.13114e-17
C8446 s_2_170 vss 3.13114e-17
C8447 s_2_169 vss 3.13114e-17
C8448 s_2_171 vss 1.40901e-17
C8449 s_2_170 vss 1.40901e-17
C8450 s_2_172 vss 3.60081e-16
C8451 s_2_352 vss 3.60081e-16
C8452 s_2_173 vss 3.13114e-17
C8453 s_2_172 vss 3.13114e-17
C8454 s_2_174 vss 3.13114e-17
C8455 s_2_173 vss 3.13114e-17
C8456 s_2_175 vss 3.13114e-17
C8457 s_2_174 vss 3.13114e-17
C8458 s_2_176 vss 3.13114e-17
C8459 s_2_175 vss 3.13114e-17
C8460 s_2_177 vss 3.13114e-17
C8461 s_2_176 vss 3.13114e-17
C8462 s_2_178 vss 3.13114e-17
C8463 s_2_177 vss 3.13114e-17
C8464 s_2_179 vss 3.13114e-17
C8465 s_2_178 vss 3.13114e-17
C8466 s_2_180 vss 2.42663e-16
C8467 s_2_179 vss 2.42663e-16
C8468 s_2_181 vss 3.13114e-17
C8469 s_2_180 vss 3.13114e-17
C8470 s_2_182 vss 3.13114e-17
C8471 s_2_181 vss 3.13114e-17
C8472 s_2_183 vss 3.13114e-17
C8473 s_2_182 vss 3.13114e-17
C8474 s_2_184 vss 3.13114e-17
C8475 s_2_183 vss 3.13114e-17
C8476 s_2_185 vss 3.13114e-17
C8477 s_2_184 vss 3.13114e-17
C8478 s_2_186 vss 3.13114e-17
C8479 s_2_185 vss 3.13114e-17
C8480 s_2_187 vss 3.13114e-17
C8481 s_2_186 vss 3.13114e-17
C8482 s_2_188 vss 3.13114e-17
C8483 s_2_187 vss 3.13114e-17
C8484 s_2_189 vss 3.13114e-17
C8485 s_2_188 vss 3.13114e-17
C8486 s_2_190 vss 3.13114e-17
C8487 s_2_189 vss 3.13114e-17
C8488 s_2_191 vss 3.13114e-17
C8489 s_2_190 vss 3.13114e-17
C8490 s_2_192 vss 3.13114e-17
C8491 s_2_191 vss 3.13114e-17
C8492 s_2_193 vss 3.13114e-17
C8493 s_2_192 vss 3.13114e-17
C8494 s_2_194 vss 3.13114e-17
C8495 s_2_193 vss 3.13114e-17
C8496 s_2_195 vss 3.13114e-17
C8497 s_2_194 vss 3.13114e-17
C8498 s_2_196 vss 3.13114e-17
C8499 s_2_195 vss 3.13114e-17
C8500 s_2_197 vss 3.13114e-17
C8501 s_2_196 vss 3.13114e-17
C8502 s_2_198 vss 3.13114e-17
C8503 s_2_197 vss 3.13114e-17
C8504 s_2_199 vss 3.13114e-17
C8505 s_2_198 vss 3.13114e-17
C8506 s_2_200 vss 1.40901e-17
C8507 s_2_199 vss 1.40901e-17
C8508 s_2_201 vss 3.60081e-16
C8509 s_2_352 vss 3.60081e-16
C8510 s_2_202 vss 3.13114e-17
C8511 s_2_201 vss 3.13114e-17
C8512 s_2_203 vss 3.13114e-17
C8513 s_2_202 vss 3.13114e-17
C8514 s_2_204 vss 3.13114e-17
C8515 s_2_203 vss 3.13114e-17
C8516 s_2_205 vss 3.13114e-17
C8517 s_2_204 vss 3.13114e-17
C8518 s_2_206 vss 3.13114e-17
C8519 s_2_205 vss 3.13114e-17
C8520 s_2_207 vss 3.13114e-17
C8521 s_2_206 vss 3.13114e-17
C8522 s_2_208 vss 3.13114e-17
C8523 s_2_207 vss 3.13114e-17
C8524 s_2_209 vss 2.42663e-16
C8525 s_2_208 vss 2.42663e-16
C8526 s_2_210 vss 3.13114e-17
C8527 s_2_209 vss 3.13114e-17
C8528 s_2_211 vss 3.13114e-17
C8529 s_2_210 vss 3.13114e-17
C8530 s_2_212 vss 3.13114e-17
C8531 s_2_211 vss 3.13114e-17
C8532 s_2_213 vss 3.13114e-17
C8533 s_2_212 vss 3.13114e-17
C8534 s_2_214 vss 3.13114e-17
C8535 s_2_213 vss 3.13114e-17
C8536 s_2_215 vss 3.13114e-17
C8537 s_2_214 vss 3.13114e-17
C8538 s_2_216 vss 3.13114e-17
C8539 s_2_215 vss 3.13114e-17
C8540 s_2_217 vss 3.13114e-17
C8541 s_2_216 vss 3.13114e-17
C8542 s_2_218 vss 3.13114e-17
C8543 s_2_217 vss 3.13114e-17
C8544 s_2_219 vss 3.13114e-17
C8545 s_2_218 vss 3.13114e-17
C8546 s_2_220 vss 3.13114e-17
C8547 s_2_219 vss 3.13114e-17
C8548 s_2_221 vss 3.13114e-17
C8549 s_2_220 vss 3.13114e-17
C8550 s_2_222 vss 3.13114e-17
C8551 s_2_221 vss 3.13114e-17
C8552 s_2_223 vss 3.13114e-17
C8553 s_2_222 vss 3.13114e-17
C8554 s_2_224 vss 3.13114e-17
C8555 s_2_223 vss 3.13114e-17
C8556 s_2_225 vss 3.13114e-17
C8557 s_2_224 vss 3.13114e-17
C8558 s_2_226 vss 3.13114e-17
C8559 s_2_225 vss 3.13114e-17
C8560 s_2_227 vss 3.13114e-17
C8561 s_2_226 vss 3.13114e-17
C8562 s_2_228 vss 3.13114e-17
C8563 s_2_227 vss 3.13114e-17
C8564 s_2_229 vss 1.40901e-17
C8565 s_2_228 vss 1.40901e-17
C8566 s_2_230 vss 3.60081e-16
C8567 s_2_352 vss 3.60081e-16
C8568 s_2_231 vss 3.13114e-17
C8569 s_2_230 vss 3.13114e-17
C8570 s_2_232 vss 3.13114e-17
C8571 s_2_231 vss 3.13114e-17
C8572 s_2_233 vss 3.13114e-17
C8573 s_2_232 vss 3.13114e-17
C8574 s_2_234 vss 3.13114e-17
C8575 s_2_233 vss 3.13114e-17
C8576 s_2_235 vss 3.13114e-17
C8577 s_2_234 vss 3.13114e-17
C8578 s_2_236 vss 3.13114e-17
C8579 s_2_235 vss 3.13114e-17
C8580 s_2_237 vss 3.13114e-17
C8581 s_2_236 vss 3.13114e-17
C8582 s_2_238 vss 2.42663e-16
C8583 s_2_237 vss 2.42663e-16
C8584 s_2_239 vss 3.13114e-17
C8585 s_2_238 vss 3.13114e-17
C8586 s_2_240 vss 3.13114e-17
C8587 s_2_239 vss 3.13114e-17
C8588 s_2_241 vss 3.13114e-17
C8589 s_2_240 vss 3.13114e-17
C8590 s_2_242 vss 3.13114e-17
C8591 s_2_241 vss 3.13114e-17
C8592 s_2_243 vss 3.13114e-17
C8593 s_2_242 vss 3.13114e-17
C8594 s_2_244 vss 3.13114e-17
C8595 s_2_243 vss 3.13114e-17
C8596 s_2_245 vss 3.13114e-17
C8597 s_2_244 vss 3.13114e-17
C8598 s_2_246 vss 3.13114e-17
C8599 s_2_245 vss 3.13114e-17
C8600 s_2_247 vss 3.13114e-17
C8601 s_2_246 vss 3.13114e-17
C8602 s_2_248 vss 3.13114e-17
C8603 s_2_247 vss 3.13114e-17
C8604 s_2_249 vss 3.13114e-17
C8605 s_2_248 vss 3.13114e-17
C8606 s_2_250 vss 3.13114e-17
C8607 s_2_249 vss 3.13114e-17
C8608 s_2_251 vss 3.13114e-17
C8609 s_2_250 vss 3.13114e-17
C8610 s_2_252 vss 3.13114e-17
C8611 s_2_251 vss 3.13114e-17
C8612 s_2_253 vss 3.13114e-17
C8613 s_2_252 vss 3.13114e-17
C8614 s_2_254 vss 3.13114e-17
C8615 s_2_253 vss 3.13114e-17
C8616 s_2_255 vss 3.13114e-17
C8617 s_2_254 vss 3.13114e-17
C8618 s_2_256 vss 3.13114e-17
C8619 s_2_255 vss 3.13114e-17
C8620 s_2_257 vss 3.13114e-17
C8621 s_2_256 vss 3.13114e-17
C8622 s_2_258 vss 1.40901e-17
C8623 s_2_257 vss 1.40901e-17
C8624 s_2_259 vss 3.60081e-16
C8625 s_2_352 vss 3.60081e-16
C8626 s_2_260 vss 3.13114e-17
C8627 s_2_259 vss 3.13114e-17
C8628 s_2_261 vss 3.13114e-17
C8629 s_2_260 vss 3.13114e-17
C8630 s_2_262 vss 3.13114e-17
C8631 s_2_261 vss 3.13114e-17
C8632 s_2_263 vss 3.13114e-17
C8633 s_2_262 vss 3.13114e-17
C8634 s_2_264 vss 3.13114e-17
C8635 s_2_263 vss 3.13114e-17
C8636 s_2_265 vss 3.13114e-17
C8637 s_2_264 vss 3.13114e-17
C8638 s_2_266 vss 3.13114e-17
C8639 s_2_265 vss 3.13114e-17
C8640 s_2_267 vss 2.42663e-16
C8641 s_2_266 vss 2.42663e-16
C8642 s_2_268 vss 3.13114e-17
C8643 s_2_267 vss 3.13114e-17
C8644 s_2_269 vss 3.13114e-17
C8645 s_2_268 vss 3.13114e-17
C8646 s_2_270 vss 3.13114e-17
C8647 s_2_269 vss 3.13114e-17
C8648 s_2_271 vss 3.13114e-17
C8649 s_2_270 vss 3.13114e-17
C8650 s_2_272 vss 3.13114e-17
C8651 s_2_271 vss 3.13114e-17
C8652 s_2_273 vss 3.13114e-17
C8653 s_2_272 vss 3.13114e-17
C8654 s_2_274 vss 3.13114e-17
C8655 s_2_273 vss 3.13114e-17
C8656 s_2_275 vss 3.13114e-17
C8657 s_2_274 vss 3.13114e-17
C8658 s_2_276 vss 3.13114e-17
C8659 s_2_275 vss 3.13114e-17
C8660 s_2_277 vss 3.13114e-17
C8661 s_2_276 vss 3.13114e-17
C8662 s_2_278 vss 3.13114e-17
C8663 s_2_277 vss 3.13114e-17
C8664 s_2_279 vss 3.13114e-17
C8665 s_2_278 vss 3.13114e-17
C8666 s_2_280 vss 3.13114e-17
C8667 s_2_279 vss 3.13114e-17
C8668 s_2_281 vss 3.13114e-17
C8669 s_2_280 vss 3.13114e-17
C8670 s_2_282 vss 3.13114e-17
C8671 s_2_281 vss 3.13114e-17
C8672 s_2_283 vss 3.13114e-17
C8673 s_2_282 vss 3.13114e-17
C8674 s_2_284 vss 3.13114e-17
C8675 s_2_283 vss 3.13114e-17
C8676 s_2_285 vss 3.13114e-17
C8677 s_2_284 vss 3.13114e-17
C8678 s_2_286 vss 3.13114e-17
C8679 s_2_285 vss 3.13114e-17
C8680 s_2_287 vss 1.40901e-17
C8681 s_2_286 vss 1.40901e-17
C8682 s_2_288 vss 1.40901e-16
C8683 s_2_346 vss 1.40901e-16
C8684 s_2_289 vss 3.13114e-17
C8685 s_2_288 vss 3.13114e-17
C8686 s_2_290 vss 3.13114e-17
C8687 s_2_289 vss 3.13114e-17
C8688 s_2_291 vss 3.13114e-17
C8689 s_2_290 vss 3.13114e-17
C8690 s_2_292 vss 3.13114e-17
C8691 s_2_291 vss 3.13114e-17
C8692 s_2_293 vss 3.13114e-17
C8693 s_2_292 vss 3.13114e-17
C8694 s_2_294 vss 3.13114e-17
C8695 s_2_293 vss 3.13114e-17
C8696 s_2_295 vss 3.13114e-17
C8697 s_2_294 vss 3.13114e-17
C8698 s_2_296 vss 2.42663e-16
C8699 s_2_295 vss 2.42663e-16
C8700 s_2_297 vss 3.13114e-17
C8701 s_2_296 vss 3.13114e-17
C8702 s_2_298 vss 3.13114e-17
C8703 s_2_297 vss 3.13114e-17
C8704 s_2_299 vss 3.13114e-17
C8705 s_2_298 vss 3.13114e-17
C8706 s_2_300 vss 3.13114e-17
C8707 s_2_299 vss 3.13114e-17
C8708 s_2_301 vss 3.13114e-17
C8709 s_2_300 vss 3.13114e-17
C8710 s_2_302 vss 3.13114e-17
C8711 s_2_301 vss 3.13114e-17
C8712 s_2_303 vss 3.13114e-17
C8713 s_2_302 vss 3.13114e-17
C8714 s_2_304 vss 3.13114e-17
C8715 s_2_303 vss 3.13114e-17
C8716 s_2_305 vss 3.13114e-17
C8717 s_2_304 vss 3.13114e-17
C8718 s_2_306 vss 3.13114e-17
C8719 s_2_305 vss 3.13114e-17
C8720 s_2_307 vss 3.13114e-17
C8721 s_2_306 vss 3.13114e-17
C8722 s_2_308 vss 3.13114e-17
C8723 s_2_307 vss 3.13114e-17
C8724 s_2_309 vss 3.13114e-17
C8725 s_2_308 vss 3.13114e-17
C8726 s_2_310 vss 3.13114e-17
C8727 s_2_309 vss 3.13114e-17
C8728 s_2_311 vss 3.13114e-17
C8729 s_2_310 vss 3.13114e-17
C8730 s_2_312 vss 3.13114e-17
C8731 s_2_311 vss 3.13114e-17
C8732 s_2_313 vss 3.13114e-17
C8733 s_2_312 vss 3.13114e-17
C8734 s_2_314 vss 3.13114e-17
C8735 s_2_313 vss 3.13114e-17
C8736 s_2_315 vss 3.13114e-17
C8737 s_2_314 vss 3.13114e-17
C8738 s_2_316 vss 1.40901e-17
C8739 s_2_315 vss 1.40901e-17
C8740 s_2_317 vss 1.40901e-16
C8741 s_2_348 vss 1.40901e-16
C8742 s_2_318 vss 3.13114e-17
C8743 s_2_317 vss 3.13114e-17
C8744 s_2_319 vss 3.13114e-17
C8745 s_2_318 vss 3.13114e-17
C8746 s_2_320 vss 3.13114e-17
C8747 s_2_319 vss 3.13114e-17
C8748 s_2_321 vss 3.13114e-17
C8749 s_2_320 vss 3.13114e-17
C8750 s_2_322 vss 3.13114e-17
C8751 s_2_321 vss 3.13114e-17
C8752 s_2_323 vss 3.13114e-17
C8753 s_2_322 vss 3.13114e-17
C8754 s_2_324 vss 3.13114e-17
C8755 s_2_323 vss 3.13114e-17
C8756 s_2_325 vss 2.42663e-16
C8757 s_2_324 vss 2.42663e-16
C8758 s_2_326 vss 3.13114e-17
C8759 s_2_325 vss 3.13114e-17
C8760 s_2_327 vss 3.13114e-17
C8761 s_2_326 vss 3.13114e-17
C8762 s_2_328 vss 3.13114e-17
C8763 s_2_327 vss 3.13114e-17
C8764 s_2_329 vss 3.13114e-17
C8765 s_2_328 vss 3.13114e-17
C8766 s_2_330 vss 3.13114e-17
C8767 s_2_329 vss 3.13114e-17
C8768 s_2_331 vss 3.13114e-17
C8769 s_2_330 vss 3.13114e-17
C8770 s_2_332 vss 3.13114e-17
C8771 s_2_331 vss 3.13114e-17
C8772 s_2_333 vss 3.13114e-17
C8773 s_2_332 vss 3.13114e-17
C8774 s_2_334 vss 3.13114e-17
C8775 s_2_333 vss 3.13114e-17
C8776 s_2_335 vss 3.13114e-17
C8777 s_2_334 vss 3.13114e-17
C8778 s_2_336 vss 3.13114e-17
C8779 s_2_335 vss 3.13114e-17
C8780 s_2_337 vss 3.13114e-17
C8781 s_2_336 vss 3.13114e-17
C8782 s_2_338 vss 3.13114e-17
C8783 s_2_337 vss 3.13114e-17
C8784 s_2_339 vss 3.13114e-17
C8785 s_2_338 vss 3.13114e-17
C8786 s_2_340 vss 3.13114e-17
C8787 s_2_339 vss 3.13114e-17
C8788 s_2_341 vss 3.13114e-17
C8789 s_2_340 vss 3.13114e-17
C8790 s_2_342 vss 3.13114e-17
C8791 s_2_341 vss 3.13114e-17
C8792 s_2_343 vss 3.13114e-17
C8793 s_2_342 vss 3.13114e-17
C8794 s_2_344 vss 3.13114e-17
C8795 s_2_343 vss 3.13114e-17
C8796 s_2_345 vss 1.40901e-17
C8797 s_2_344 vss 1.40901e-17
C8798 s_2_347 vss 2.95333e-17
C8799 s_2_346 vss 2.95333e-17
C8800 s_2_348 vss 3.71708e-16
C8801 s_2_347 vss 3.71708e-16
C8802 s_2_352 vss 2.15831e-15
C8803 s_2_348 vss 2.15831e-15
C8804 s_2_349 vss 2.15831e-15
C8805 s_2_352 vss 2.15831e-15
C8806 s_2_350 vss 3.71708e-16
C8807 s_2_349 vss 3.71708e-16
C8808 s_2_351 vss 2.95333e-17
C8809 s_2_350 vss 2.95333e-17
C8810 s_2_353 vss 3.60081e-16
C8811 s_2_352 vss 3.60081e-16
C8812 s_2_354 vss 3.13114e-17
C8813 s_2_353 vss 3.13114e-17
C8814 s_2_355 vss 3.13114e-17
C8815 s_2_354 vss 3.13114e-17
C8816 s_2_356 vss 3.13114e-17
C8817 s_2_355 vss 3.13114e-17
C8818 s_2_357 vss 3.13114e-17
C8819 s_2_356 vss 3.13114e-17
C8820 s_2_358 vss 3.13114e-17
C8821 s_2_357 vss 3.13114e-17
C8822 s_2_359 vss 3.13114e-17
C8823 s_2_358 vss 3.13114e-17
C8824 s_2_360 vss 3.13114e-17
C8825 s_2_359 vss 3.13114e-17
C8826 s_2_361 vss 2.42663e-16
C8827 s_2_360 vss 2.42663e-16
C8828 s_2_362 vss 3.13114e-17
C8829 s_2_361 vss 3.13114e-17
C8830 s_2_363 vss 3.13114e-17
C8831 s_2_362 vss 3.13114e-17
C8832 s_2_364 vss 3.13114e-17
C8833 s_2_363 vss 3.13114e-17
C8834 s_2_365 vss 3.13114e-17
C8835 s_2_364 vss 3.13114e-17
C8836 s_2_366 vss 3.13114e-17
C8837 s_2_365 vss 3.13114e-17
C8838 s_2_367 vss 3.13114e-17
C8839 s_2_366 vss 3.13114e-17
C8840 s_2_368 vss 3.13114e-17
C8841 s_2_367 vss 3.13114e-17
C8842 s_2_369 vss 3.13114e-17
C8843 s_2_368 vss 3.13114e-17
C8844 s_2_370 vss 3.13114e-17
C8845 s_2_369 vss 3.13114e-17
C8846 s_2_371 vss 3.13114e-17
C8847 s_2_370 vss 3.13114e-17
C8848 s_2_372 vss 3.13114e-17
C8849 s_2_371 vss 3.13114e-17
C8850 s_2_373 vss 3.13114e-17
C8851 s_2_372 vss 3.13114e-17
C8852 s_2_374 vss 3.13114e-17
C8853 s_2_373 vss 3.13114e-17
C8854 s_2_375 vss 3.13114e-17
C8855 s_2_374 vss 3.13114e-17
C8856 s_2_376 vss 3.13114e-17
C8857 s_2_375 vss 3.13114e-17
C8858 s_2_377 vss 3.13114e-17
C8859 s_2_376 vss 3.13114e-17
C8860 s_2_378 vss 3.13114e-17
C8861 s_2_377 vss 3.13114e-17
C8862 s_2_379 vss 3.13114e-17
C8863 s_2_378 vss 3.13114e-17
C8864 s_2_380 vss 3.13114e-17
C8865 s_2_379 vss 3.13114e-17
C8866 s_2_381 vss 1.40901e-17
C8867 s_2_380 vss 1.40901e-17

R159_1 n5912_3 n5912_153 0.001
R159_2 n5912_123 n5912_8 0.001
R159_3 n5912_7 n5912_11 0.001
R159_4 n5912_152 n5912_18 0.001
R159_5 n5912_115 n5912_27 0.001
R159_6 n5912_26 n5912 0.001
R159_7 n5912_29 n5912 0.001
R159_8 n5912_28 n5912 0.001
R159_9 n5912_23 n5912 0.001
R159_10 n5912_25 n5912 0.001
R159_11 n5912_24 n5912 0.001
R159_12 n5912_140 n5912_31 0.001
R159_13 n5912_141 n5912_31 0.001
R159_14 n5912_143 n5912_31 0.001
R159_15 n5912_142 n5912_31 0.001
R159_16 n5912_139 n5912_31 0.001
R159_17 n5912_136 n5912_31 0.001
R159_18 n5912_137 n5912_31 0.001
R159_19 n5912_138 n5912_31 0.001
R159_20 n5912_132 n5912_31 0.001
R159_21 n5912_134 n5912_31 0.001
R159_22 n5912_135 n5912_31 0.001
R159_23 n5912_133 n5912_31 0.001
R159_24 n5912_129 n5912_31 0.001
R159_25 n5912_130 n5912_31 0.001
R159_26 n5912_131 n5912_31 0.001
R159_27 n5912_122 n5912_33 0.001
R159_28 n5912_32 n5912_36 0.001
R159_29 n5912_114 n5912_46 0.001
R159_30 n5912_45 n5912_41 0.001
R159_31 n5912_47 n5912_41 0.001
R159_32 n5912_48 n5912_41 0.001
R159_33 n5912_44 n5912_41 0.001
R159_34 n5912_43 n5912_41 0.001
R159_35 n5912_42 n5912_41 0.001
R159_36 n5912_166 n5912_50 0.001
R159_37 n5912_167 n5912_50 0.001
R159_38 n5912_168 n5912_50 0.001
R159_39 n5912_169 n5912_50 0.001
R159_40 n5912_162 n5912_50 0.001
R159_41 n5912_163 n5912_50 0.001
R159_42 n5912_164 n5912_50 0.001
R159_43 n5912_165 n5912_50 0.001
R159_44 n5912_158 n5912_50 0.001
R159_45 n5912_161 n5912_50 0.001
R159_46 n5912_159 n5912_50 0.001
R159_47 n5912_160 n5912_50 0.001
R159_48 n5912_155 n5912_50 0.001
R159_49 n5912_156 n5912_50 0.001
R159_50 n5912_157 n5912_50 0.001
R159_51 n5912_150 n5912_53 0.001
R159_52 n5912_121 n5912_58 0.001
R159_53 n5912_57 n5912_61 0.001
R159_54 n5912_149 n5912_68 0.001
R159_55 n5912_120 n5912_73 0.001
R159_56 n5912_72 n5912_76 0.001
R159_57 n5912_148 n5912_83 0.001
R159_58 n5912_119 n5912_88 0.001
R159_59 n5912_87 n5912_91 0.001
R159_60 n5912_147 n5912_98 0.001
R159_61 n5912_118 n5912_103 0.001
R159_62 n5912_102 n5912_106 0.001
R159_63 n5912_145 n5912_111 0.001
R159_64 n5912_124 n5912_112 0.001
R159_65 n5912_125 n5912_113 0.001
R159_66 n5912_144 n5912_116 0.001
R159_67 n5912_127 n5912_117 0.001
R159_68 n5912_10 n5912_9 21.6
R159_69 n5912_13 n5912_10 21.6
R159_70 n5912_14 n5912_13 43.2
R159_71 n5912_15 n5912_14 43.2
R159_72 n5912_35 n5912_34 21.6
R159_73 n5912_38 n5912_35 21.6
R159_74 n5912_39 n5912_38 43.2
R159_75 n5912_40 n5912_39 43.2
R159_76 n5912_60 n5912_59 21.6
R159_77 n5912_63 n5912_60 21.6
R159_78 n5912_64 n5912_63 43.2
R159_79 n5912_65 n5912_64 43.2
R159_80 n5912_90 n5912_89 21.6
R159_81 n5912_93 n5912_90 21.6
R159_82 n5912_94 n5912_93 43.2
R159_83 n5912_95 n5912_94 43.2
R159_84 n5912_75 n5912_74 21.6
R159_85 n5912_78 n5912_75 21.6
R159_86 n5912_79 n5912_78 43.2
R159_87 n5912_80 n5912_79 43.2
R159_88 n5912_105 n5912_104 21.6
R159_89 n5912_108 n5912_105 21.6
R159_90 n5912_109 n5912_108 43.2
R159_91 n5912_110 n5912_109 43.2
R159_92 n5912_12 n5912_10 28.8
R159_93 n5912_37 n5912_35 28.8
R159_94 n5912_62 n5912_60 28.8
R159_95 n5912_92 n5912_90 28.8
R159_96 n5912_77 n5912_75 28.8
R159_97 n5912_107 n5912_105 28.8
R159_98 n5912_12 n5912_11 7.2
R159_99 n5912_37 n5912_36 7.2
R159_100 n5912_62 n5912_61 7.2
R159_101 n5912_92 n5912_91 7.2
R159_102 n5912_77 n5912_76 7.2
R159_103 n5912_107 n5912_106 7.2
R159_104 n5912_24 n5912_23 0.108
R159_105 n5912_25 n5912_24 0.108
R159_106 n5912_26 n5912_25 0.108
R159_107 n5912_27 n5912_26 0.108
R159_108 n5912_28 n5912_27 0.108
R159_109 n5912_29 n5912_28 0.108
R159_110 n5912_30 n5912_29 0.001
R159_111 n5912_43 n5912_42 0.108
R159_112 n5912_44 n5912_43 0.108
R159_113 n5912_45 n5912_44 0.108
R159_114 n5912_46 n5912_45 0.108
R159_115 n5912_47 n5912_46 0.108
R159_116 n5912_48 n5912_47 0.108
R159_117 n5912_49 n5912_48 0.001
R159_118 n5912_8 n5912_7 0.216
R159_119 n5912_33 n5912_32 0.216
R159_120 n5912_58 n5912_57 0.216
R159_121 n5912_88 n5912_87 0.216
R159_122 n5912_73 n5912_72 0.216
R159_123 n5912_103 n5912_102 0.216
R159_124 n5912_17 n5912_16 21.6
R159_125 n5912_19 n5912_17 21.6
R159_126 n5912_20 n5912_19 43.2
R159_127 n5912_21 n5912_20 43.2
R159_128 n5912_67 n5912_66 21.6
R159_129 n5912_69 n5912_67 21.6
R159_130 n5912_70 n5912_69 43.2
R159_131 n5912_71 n5912_70 43.2
R159_132 n5912_52 n5912_51 21.6
R159_133 n5912_54 n5912_52 21.6
R159_134 n5912_55 n5912_54 43.2
R159_135 n5912_56 n5912_55 43.2
R159_136 n5912_82 n5912_81 21.6
R159_137 n5912_84 n5912_82 21.6
R159_138 n5912_85 n5912_84 43.2
R159_139 n5912_86 n5912_85 43.2
R159_140 n5912_97 n5912_96 21.6
R159_141 n5912_99 n5912_97 21.6
R159_142 n5912_100 n5912_99 43.2
R159_143 n5912_101 n5912_100 43.2
R159_144 n5912_18 n5912_17 28.8
R159_145 n5912_68 n5912_67 28.8
R159_146 n5912_53 n5912_52 28.8
R159_147 n5912_83 n5912_82 28.8
R159_148 n5912_98 n5912_97 28.8
R159_149 n5912_112 n5912_111 0.054
R159_150 n5912_113 n5912_112 0.054
R159_151 n5912_114 n5912_113 1.458
R159_152 n5912_115 n5912_114 0.216
R159_153 n5912_117 n5912_116 0.054
R159_154 n5912_118 n5912_117 0.108
R159_155 n5912_119 n5912_118 0.432
R159_156 n5912_120 n5912_119 0.432
R159_157 n5912_121 n5912_120 0.432
R159_158 n5912_122 n5912_121 0.432
R159_159 n5912_123 n5912_122 0.432
R159_160 n5912_124 n5912_145 0.108
R159_161 n5912_125 n5912_124 0.108
R159_162 n5912_126 n5912_125 0.001
R159_163 n5912_127 n5912_144 0.108
R159_164 n5912_128 n5912_127 0.001
R159_165 n5912_129 n5912_151 0.648
R159_166 n5912_130 n5912_129 0.108
R159_167 n5912_131 n5912_130 0.108
R159_168 n5912_132 n5912_131 0.108
R159_169 n5912_133 n5912_132 0.108
R159_170 n5912_134 n5912_133 0.108
R159_171 n5912_135 n5912_134 0.108
R159_172 n5912_136 n5912_135 0.108
R159_173 n5912_137 n5912_136 0.108
R159_174 n5912_138 n5912_137 0.108
R159_175 n5912_139 n5912_138 0.108
R159_176 n5912_140 n5912_139 0.108
R159_177 n5912_141 n5912_140 0.108
R159_178 n5912_142 n5912_141 0.108
R159_179 n5912_143 n5912_142 0.108
R159_180 n5912_155 n5912_150 0.648
R159_181 n5912_156 n5912_155 0.108
R159_182 n5912_157 n5912_156 0.108
R159_183 n5912_158 n5912_157 0.108
R159_184 n5912_159 n5912_158 0.108
R159_185 n5912_160 n5912_159 0.108
R159_186 n5912_161 n5912_160 0.108
R159_187 n5912_162 n5912_161 0.108
R159_188 n5912_163 n5912_162 0.108
R159_189 n5912_164 n5912_163 0.108
R159_190 n5912_165 n5912_164 0.108
R159_191 n5912_166 n5912_165 0.108
R159_192 n5912_167 n5912_166 0.108
R159_193 n5912_168 n5912_167 0.108
R159_194 n5912_169 n5912_168 0.108
R159_195 n5912_146 n5912_144 3.024
R159_196 n5912_145 n5912_146 3.348
R159_197 n5912_147 n5912_146 0.432
R159_198 n5912_148 n5912_147 0.648
R159_199 n5912_149 n5912_148 0.648
R159_200 n5912_150 n5912_149 0.648
R159_201 n5912_151 n5912_150 0.324
R159_202 n5912_152 n5912_151 0.216
R159_203 n5912_153 n5912_152 0.648
R159_204 n5912_154 n5912_153 0.001
R159_205 n5912_2 n5912_1 21.6
R159_206 n5912_4 n5912_2 21.6
R159_207 n5912_5 n5912_4 43.2
R159_208 n5912_6 n5912_5 43.2
R159_209 n5912_3 n5912_2 28.8

C8868 n5912_10 vss 2.34738e-17
C8869 n5912_9 vss 2.34738e-17
C8870 n5912_13 vss 2.34738e-17
C8871 n5912_10 vss 2.34738e-17
C8872 n5912_14 vss 4.69476e-17
C8873 n5912_13 vss 4.69476e-17
C8874 n5912_15 vss 4.69476e-17
C8875 n5912_14 vss 4.69476e-17
C8876 n5912_35 vss 2.34738e-17
C8877 n5912_34 vss 2.34738e-17
C8878 n5912_38 vss 2.34738e-17
C8879 n5912_35 vss 2.34738e-17
C8880 n5912_39 vss 4.69476e-17
C8881 n5912_38 vss 4.69476e-17
C8882 n5912_40 vss 4.69476e-17
C8883 n5912_39 vss 4.69476e-17
C8884 n5912_60 vss 2.34738e-17
C8885 n5912_59 vss 2.34738e-17
C8886 n5912_63 vss 2.34738e-17
C8887 n5912_60 vss 2.34738e-17
C8888 n5912_64 vss 4.69476e-17
C8889 n5912_63 vss 4.69476e-17
C8890 n5912_65 vss 4.69476e-17
C8891 n5912_64 vss 4.69476e-17
C8892 n5912_90 vss 2.34738e-17
C8893 n5912_89 vss 2.34738e-17
C8894 n5912_93 vss 2.34738e-17
C8895 n5912_90 vss 2.34738e-17
C8896 n5912_94 vss 4.69476e-17
C8897 n5912_93 vss 4.69476e-17
C8898 n5912_95 vss 4.69476e-17
C8899 n5912_94 vss 4.69476e-17
C8900 n5912_75 vss 2.34738e-17
C8901 n5912_74 vss 2.34738e-17
C8902 n5912_78 vss 2.34738e-17
C8903 n5912_75 vss 2.34738e-17
C8904 n5912_79 vss 4.69476e-17
C8905 n5912_78 vss 4.69476e-17
C8906 n5912_80 vss 4.69476e-17
C8907 n5912_79 vss 4.69476e-17
C8908 n5912_105 vss 2.34738e-17
C8909 n5912_104 vss 2.34738e-17
C8910 n5912_108 vss 2.34738e-17
C8911 n5912_105 vss 2.34738e-17
C8912 n5912_109 vss 4.69476e-17
C8913 n5912_108 vss 4.69476e-17
C8914 n5912_110 vss 4.69476e-17
C8915 n5912_109 vss 4.69476e-17
C8916 n5912_12 vss 7.33536e-17
C8917 n5912_10 vss 7.33536e-17
C8918 n5912_37 vss 7.33536e-17
C8919 n5912_35 vss 7.33536e-17
C8920 n5912_62 vss 7.33536e-17
C8921 n5912_60 vss 7.33536e-17
C8922 n5912_92 vss 7.33536e-17
C8923 n5912_90 vss 7.33536e-17
C8924 n5912_77 vss 7.33536e-17
C8925 n5912_75 vss 7.33536e-17
C8926 n5912_107 vss 7.33536e-17
C8927 n5912_105 vss 7.33536e-17
C8928 n5912_12 vss 5.2569e-17
C8929 n5912_11 vss 5.2569e-17
C8930 n5912_37 vss 5.2569e-17
C8931 n5912_36 vss 5.2569e-17
C8932 n5912_62 vss 5.2569e-17
C8933 n5912_61 vss 5.2569e-17
C8934 n5912_92 vss 5.2569e-17
C8935 n5912_91 vss 5.2569e-17
C8936 n5912_77 vss 5.2569e-17
C8937 n5912_76 vss 5.2569e-17
C8938 n5912_107 vss 5.2569e-17
C8939 n5912_106 vss 5.2569e-17
C8940 n5912_24 vss 2.92378e-17
C8941 n5912_23 vss 2.92378e-17
C8942 n5912_25 vss 2.92378e-17
C8943 n5912_24 vss 2.92378e-17
C8944 n5912_26 vss 2.92378e-17
C8945 n5912_25 vss 2.92378e-17
C8946 n5912_27 vss 3.65472e-17
C8947 n5912_26 vss 3.65472e-17
C8948 n5912_28 vss 2.92378e-17
C8949 n5912_27 vss 2.92378e-17
C8950 n5912_29 vss 3.65472e-17
C8951 n5912_28 vss 3.65472e-17
C8952 n5912_30 vss 1.3157e-17
C8953 n5912_29 vss 1.3157e-17
C8954 n5912_43 vss 2.92378e-17
C8955 n5912_42 vss 2.92378e-17
C8956 n5912_44 vss 2.92378e-17
C8957 n5912_43 vss 2.92378e-17
C8958 n5912_45 vss 2.92378e-17
C8959 n5912_44 vss 2.92378e-17
C8960 n5912_46 vss 3.65472e-17
C8961 n5912_45 vss 3.65472e-17
C8962 n5912_47 vss 2.92378e-17
C8963 n5912_46 vss 2.92378e-17
C8964 n5912_48 vss 3.65472e-17
C8965 n5912_47 vss 3.65472e-17
C8966 n5912_49 vss 1.3157e-17
C8967 n5912_48 vss 1.3157e-17
C8968 n5912_8 vss 4.38566e-17
C8969 n5912_7 vss 4.38566e-17
C8970 n5912_33 vss 4.38566e-17
C8971 n5912_32 vss 4.38566e-17
C8972 n5912_58 vss 4.38566e-17
C8973 n5912_57 vss 4.38566e-17
C8974 n5912_88 vss 4.38566e-17
C8975 n5912_87 vss 4.38566e-17
C8976 n5912_73 vss 4.38566e-17
C8977 n5912_72 vss 4.38566e-17
C8978 n5912_103 vss 4.38566e-17
C8979 n5912_102 vss 4.38566e-17
C8980 n5912_17 vss 2.34738e-17
C8981 n5912_16 vss 2.34738e-17
C8982 n5912_19 vss 2.34738e-17
C8983 n5912_17 vss 2.34738e-17
C8984 n5912_20 vss 4.69476e-17
C8985 n5912_19 vss 4.69476e-17
C8986 n5912_21 vss 4.69476e-17
C8987 n5912_20 vss 4.69476e-17
C8988 n5912_67 vss 2.34738e-17
C8989 n5912_66 vss 2.34738e-17
C8990 n5912_69 vss 2.34738e-17
C8991 n5912_67 vss 2.34738e-17
C8992 n5912_70 vss 4.69476e-17
C8993 n5912_69 vss 4.69476e-17
C8994 n5912_71 vss 4.69476e-17
C8995 n5912_70 vss 4.69476e-17
C8996 n5912_52 vss 2.34738e-17
C8997 n5912_51 vss 2.34738e-17
C8998 n5912_54 vss 2.34738e-17
C8999 n5912_52 vss 2.34738e-17
C9000 n5912_55 vss 4.69476e-17
C9001 n5912_54 vss 4.69476e-17
C9002 n5912_56 vss 4.69476e-17
C9003 n5912_55 vss 4.69476e-17
C9004 n5912_82 vss 2.34738e-17
C9005 n5912_81 vss 2.34738e-17
C9006 n5912_84 vss 2.34738e-17
C9007 n5912_82 vss 2.34738e-17
C9008 n5912_85 vss 4.69476e-17
C9009 n5912_84 vss 4.69476e-17
C9010 n5912_86 vss 4.69476e-17
C9011 n5912_85 vss 4.69476e-17
C9012 n5912_97 vss 2.34738e-17
C9013 n5912_96 vss 2.34738e-17
C9014 n5912_99 vss 2.34738e-17
C9015 n5912_97 vss 2.34738e-17
C9016 n5912_100 vss 4.69476e-17
C9017 n5912_99 vss 4.69476e-17
C9018 n5912_101 vss 4.69476e-17
C9019 n5912_100 vss 4.69476e-17
C9020 n5912_18 vss 7.33536e-17
C9021 n5912_17 vss 7.33536e-17
C9022 n5912_68 vss 7.33536e-17
C9023 n5912_67 vss 7.33536e-17
C9024 n5912_53 vss 7.33536e-17
C9025 n5912_52 vss 7.33536e-17
C9026 n5912_83 vss 7.33536e-17
C9027 n5912_82 vss 7.33536e-17
C9028 n5912_98 vss 7.33536e-17
C9029 n5912_97 vss 7.33536e-17
C9030 n5912_112 vss 2.60496e-17
C9031 n5912_111 vss 2.60496e-17
C9032 n5912_113 vss 2.60496e-17
C9033 n5912_112 vss 2.60496e-17
C9034 n5912_114 vss 5.40529e-16
C9035 n5912_113 vss 5.40529e-16
C9036 n5912_115 vss 7.81488e-17
C9037 n5912_114 vss 7.81488e-17
C9038 n5912_117 vss 3.2562e-17
C9039 n5912_116 vss 3.2562e-17
C9040 n5912_118 vss 4.55868e-17
C9041 n5912_117 vss 4.55868e-17
C9042 n5912_119 vss 1.56298e-16
C9043 n5912_118 vss 1.56298e-16
C9044 n5912_120 vss 1.56298e-16
C9045 n5912_119 vss 1.56298e-16
C9046 n5912_121 vss 1.56298e-16
C9047 n5912_120 vss 1.56298e-16
C9048 n5912_122 vss 1.56298e-16
C9049 n5912_121 vss 1.56298e-16
C9050 n5912_123 vss 1.56298e-16
C9051 n5912_122 vss 1.56298e-16
C9052 n5912_124 vss 3.13114e-17
C9053 n5912_145 vss 3.13114e-17
C9054 n5912_125 vss 3.13114e-17
C9055 n5912_124 vss 3.13114e-17
C9056 n5912_126 vss 1.40901e-17
C9057 n5912_125 vss 1.40901e-17
C9058 n5912_127 vss 3.91392e-17
C9059 n5912_144 vss 3.91392e-17
C9060 n5912_128 vss 1.40901e-17
C9061 n5912_127 vss 1.40901e-17
C9062 n5912_129 vss 1.20606e-16
C9063 n5912_151 vss 1.20606e-16
C9064 n5912_130 vss 2.92378e-17
C9065 n5912_129 vss 2.92378e-17
C9066 n5912_131 vss 2.92378e-17
C9067 n5912_130 vss 2.92378e-17
C9068 n5912_132 vss 2.92378e-17
C9069 n5912_131 vss 2.92378e-17
C9070 n5912_133 vss 2.92378e-17
C9071 n5912_132 vss 2.92378e-17
C9072 n5912_134 vss 2.92378e-17
C9073 n5912_133 vss 2.92378e-17
C9074 n5912_135 vss 2.92378e-17
C9075 n5912_134 vss 2.92378e-17
C9076 n5912_136 vss 2.92378e-17
C9077 n5912_135 vss 2.92378e-17
C9078 n5912_137 vss 2.92378e-17
C9079 n5912_136 vss 2.92378e-17
C9080 n5912_138 vss 2.92378e-17
C9081 n5912_137 vss 2.92378e-17
C9082 n5912_139 vss 2.92378e-17
C9083 n5912_138 vss 2.92378e-17
C9084 n5912_140 vss 2.92378e-17
C9085 n5912_139 vss 2.92378e-17
C9086 n5912_141 vss 2.92378e-17
C9087 n5912_140 vss 2.92378e-17
C9088 n5912_142 vss 2.92378e-17
C9089 n5912_141 vss 2.92378e-17
C9090 n5912_143 vss 2.92378e-17
C9091 n5912_142 vss 2.92378e-17
C9092 n5912_155 vss 1.20606e-16
C9093 n5912_150 vss 1.20606e-16
C9094 n5912_156 vss 2.92378e-17
C9095 n5912_155 vss 2.92378e-17
C9096 n5912_157 vss 2.92378e-17
C9097 n5912_156 vss 2.92378e-17
C9098 n5912_158 vss 2.92378e-17
C9099 n5912_157 vss 2.92378e-17
C9100 n5912_159 vss 2.92378e-17
C9101 n5912_158 vss 2.92378e-17
C9102 n5912_160 vss 2.92378e-17
C9103 n5912_159 vss 2.92378e-17
C9104 n5912_161 vss 2.92378e-17
C9105 n5912_160 vss 2.92378e-17
C9106 n5912_162 vss 2.92378e-17
C9107 n5912_161 vss 2.92378e-17
C9108 n5912_163 vss 2.92378e-17
C9109 n5912_162 vss 2.92378e-17
C9110 n5912_164 vss 2.92378e-17
C9111 n5912_163 vss 2.92378e-17
C9112 n5912_165 vss 2.92378e-17
C9113 n5912_164 vss 2.92378e-17
C9114 n5912_166 vss 2.92378e-17
C9115 n5912_165 vss 2.92378e-17
C9116 n5912_167 vss 2.92378e-17
C9117 n5912_166 vss 2.92378e-17
C9118 n5912_168 vss 2.92378e-17
C9119 n5912_167 vss 2.92378e-17
C9120 n5912_169 vss 2.92378e-17
C9121 n5912_168 vss 2.92378e-17
C9122 n5912_146 vss 7.94526e-16
C9123 n5912_144 vss 7.94526e-16
C9124 n5912_145 vss 8.96288e-16
C9125 n5912_146 vss 8.96288e-16
C9126 n5912_147 vss 1.33073e-16
C9127 n5912_146 vss 1.33073e-16
C9128 n5912_148 vss 1.87868e-16
C9129 n5912_147 vss 1.87868e-16
C9130 n5912_149 vss 1.87868e-16
C9131 n5912_148 vss 1.87868e-16
C9132 n5912_150 vss 1.95696e-16
C9133 n5912_149 vss 1.95696e-16
C9134 n5912_151 vss 1.01762e-16
C9135 n5912_150 vss 1.01762e-16
C9136 n5912_152 vss 7.82784e-17
C9137 n5912_151 vss 7.82784e-17
C9138 n5912_153 vss 1.87868e-16
C9139 n5912_152 vss 1.87868e-16
C9140 n5912_154 vss 1.40901e-17
C9141 n5912_153 vss 1.40901e-17
C9142 n5912_2 vss 2.34738e-17
C9143 n5912_1 vss 2.34738e-17
C9144 n5912_4 vss 2.34738e-17
C9145 n5912_2 vss 2.34738e-17
C9146 n5912_5 vss 4.69476e-17
C9147 n5912_4 vss 4.69476e-17
C9148 n5912_6 vss 4.69476e-17
C9149 n5912_5 vss 4.69476e-17
C9150 n5912_3 vss 7.33536e-17
C9151 n5912_2 vss 7.33536e-17

R160_1 ss_2_2 ss_2_5 0.001
R160_2 ss_2_6 ss_2_3 0.001
R160_3 ss_2_4 ss_2_10 0.001
R160_4 ss_2_8 ss_2_14 0.001
R160_5 ss_2_9 ss_2_7 0.001
R160_6 ss_2_12 ss_2_22 0.001
R160_7 ss_2_25 ss_2_29 0.001
R160_8 ss_2_20 ss_2_15 0.001
R160_9 ss_2_16 ss_2_18 0.001
R160_10 ss_2_28 ss_2_32 0.001
R160_11 ss_2_30 ss_2_40 0.001
R160_12 ss_2_38 ss_2_35 0.001
R160_13 ss_2_39 ss_2_35 0.001
R160_14 ss_2_37 ss_2_36 0.001
R160_15 ss_2_13 ss_2_11 0.001
R160_16 ss_2_37 ss_2_41 0.324
R160_17 ss_2_39 ss_2_38 0.216
R160_18 ss_2_40 ss_2_39 0.216
R160_19 ss_2_41 ss_2_40 0.108
R160_20 ss_2_18 ss_2_17 108
R160_21 ss_2 ss_2_18 50.4
R160_22 ss_2_30 ss_2_34 0.594
R160_23 ss_2_31 ss_2_30 0.54
R160_24 ss_2_33 ss_2_32 0.108
R160_25 ss_2_34 ss_2_33 0.054
R160_26 ss_2_16 ss_2_15 0.216
R160_27 ss_2_29 ss_2_28 18.576
R160_28 ss_2_20 ss_2_27 0.54
R160_29 ss_2_21 ss_2_20 0.54
R160_30 ss_2_25 ss_2_24 0.27
R160_31 ss_2_26 ss_2_25 0.108
R160_32 ss_2_27 ss_2_26 0.054
R160_33 ss_2_23 ss_2_22 0.216
R160_34 ss_2_24 ss_2_23 0.054
R160_35 ss_2_12 ss_2_11 27.648
R160_36 ss_2_14 ss_2_13 4.698
R160_37 ss_2_8 ss_2_7 5.724
R160_38 ss_2_10 ss_2_9 5.832
R160_39 ss_2_4 ss_2_6 0.324
R160_40 ss_2_6 ss_2_5 0.324
R160_41 ss_2_2 ss_2_1 475.2

C9152 ss_2_37 vss 4.07462e-17
C9153 ss_2_41 vss 4.07462e-17
C9154 ss_2_39 vss 4.38566e-17
C9155 ss_2_38 vss 4.38566e-17
C9156 ss_2_40 vss 4.38566e-17
C9157 ss_2_39 vss 4.38566e-17
C9158 ss_2_41 vss 3.65472e-17
C9159 ss_2_40 vss 3.65472e-17
C9160 ss_2_18 vss 1.21281e-16
C9161 ss_2_17 vss 1.21281e-16
C9162 ss_2 vss 5.86844e-17
C9163 ss_2_18 vss 5.86844e-17
C9164 ss_2_30 vss 1.35432e-16
C9165 ss_2_34 vss 1.35432e-16
C9166 ss_2_31 vss 1.2312e-16
C9167 ss_2_30 vss 1.2312e-16
C9168 ss_2_33 vss 3.078e-17
C9169 ss_2_32 vss 3.078e-17
C9170 ss_2_34 vss 1.2312e-17
C9171 ss_2_33 vss 1.2312e-17
C9172 ss_2_16 vss 2.71642e-17
C9173 ss_2_15 vss 2.71642e-17
C9174 ss_2_29 vss 1.87433e-15
C9175 ss_2_28 vss 1.87433e-15
C9176 ss_2_20 vss 1.29276e-16
C9177 ss_2_27 vss 1.29276e-16
C9178 ss_2_21 vss 1.29276e-16
C9179 ss_2_20 vss 1.29276e-16
C9180 ss_2_25 vss 6.156e-17
C9181 ss_2_24 vss 6.156e-17
C9182 ss_2_26 vss 3.078e-17
C9183 ss_2_25 vss 3.078e-17
C9184 ss_2_27 vss 1.2312e-17
C9185 ss_2_26 vss 1.2312e-17
C9186 ss_2_23 vss 5.5404e-17
C9187 ss_2_22 vss 5.5404e-17
C9188 ss_2_24 vss 1.2312e-17
C9189 ss_2_23 vss 1.2312e-17
C9190 ss_2_12 vss 2.78433e-15
C9191 ss_2_11 vss 2.78433e-15
C9192 ss_2_14 vss 1.0773e-15
C9193 ss_2_13 vss 1.0773e-15
C9194 ss_2_8 vss 1.02332e-15
C9195 ss_2_7 vss 1.02332e-15
C9196 ss_2_10 vss 1.33585e-15
C9197 ss_2_9 vss 1.33585e-15
C9198 ss_2_4 vss 7.30944e-17
C9199 ss_2_6 vss 7.30944e-17
C9200 ss_2_6 vss 7.30944e-17
C9201 ss_2_5 vss 7.30944e-17
C9202 ss_2_2 vss 5.18379e-16
C9203 ss_2_1 vss 5.18379e-16

R161_1 n5983_2 n5983_33 0.001
R161_2 n5983_20 n5983_6 0.001
R161_3 n5983_1 n5983_32 0.001
R161_4 n5983_29 n5983_5 0.001
R161_5 n5983_38 n5983_9 0.001
R161_6 n5983_39 n5983_9 0.001
R161_7 n5983_37 n5983_9 0.001
R161_8 n5983_36 n5983_9 0.001
R161_9 n5983_35 n5983_9 0.001
R161_10 n5983_27 n5983_10 0.001
R161_11 n5983_28 n5983_10 0.001
R161_12 n5983_26 n5983_10 0.001
R161_13 n5983_24 n5983_10 0.001
R161_14 n5983_25 n5983_12 0.001
R161_15 n5983_18 n5983_13 0.001
R161_16 n5983_17 n5983_13 0.001
R161_17 n5983_16 n5983_13 0.001
R161_18 n5983_11 n5983_15 0.001
R161_19 n5983_14 n5983_13 0.001
R161_20 n5983_6 n5983_5 7.2
R161_21 n5983_7 n5983_6 21.6
R161_22 n5983 n5983_7 0.001
R161_23 n5983_14 n5983_22 0.324
R161_24 n5983_15 n5983_14 0.108
R161_25 n5983_16 n5983_15 0.108
R161_26 n5983_17 n5983_16 0.108
R161_27 n5983_18 n5983_17 0.108
R161_28 n5983_19 n5983_18 0.001
R161_29 n5983_12 n5983_11 0.216
R161_30 n5983_20 n5983_29 0.108
R161_31 n5983_21 n5983_20 0.001
R161_32 n5983_23 n5983_22 0.324
R161_33 n5983_24 n5983_23 0.324
R161_34 n5983_25 n5983_24 0.108
R161_35 n5983_26 n5983_25 0.108
R161_36 n5983_27 n5983_26 0.108
R161_37 n5983_28 n5983_27 0.108
R161_38 n5983_29 n5983_28 0.108
R161_39 n5983_30 n5983_29 0.216
R161_40 n5983_31 n5983_30 0.108
R161_41 n5983_32 n5983_31 0.216
R161_42 n5983_35 n5983_32 0.108
R161_43 n5983_36 n5983_35 0.108
R161_44 n5983_37 n5983_36 0.108
R161_45 n5983_38 n5983_37 0.108
R161_46 n5983_39 n5983_38 0.108
R161_47 n5983_40 n5983_39 0.001
R161_48 n5983_33 n5983_32 0.108
R161_49 n5983_34 n5983_33 0.001
R161_50 n5983_2 n5983_1 7.2
R161_51 n5983_3 n5983_2 21.6
R161_52 n5983_4 n5983_3 0.001

C9204 n5983_6 vss 4.20552e-17
C9205 n5983_5 vss 4.20552e-17
C9206 n5983_7 vss 9.46242e-17
C9207 n5983_6 vss 9.46242e-17
C9208 n5983 vss 3.05111e-16
C9209 n5983_7 vss 3.05111e-16
C9210 n5983_14 vss 1.0959e-16
C9211 n5983_22 vss 1.0959e-16
C9212 n5983_15 vss 3.91392e-17
C9213 n5983_14 vss 3.91392e-17
C9214 n5983_16 vss 3.91392e-17
C9215 n5983_15 vss 3.91392e-17
C9216 n5983_17 vss 3.91392e-17
C9217 n5983_16 vss 3.91392e-17
C9218 n5983_18 vss 3.91392e-17
C9219 n5983_17 vss 3.91392e-17
C9220 n5983_19 vss 1.40901e-17
C9221 n5983_18 vss 1.40901e-17
C9222 n5983_12 vss 7.81488e-17
C9223 n5983_11 vss 7.81488e-17
C9224 n5983_20 vss 3.71822e-17
C9225 n5983_29 vss 3.71822e-17
C9226 n5983_21 vss 1.40901e-17
C9227 n5983_20 vss 1.40901e-17
C9228 n5983_23 vss 9.39341e-17
C9229 n5983_22 vss 9.39341e-17
C9230 n5983_24 vss 1.0959e-16
C9231 n5983_23 vss 1.0959e-16
C9232 n5983_25 vss 3.91392e-17
C9233 n5983_24 vss 3.91392e-17
C9234 n5983_26 vss 3.91392e-17
C9235 n5983_25 vss 3.91392e-17
C9236 n5983_27 vss 3.91392e-17
C9237 n5983_26 vss 3.91392e-17
C9238 n5983_28 vss 3.91392e-17
C9239 n5983_27 vss 3.91392e-17
C9240 n5983_29 vss 4.6967e-17
C9241 n5983_28 vss 4.6967e-17
C9242 n5983_30 vss 5.63604e-17
C9243 n5983_29 vss 5.63604e-17
C9244 n5983_31 vss 2.81802e-17
C9245 n5983_30 vss 2.81802e-17
C9246 n5983_32 vss 6.41883e-17
C9247 n5983_31 vss 6.41883e-17
C9248 n5983_35 vss 4.6967e-17
C9249 n5983_32 vss 4.6967e-17
C9250 n5983_36 vss 3.91392e-17
C9251 n5983_35 vss 3.91392e-17
C9252 n5983_37 vss 4.6967e-17
C9253 n5983_36 vss 4.6967e-17
C9254 n5983_38 vss 3.91392e-17
C9255 n5983_37 vss 3.91392e-17
C9256 n5983_39 vss 3.91392e-17
C9257 n5983_38 vss 3.91392e-17
C9258 n5983_40 vss 1.40901e-17
C9259 n5983_39 vss 1.40901e-17
C9260 n5983_33 vss 3.71822e-17
C9261 n5983_32 vss 3.71822e-17
C9262 n5983_34 vss 1.40901e-17
C9263 n5983_33 vss 1.40901e-17
C9264 n5983_2 vss 4.20552e-17
C9265 n5983_1 vss 4.20552e-17
C9266 n5983_3 vss 9.46242e-17
C9267 n5983_2 vss 9.46242e-17
C9268 n5983_4 vss 5.47139e-16
C9269 n5983_3 vss 5.47139e-16

R162_1 aa_0_1 aa_0_37 0.001
R162_2 aa_0_1 aa_0_35 0.001
R162_3 aa_0_1 aa_0_36 0.001
R162_4 aa_0_1 aa_0_34 0.001
R162_5 aa_0_1 aa_0_38 0.001
R162_6 aa_0_1 aa_0_39 0.001
R162_7 aa_0_1 aa_0_40 0.001
R162_8 aa_0_1 aa_0_41 0.001
R162_9 aa_0_1 aa_0_46 0.001
R162_10 aa_0_1 aa_0_45 0.001
R162_11 aa_0_1 aa_0_44 0.001
R162_12 aa_0_1 aa_0_43 0.001
R162_13 aa_0_1 aa_0_42 0.001
R162_14 aa_0_1 aa_0_33 0.001
R162_15 aa_0_29 aa_0_2 0.001
R162_16 aa_0_31 aa_0_2 0.001
R162_17 aa_0_32 aa_0_2 0.001
R162_18 aa_0_30 aa_0_2 0.001
R162_19 aa_0_28 aa_0_4 0.001
R162_20 aa_0_26 aa_0_7 0.001
R162_21 aa_0_6 aa_0_9 0.001
R162_22 aa_0_8 aa_0_10 0.001
R162_23 aa_0_11 aa_0_13 0.001
R162_24 aa_0_12 aa_0_25 0.001
R162_25 aa_0_20 aa_0_15 0.001
R162_26 aa_0_14 aa_0_17 0.001
R162_27 aa_0_17 aa_0_16 72
R162_28 aa_0 aa_0_17 43.2
R162_29 aa_0_15 aa_0_14 0.108
R162_30 aa_0_20 aa_0_19 0.756
R162_31 aa_0_21 aa_0_20 0.324
R162_32 aa_0_22 aa_0_21 0.054
R162_33 aa_0_23 aa_0_22 0.648
R162_34 aa_0_24 aa_0_23 0.054
R162_35 aa_0_25 aa_0_24 0.648
R162_36 aa_0_13 aa_0_12 9.936
R162_37 aa_0_11 aa_0_10 0.81
R162_38 aa_0_9 aa_0_8 9.072
R162_39 aa_0_7 aa_0_6 7.236
R162_40 aa_0_4 aa_0_3 0.054
R162_41 aa_0_5 aa_0_4 0.001
R162_42 aa_0_27 aa_0_26 0.54
R162_43 aa_0_28 aa_0_27 0.001
R162_44 aa_0_29 aa_0_28 0.54
R162_45 aa_0_30 aa_0_29 0.108
R162_46 aa_0_31 aa_0_30 0.108
R162_47 aa_0_32 aa_0_31 0.108
R162_48 aa_0_33 aa_0_32 0.864
R162_49 aa_0_34 aa_0_33 0.108
R162_50 aa_0_35 aa_0_34 0.108
R162_51 aa_0_36 aa_0_35 0.108
R162_52 aa_0_37 aa_0_36 0.108
R162_53 aa_0_38 aa_0_37 0.108
R162_54 aa_0_39 aa_0_38 0.108
R162_55 aa_0_40 aa_0_39 0.108
R162_56 aa_0_41 aa_0_40 0.108
R162_57 aa_0_42 aa_0_41 0.108
R162_58 aa_0_43 aa_0_42 0.108
R162_59 aa_0_44 aa_0_43 0.108
R162_60 aa_0_45 aa_0_44 0.108
R162_61 aa_0_46 aa_0_45 0.108
R162_62 aa_0_47 aa_0_46 0.001

C9270 aa_0_17 vss 8.21582e-17
C9271 aa_0_16 vss 8.21582e-17
C9272 aa_0 vss 5.086e-17
C9273 aa_0_17 vss 5.086e-17
C9274 aa_0_15 vss 3.65472e-17
C9275 aa_0_14 vss 3.65472e-17
C9276 aa_0_20 vss 1.78524e-16
C9277 aa_0_19 vss 1.78524e-16
C9278 aa_0_21 vss 8.0028e-17
C9279 aa_0_20 vss 8.0028e-17
C9280 aa_0_22 vss 1.2312e-17
C9281 aa_0_21 vss 1.2312e-17
C9282 aa_0_23 vss 1.539e-16
C9283 aa_0_22 vss 1.539e-16
C9284 aa_0_24 vss 1.2312e-17
C9285 aa_0_23 vss 1.2312e-17
C9286 aa_0_25 vss 1.47744e-16
C9287 aa_0_24 vss 1.47744e-16
C9288 aa_0_13 vss 1.00507e-15
C9289 aa_0_12 vss 1.00507e-15
C9290 aa_0_11 vss 1.8468e-16
C9291 aa_0_10 vss 1.8468e-16
C9292 aa_0_9 vss 9.1679e-16
C9293 aa_0_8 vss 9.1679e-16
C9294 aa_0_7 vss 1.64981e-15
C9295 aa_0_6 vss 1.64981e-15
C9296 aa_0_4 vss 1.95372e-17
C9297 aa_0_3 vss 1.95372e-17
C9298 aa_0_5 vss 1.30248e-17
C9299 aa_0_4 vss 1.30248e-17
C9300 aa_0_27 vss 6.24776e-17
C9301 aa_0_26 vss 6.24776e-17
C9302 aa_0_28 vss 2.1918e-17
C9303 aa_0_27 vss 2.1918e-17
C9304 aa_0_29 vss 1.64385e-16
C9305 aa_0_28 vss 1.64385e-16
C9306 aa_0_30 vss 3.91392e-17
C9307 aa_0_29 vss 3.91392e-17
C9308 aa_0_31 vss 3.91392e-17
C9309 aa_0_30 vss 3.91392e-17
C9310 aa_0_32 vss 3.91392e-17
C9311 aa_0_31 vss 3.91392e-17
C9312 aa_0_33 vss 2.42663e-16
C9313 aa_0_32 vss 2.42663e-16
C9314 aa_0_34 vss 3.13114e-17
C9315 aa_0_33 vss 3.13114e-17
C9316 aa_0_35 vss 3.13114e-17
C9317 aa_0_34 vss 3.13114e-17
C9318 aa_0_36 vss 3.13114e-17
C9319 aa_0_35 vss 3.13114e-17
C9320 aa_0_37 vss 3.13114e-17
C9321 aa_0_36 vss 3.13114e-17
C9322 aa_0_38 vss 3.13114e-17
C9323 aa_0_37 vss 3.13114e-17
C9324 aa_0_39 vss 3.13114e-17
C9325 aa_0_38 vss 3.13114e-17
C9326 aa_0_40 vss 3.13114e-17
C9327 aa_0_39 vss 3.13114e-17
C9328 aa_0_41 vss 3.13114e-17
C9329 aa_0_40 vss 3.13114e-17
C9330 aa_0_42 vss 3.13114e-17
C9331 aa_0_41 vss 3.13114e-17
C9332 aa_0_43 vss 3.13114e-17
C9333 aa_0_42 vss 3.13114e-17
C9334 aa_0_44 vss 3.13114e-17
C9335 aa_0_43 vss 3.13114e-17
C9336 aa_0_45 vss 3.13114e-17
C9337 aa_0_44 vss 3.13114e-17
C9338 aa_0_46 vss 3.13114e-17
C9339 aa_0_45 vss 3.13114e-17
C9340 aa_0_47 vss 1.40901e-17
C9341 aa_0_46 vss 1.40901e-17

R5_1 a_0_50 a_0_1 0.001
R5_2 a_0_48 a_0_1 0.001
R5_3 a_0_49 a_0_1 0.001
R5_4 a_0_47 a_0_1 0.001
R5_5 a_0_46 a_0_1 0.001
R5_6 a_0_45 a_0_1 0.001
R5_7 a_0_44 a_0_1 0.001
R5_8 a_0_43 a_0_1 0.001
R5_9 a_0_41 a_0_2 0.001
R5_10 a_0_42 a_0_2 0.001
R5_11 a_0_39 a_0_2 0.001
R5_12 a_0_40 a_0_2 0.001
R5_13 a_0_36 a_0_2 0.001
R5_14 a_0_37 a_0_2 0.001
R5_15 a_0_38 a_0_2 0.001
R5_16 a_0_35 a_0_2 0.001
R5_17 a_0_34 a_0_2 0.001
R5_18 a_0_33 a_0_2 0.001
R5_19 a_0_32 a_0_2 0.001
R5_20 a_0_30 a_0_2 0.001
R5_21 a_0_31 a_0_2 0.001
R5_22 a_0_28 a_0_2 0.001
R5_23 a_0_29 a_0_2 0.001
R5_24 a_0_27 a_0_2 0.001
R5_25 a_0_26 a_0_2 0.001
R5_26 a_0_24 a_0_2 0.001
R5_27 a_0_25 a_0_2 0.001
R5_28 a_0_23 a_0_2 0.001
R5_29 a_0_79 a_0_3 0.001
R5_30 a_0_77 a_0_3 0.001
R5_31 a_0_78 a_0_3 0.001
R5_32 a_0_76 a_0_3 0.001
R5_33 a_0_75 a_0_3 0.001
R5_34 a_0_73 a_0_3 0.001
R5_35 a_0_74 a_0_3 0.001
R5_36 a_0_72 a_0_3 0.001
R5_37 a_0_70 a_0_4 0.001
R5_38 a_0_71 a_0_4 0.001
R5_39 a_0_68 a_0_4 0.001
R5_40 a_0_69 a_0_4 0.001
R5_41 a_0_66 a_0_4 0.001
R5_42 a_0_65 a_0_4 0.001
R5_43 a_0_67 a_0_4 0.001
R5_44 a_0_63 a_0_4 0.001
R5_45 a_0_64 a_0_4 0.001
R5_46 a_0_62 a_0_4 0.001
R5_47 a_0_61 a_0_4 0.001
R5_48 a_0_59 a_0_4 0.001
R5_49 a_0_60 a_0_4 0.001
R5_50 a_0_58 a_0_4 0.001
R5_51 a_0_57 a_0_4 0.001
R5_52 a_0_55 a_0_4 0.001
R5_53 a_0_56 a_0_4 0.001
R5_54 a_0_54 a_0_4 0.001
R5_55 a_0_53 a_0_4 0.001
R5_56 a_0_52 a_0_4 0.001
R5_57 a_0_14 a_0_5 0.001
R5_58 a_0_13 a_0_8 0.001
R5_59 a_0 a_0_11 0.001
R5_60 a_0_6 a_0_5 21.6
R5_61 a_0_8 a_0_7 7.2
R5_62 a_0_9 a_0_8 7.2
R5_63 a_0_10 a_0_9 14.4
R5_64 a_0_13 a_0_12 0.001
R5_65 a_0_16 a_0_13 0.216
R5_66 a_0_14 a_0_16 0.216
R5_67 a_0_15 a_0_14 0.001
R5_68 a_0_16 a_0_17 0.324
R5_69 a_0_18 a_0_17 2.268
R5_70 a_0_19 a_0_18 1.08
R5_71 a_0_20 a_0_19 0.001
R5_72 a_0_21 a_0_20 0.001
R5_73 a_0_51 a_0_21 0.216
R5_74 a_0_23 a_0_22 0.001
R5_75 a_0_24 a_0_23 0.108
R5_76 a_0_25 a_0_24 0.108
R5_77 a_0_26 a_0_25 0.108
R5_78 a_0_27 a_0_26 0.108
R5_79 a_0_28 a_0_27 0.108
R5_80 a_0_29 a_0_28 0.108
R5_81 a_0_30 a_0_29 0.108
R5_82 a_0_31 a_0_30 0.108
R5_83 a_0_32 a_0_31 0.108
R5_84 a_0_33 a_0_32 0.108
R5_85 a_0_34 a_0_33 0.108
R5_86 a_0_35 a_0_34 0.108
R5_87 a_0_36 a_0_35 0.108
R5_88 a_0_37 a_0_36 0.108
R5_89 a_0_38 a_0_37 0.108
R5_90 a_0_39 a_0_38 0.108
R5_91 a_0_40 a_0_39 0.108
R5_92 a_0_41 a_0_40 0.108
R5_93 a_0_42 a_0_41 0.108
R5_94 a_0_43 a_0_42 0.864
R5_95 a_0_44 a_0_43 0.108
R5_96 a_0_45 a_0_44 0.108
R5_97 a_0_46 a_0_45 0.108
R5_98 a_0_47 a_0_46 0.108
R5_99 a_0_48 a_0_47 0.108
R5_100 a_0_49 a_0_48 0.108
R5_101 a_0_50 a_0_49 0.108
R5_102 a_0_81 a_0_50 0.54
R5_103 a_0_52 a_0_51 0.001
R5_104 a_0_53 a_0_52 0.108
R5_105 a_0_54 a_0_53 0.108
R5_106 a_0_55 a_0_54 0.108
R5_107 a_0_56 a_0_55 0.108
R5_108 a_0_57 a_0_56 0.108
R5_109 a_0_58 a_0_57 0.108
R5_110 a_0_59 a_0_58 0.108
R5_111 a_0_60 a_0_59 0.108
R5_112 a_0_61 a_0_60 0.108
R5_113 a_0_62 a_0_61 0.108
R5_114 a_0_63 a_0_62 0.108
R5_115 a_0_64 a_0_63 0.108
R5_116 a_0_65 a_0_64 0.108
R5_117 a_0_66 a_0_65 0.108
R5_118 a_0_67 a_0_66 0.108
R5_119 a_0_68 a_0_67 0.108
R5_120 a_0_69 a_0_68 0.108
R5_121 a_0_70 a_0_69 0.108
R5_122 a_0_71 a_0_70 0.108
R5_123 a_0_72 a_0_71 0.864
R5_124 a_0_73 a_0_72 0.108
R5_125 a_0_74 a_0_73 0.108
R5_126 a_0_75 a_0_74 0.108
R5_127 a_0_76 a_0_75 0.108
R5_128 a_0_77 a_0_76 0.108
R5_129 a_0_78 a_0_77 0.108
R5_130 a_0_79 a_0_78 0.108
R5_131 a_0_82 a_0_79 0.54
R5_132 a_0_82 a_0_80 0.001
R5_133 a_0_81 a_0_82 0.108
R5_134 a_0_83 a_0_82 0.54
R5_135 a_0_84 a_0_83 0.001
R5_136 a_0 a_0_84 0.001

C9342 a_0_6 vss 9.46242e-17
C9343 a_0_5 vss 9.46242e-17
C9344 a_0_8 vss 3.15414e-17
C9345 a_0_7 vss 3.15414e-17
C9346 a_0_9 vss 3.15414e-17
C9347 a_0_8 vss 3.15414e-17
C9348 a_0_10 vss 6.30828e-17
C9349 a_0_9 vss 6.30828e-17
C9350 a_0_13 vss 1.40901e-17
C9351 a_0_12 vss 1.40901e-17
C9352 a_0_16 vss 7.82784e-17
C9353 a_0_13 vss 7.82784e-17
C9354 a_0_14 vss 7.04506e-17
C9355 a_0_16 vss 7.04506e-17
C9356 a_0_15 vss 1.40901e-17
C9357 a_0_14 vss 1.40901e-17
C9358 a_0_16 vss 9.39341e-17
C9359 a_0_17 vss 9.39341e-17
C9360 a_0_18 vss 6.18399e-16
C9361 a_0_17 vss 6.18399e-16
C9362 a_0_19 vss 2.97458e-16
C9363 a_0_18 vss 2.97458e-16
C9364 a_0_20 vss 2.50491e-17
C9365 a_0_19 vss 2.50491e-17
C9366 a_0_21 vss 1.25245e-17
C9367 a_0_20 vss 1.25245e-17
C9368 a_0_51 vss 8.14095e-17
C9369 a_0_21 vss 8.14095e-17
C9370 a_0_23 vss 1.40901e-17
C9371 a_0_22 vss 1.40901e-17
C9372 a_0_24 vss 3.13114e-17
C9373 a_0_23 vss 3.13114e-17
C9374 a_0_25 vss 3.13114e-17
C9375 a_0_24 vss 3.13114e-17
C9376 a_0_26 vss 3.13114e-17
C9377 a_0_25 vss 3.13114e-17
C9378 a_0_27 vss 3.13114e-17
C9379 a_0_26 vss 3.13114e-17
C9380 a_0_28 vss 3.13114e-17
C9381 a_0_27 vss 3.13114e-17
C9382 a_0_29 vss 3.13114e-17
C9383 a_0_28 vss 3.13114e-17
C9384 a_0_30 vss 3.13114e-17
C9385 a_0_29 vss 3.13114e-17
C9386 a_0_31 vss 3.13114e-17
C9387 a_0_30 vss 3.13114e-17
C9388 a_0_32 vss 3.13114e-17
C9389 a_0_31 vss 3.13114e-17
C9390 a_0_33 vss 3.13114e-17
C9391 a_0_32 vss 3.13114e-17
C9392 a_0_34 vss 3.13114e-17
C9393 a_0_33 vss 3.13114e-17
C9394 a_0_35 vss 3.13114e-17
C9395 a_0_34 vss 3.13114e-17
C9396 a_0_36 vss 3.13114e-17
C9397 a_0_35 vss 3.13114e-17
C9398 a_0_37 vss 3.13114e-17
C9399 a_0_36 vss 3.13114e-17
C9400 a_0_38 vss 3.13114e-17
C9401 a_0_37 vss 3.13114e-17
C9402 a_0_39 vss 3.13114e-17
C9403 a_0_38 vss 3.13114e-17
C9404 a_0_40 vss 3.13114e-17
C9405 a_0_39 vss 3.13114e-17
C9406 a_0_41 vss 3.13114e-17
C9407 a_0_40 vss 3.13114e-17
C9408 a_0_42 vss 3.13114e-17
C9409 a_0_41 vss 3.13114e-17
C9410 a_0_43 vss 2.42663e-16
C9411 a_0_42 vss 2.42663e-16
C9412 a_0_44 vss 3.13114e-17
C9413 a_0_43 vss 3.13114e-17
C9414 a_0_45 vss 3.13114e-17
C9415 a_0_44 vss 3.13114e-17
C9416 a_0_46 vss 3.13114e-17
C9417 a_0_45 vss 3.13114e-17
C9418 a_0_47 vss 3.13114e-17
C9419 a_0_46 vss 3.13114e-17
C9420 a_0_48 vss 3.13114e-17
C9421 a_0_47 vss 3.13114e-17
C9422 a_0_49 vss 3.13114e-17
C9423 a_0_48 vss 3.13114e-17
C9424 a_0_50 vss 3.13114e-17
C9425 a_0_49 vss 3.13114e-17
C9426 a_0_81 vss 1.40901e-16
C9427 a_0_50 vss 1.40901e-16
C9428 a_0_52 vss 1.40901e-17
C9429 a_0_51 vss 1.40901e-17
C9430 a_0_53 vss 3.13114e-17
C9431 a_0_52 vss 3.13114e-17
C9432 a_0_54 vss 3.13114e-17
C9433 a_0_53 vss 3.13114e-17
C9434 a_0_55 vss 3.13114e-17
C9435 a_0_54 vss 3.13114e-17
C9436 a_0_56 vss 3.13114e-17
C9437 a_0_55 vss 3.13114e-17
C9438 a_0_57 vss 3.13114e-17
C9439 a_0_56 vss 3.13114e-17
C9440 a_0_58 vss 3.13114e-17
C9441 a_0_57 vss 3.13114e-17
C9442 a_0_59 vss 3.13114e-17
C9443 a_0_58 vss 3.13114e-17
C9444 a_0_60 vss 3.13114e-17
C9445 a_0_59 vss 3.13114e-17
C9446 a_0_61 vss 3.13114e-17
C9447 a_0_60 vss 3.13114e-17
C9448 a_0_62 vss 3.13114e-17
C9449 a_0_61 vss 3.13114e-17
C9450 a_0_63 vss 3.13114e-17
C9451 a_0_62 vss 3.13114e-17
C9452 a_0_64 vss 3.13114e-17
C9453 a_0_63 vss 3.13114e-17
C9454 a_0_65 vss 3.13114e-17
C9455 a_0_64 vss 3.13114e-17
C9456 a_0_66 vss 3.13114e-17
C9457 a_0_65 vss 3.13114e-17
C9458 a_0_67 vss 3.13114e-17
C9459 a_0_66 vss 3.13114e-17
C9460 a_0_68 vss 3.13114e-17
C9461 a_0_67 vss 3.13114e-17
C9462 a_0_69 vss 3.13114e-17
C9463 a_0_68 vss 3.13114e-17
C9464 a_0_70 vss 3.13114e-17
C9465 a_0_69 vss 3.13114e-17
C9466 a_0_71 vss 3.13114e-17
C9467 a_0_70 vss 3.13114e-17
C9468 a_0_72 vss 2.42663e-16
C9469 a_0_71 vss 2.42663e-16
C9470 a_0_73 vss 3.13114e-17
C9471 a_0_72 vss 3.13114e-17
C9472 a_0_74 vss 3.13114e-17
C9473 a_0_73 vss 3.13114e-17
C9474 a_0_75 vss 3.13114e-17
C9475 a_0_74 vss 3.13114e-17
C9476 a_0_76 vss 3.13114e-17
C9477 a_0_75 vss 3.13114e-17
C9478 a_0_77 vss 3.13114e-17
C9479 a_0_76 vss 3.13114e-17
C9480 a_0_78 vss 3.13114e-17
C9481 a_0_77 vss 3.13114e-17
C9482 a_0_79 vss 3.13114e-17
C9483 a_0_78 vss 3.13114e-17
C9484 a_0_82 vss 1.40901e-16
C9485 a_0_79 vss 1.40901e-16
C9486 a_0_82 vss 6.34418e-17
C9487 a_0_80 vss 6.34418e-17
C9488 a_0_81 vss 1.42197e-16
C9489 a_0_82 vss 1.42197e-16
C9490 a_0_83 vss 6.8969e-16
C9491 a_0_82 vss 6.8969e-16
C9492 a_0_84 vss 3.48676e-17
C9493 a_0_83 vss 3.48676e-17
C9494 a_0 vss 4.3846e-15
C9495 a_0_84 vss 4.3846e-15

R163_1 clock_1 clock_53 0.001
R163_2 clock_1 clock_52 0.001
R163_3 clock_1 clock_51 0.001
R163_4 clock_1 clock_54 0.001
R163_5 clock_1 clock_57 0.001
R163_6 clock_1 clock_56 0.001
R163_7 clock_1 clock_55 0.001
R163_8 clock_1 clock_58 0.001
R163_9 clock_48 clock_2 0.001
R163_10 clock_41 clock_2 0.001
R163_11 clock_42 clock_2 0.001
R163_12 clock_43 clock_2 0.001
R163_13 clock_44 clock_2 0.001
R163_14 clock_45 clock_2 0.001
R163_15 clock_46 clock_2 0.001
R163_16 clock_47 clock_2 0.001
R163_17 clock_50 clock_3 0.001
R163_18 clock_27 clock_3 0.001
R163_19 clock_28 clock_3 0.001
R163_20 clock_29 clock_3 0.001
R163_21 clock_30 clock_3 0.001
R163_22 clock_31 clock_3 0.001
R163_23 clock_32 clock_3 0.001
R163_24 clock_33 clock_3 0.001
R163_25 clock_40 clock_4 0.001
R163_26 clock_36 clock_4 0.001
R163_27 clock_37 clock_4 0.001
R163_28 clock_38 clock_4 0.001
R163_29 clock_39 clock_4 0.001
R163_30 clock_23 clock_5 0.001
R163_31 clock_24 clock_5 0.001
R163_32 clock_20 clock_5 0.001
R163_33 clock_21 clock_5 0.001
R163_34 clock_22 clock_5 0.001
R163_35 clock_14 clock_6 0.001
R163_36 clock_15 clock_6 0.001
R163_37 clock_18 clock_6 0.001
R163_38 clock_17 clock_6 0.001
R163_39 clock_16 clock_6 0.001
R163_40 clock_8 clock_62 0.001
R163_41 clock_34 clock_10 0.001
R163_42 clock_9 clock_7 0.001
R163_43 clock_19 clock_11 0.001
R163_44 clock_13 clock_12 0.001
R163_45 clock_60 clock_91 0.001
R163_46 clock_61 clock_59 0.001
R163_47 clock_118 clock_70 0.001
R163_48 clock_71 clock_64 0.001
R163_49 clock_69 clock_67 0.001
R163_50 clock_82 clock_99 0.001
R163_51 clock_86 clock_79 0.001
R163_52 clock_83 clock_81 0.001
R163_53 clock_80 clock_73 0.001
R163_54 clock_78 clock_76 0.001
R163_55 clock_93 clock_124 0.001
R163_56 clock_121 clock_116 0.001
R163_57 clock_117 clock_110 0.001
R163_58 clock_115 clock_113 0.001
R163_59 clock_98 clock_92 0.001
R163_60 clock_95 clock_107 0.001
R163_61 clock_108 clock_101 0.001
R163_62 clock_106 clock_104 0.001
R163_63 clock_67 clock_66 86.4
R163_64 clock clock_67 100.8
R163_65 clock_63 clock_65 79.2
R163_66 clock_113 clock_112 86.4
R163_67 clock_114 clock_113 100.8
R163_68 clock_109 clock_111 79.2
R163_69 clock_65 clock_64 36
R163_70 clock_111 clock_110 36
R163_71 clock_70 clock_69 0.216
R163_72 clock_116 clock_115 0.216
R163_73 clock_71 clock_70 0.648
R163_74 clock_117 clock_116 0.648
R163_75 clock_104 clock_103 86.4
R163_76 clock_105 clock_104 100.8
R163_77 clock_100 clock_102 79.2
R163_78 clock_102 clock_101 36
R163_79 clock_118 clock_126 0.594
R163_80 clock_119 clock_118 0.54
R163_81 clock_121 clock_120 0.648
R163_82 clock_122 clock_121 0.486
R163_83 clock_107 clock_106 0.216
R163_84 clock_123 clock_122 0.054
R163_85 clock_124 clock_123 0.108
R163_86 clock_125 clock_124 0.918
R163_87 clock_126 clock_125 0.054
R163_88 clock_108 clock_107 0.648
R163_89 clock_93 clock_92 9.72
R163_90 clock_95 clock_94 0.648
R163_91 clock_96 clock_95 0.486
R163_92 clock_97 clock_96 0.054
R163_93 clock_98 clock_97 0.108
R163_94 clock_99 clock_98 0.81
R163_95 clock_76 clock_75 86.4
R163_96 clock_77 clock_76 100.8
R163_97 clock_72 clock_74 79.2
R163_98 clock_74 clock_73 36
R163_99 clock_82 clock_81 19.764
R163_100 clock_79 clock_78 0.216
R163_101 clock_80 clock_79 0.648
R163_102 clock_84 clock_83 0.108
R163_103 clock_85 clock_84 0.054
R163_104 clock_86 clock_85 0.594
R163_105 clock_87 clock_86 0.486
R163_106 clock_88 clock_87 0.054
R163_107 clock_89 clock_88 0.648
R163_108 clock_90 clock_89 0.054
R163_109 clock_91 clock_90 0.486
R163_110 clock_60 clock_59 5.4
R163_111 clock_62 clock_61 8.478
R163_112 clock_8 clock_7 3.24
R163_113 clock_25 clock_13 0.864
R163_114 clock_14 clock_25 0.432
R163_115 clock_15 clock_14 0.108
R163_116 clock_16 clock_15 0.108
R163_117 clock_17 clock_16 0.108
R163_118 clock_18 clock_17 0.108
R163_119 clock_26 clock_19 0.864
R163_120 clock_20 clock_26 0.432
R163_121 clock_21 clock_20 0.108
R163_122 clock_22 clock_21 0.108
R163_123 clock_23 clock_22 0.108
R163_124 clock_24 clock_23 0.108
R163_125 clock_10 clock_9 0.27
R163_126 clock_25 clock_35 0.432
R163_127 clock_26 clock_25 0.432
R163_128 clock_27 clock_50 0.108
R163_129 clock_28 clock_27 0.108
R163_130 clock_29 clock_28 0.108
R163_131 clock_30 clock_29 0.108
R163_132 clock_31 clock_30 0.108
R163_133 clock_32 clock_31 0.108
R163_134 clock_33 clock_32 0.108
R163_135 clock_35 clock_34 0.864
R163_136 clock_36 clock_35 0.432
R163_137 clock_37 clock_36 0.108
R163_138 clock_38 clock_37 0.108
R163_139 clock_39 clock_38 0.108
R163_140 clock_40 clock_39 0.108
R163_141 clock_48 clock_40 0.864
R163_142 clock_41 clock_48 0.108
R163_143 clock_42 clock_41 0.108
R163_144 clock_43 clock_42 0.108
R163_145 clock_44 clock_43 0.108
R163_146 clock_45 clock_44 0.108
R163_147 clock_46 clock_45 0.108
R163_148 clock_47 clock_46 0.108
R163_149 clock_51 clock_48 0.432
R163_150 clock_50 clock_51 0.432
R163_151 clock_50 clock_49 0.001
R163_152 clock_52 clock_51 0.108
R163_153 clock_53 clock_52 0.108
R163_154 clock_54 clock_53 0.108
R163_155 clock_55 clock_54 0.108
R163_156 clock_56 clock_55 0.108
R163_157 clock_57 clock_56 0.108
R163_158 clock_58 clock_57 0.108

C9496 clock_67 vss 9.78074e-17
C9497 clock_66 vss 9.78074e-17
C9498 clock vss 1.09544e-16
C9499 clock_67 vss 1.09544e-16
C9500 clock_63 vss 8.9983e-17
C9501 clock_65 vss 8.9983e-17
C9502 clock_113 vss 9.78074e-17
C9503 clock_112 vss 9.78074e-17
C9504 clock_114 vss 1.09544e-16
C9505 clock_113 vss 1.09544e-16
C9506 clock_109 vss 8.9983e-17
C9507 clock_111 vss 8.9983e-17
C9508 clock_65 vss 3.9123e-17
C9509 clock_64 vss 3.9123e-17
C9510 clock_111 vss 3.9123e-17
C9511 clock_110 vss 3.9123e-17
C9512 clock_70 vss 2.54664e-17
C9513 clock_69 vss 2.54664e-17
C9514 clock_116 vss 2.54664e-17
C9515 clock_115 vss 2.54664e-17
C9516 clock_71 vss 7.30037e-17
C9517 clock_70 vss 7.30037e-17
C9518 clock_117 vss 7.30037e-17
C9519 clock_116 vss 7.30037e-17
C9520 clock_104 vss 9.78074e-17
C9521 clock_103 vss 9.78074e-17
C9522 clock_105 vss 1.09544e-16
C9523 clock_104 vss 1.09544e-16
C9524 clock_100 vss 8.9983e-17
C9525 clock_102 vss 8.9983e-17
C9526 clock_102 vss 3.9123e-17
C9527 clock_101 vss 3.9123e-17
C9528 clock_118 vss 1.35432e-16
C9529 clock_126 vss 1.35432e-16
C9530 clock_119 vss 1.2312e-16
C9531 clock_118 vss 1.2312e-16
C9532 clock_121 vss 1.47744e-16
C9533 clock_120 vss 1.47744e-16
C9534 clock_122 vss 1.10808e-16
C9535 clock_121 vss 1.10808e-16
C9536 clock_107 vss 2.54664e-17
C9537 clock_106 vss 2.54664e-17
C9538 clock_123 vss 1.2312e-17
C9539 clock_122 vss 1.2312e-17
C9540 clock_124 vss 3.078e-17
C9541 clock_123 vss 3.078e-17
C9542 clock_125 vss 2.1546e-16
C9543 clock_124 vss 2.1546e-16
C9544 clock_126 vss 1.2312e-17
C9545 clock_125 vss 1.2312e-17
C9546 clock_108 vss 7.30037e-17
C9547 clock_107 vss 7.30037e-17
C9548 clock_93 vss 9.7791e-16
C9549 clock_92 vss 9.7791e-16
C9550 clock_95 vss 1.47744e-16
C9551 clock_94 vss 1.47744e-16
C9552 clock_96 vss 1.10808e-16
C9553 clock_95 vss 1.10808e-16
C9554 clock_97 vss 1.2312e-17
C9555 clock_96 vss 1.2312e-17
C9556 clock_98 vss 3.078e-17
C9557 clock_97 vss 3.078e-17
C9558 clock_99 vss 1.8468e-16
C9559 clock_98 vss 1.8468e-16
C9560 clock_76 vss 9.78074e-17
C9561 clock_75 vss 9.78074e-17
C9562 clock_77 vss 1.09544e-16
C9563 clock_76 vss 1.09544e-16
C9564 clock_72 vss 8.9983e-17
C9565 clock_74 vss 8.9983e-17
C9566 clock_74 vss 3.9123e-17
C9567 clock_73 vss 3.9123e-17
C9568 clock_82 vss 1.99657e-15
C9569 clock_81 vss 1.99657e-15
C9570 clock_79 vss 2.54664e-17
C9571 clock_78 vss 2.54664e-17
C9572 clock_80 vss 7.30037e-17
C9573 clock_79 vss 7.30037e-17
C9574 clock_84 vss 3.078e-17
C9575 clock_83 vss 3.078e-17
C9576 clock_85 vss 1.2312e-17
C9577 clock_84 vss 1.2312e-17
C9578 clock_86 vss 1.35432e-16
C9579 clock_85 vss 1.35432e-16
C9580 clock_87 vss 1.10808e-16
C9581 clock_86 vss 1.10808e-16
C9582 clock_88 vss 1.2312e-17
C9583 clock_87 vss 1.2312e-17
C9584 clock_89 vss 1.539e-16
C9585 clock_88 vss 1.539e-16
C9586 clock_90 vss 1.2312e-17
C9587 clock_89 vss 1.2312e-17
C9588 clock_91 vss 1.16964e-16
C9589 clock_90 vss 1.16964e-16
C9590 clock_60 vss 5.50074e-16
C9591 clock_59 vss 5.50074e-16
C9592 clock_62 vss 1.93914e-15
C9593 clock_61 vss 1.93914e-15
C9594 clock_8 vss 5.77446e-16
C9595 clock_7 vss 5.77446e-16
C9596 clock_25 vss 1.68117e-16
C9597 clock_13 vss 1.68117e-16
C9598 clock_14 vss 8.77133e-17
C9599 clock_25 vss 8.77133e-17
C9600 clock_15 vss 2.92378e-17
C9601 clock_14 vss 2.92378e-17
C9602 clock_16 vss 2.92378e-17
C9603 clock_15 vss 2.92378e-17
C9604 clock_17 vss 2.92378e-17
C9605 clock_16 vss 2.92378e-17
C9606 clock_18 vss 2.92378e-17
C9607 clock_17 vss 2.92378e-17
C9608 clock_26 vss 1.68117e-16
C9609 clock_19 vss 1.68117e-16
C9610 clock_20 vss 8.77133e-17
C9611 clock_26 vss 8.77133e-17
C9612 clock_21 vss 2.92378e-17
C9613 clock_20 vss 2.92378e-17
C9614 clock_22 vss 2.92378e-17
C9615 clock_21 vss 2.92378e-17
C9616 clock_23 vss 2.92378e-17
C9617 clock_22 vss 2.92378e-17
C9618 clock_24 vss 2.92378e-17
C9619 clock_23 vss 2.92378e-17
C9620 clock_10 vss 6.156e-17
C9621 clock_9 vss 6.156e-17
C9622 clock_25 vss 8.77133e-17
C9623 clock_35 vss 8.77133e-17
C9624 clock_26 vss 8.77133e-17
C9625 clock_25 vss 8.77133e-17
C9626 clock_27 vss 3.65472e-17
C9627 clock_50 vss 3.65472e-17
C9628 clock_28 vss 2.92378e-17
C9629 clock_27 vss 2.92378e-17
C9630 clock_29 vss 2.92378e-17
C9631 clock_28 vss 2.92378e-17
C9632 clock_30 vss 2.92378e-17
C9633 clock_29 vss 2.92378e-17
C9634 clock_31 vss 2.92378e-17
C9635 clock_30 vss 2.92378e-17
C9636 clock_32 vss 2.92378e-17
C9637 clock_31 vss 2.92378e-17
C9638 clock_33 vss 2.92378e-17
C9639 clock_32 vss 2.92378e-17
C9640 clock_35 vss 1.68117e-16
C9641 clock_34 vss 1.68117e-16
C9642 clock_36 vss 8.77133e-17
C9643 clock_35 vss 8.77133e-17
C9644 clock_37 vss 2.92378e-17
C9645 clock_36 vss 2.92378e-17
C9646 clock_38 vss 2.92378e-17
C9647 clock_37 vss 2.92378e-17
C9648 clock_39 vss 2.92378e-17
C9649 clock_38 vss 2.92378e-17
C9650 clock_40 vss 2.92378e-17
C9651 clock_39 vss 2.92378e-17
C9652 clock_48 vss 1.68117e-16
C9653 clock_40 vss 1.68117e-16
C9654 clock_41 vss 3.65472e-17
C9655 clock_48 vss 3.65472e-17
C9656 clock_42 vss 2.92378e-17
C9657 clock_41 vss 2.92378e-17
C9658 clock_43 vss 2.92378e-17
C9659 clock_42 vss 2.92378e-17
C9660 clock_44 vss 2.92378e-17
C9661 clock_43 vss 2.92378e-17
C9662 clock_45 vss 2.92378e-17
C9663 clock_44 vss 2.92378e-17
C9664 clock_46 vss 2.92378e-17
C9665 clock_45 vss 2.92378e-17
C9666 clock_47 vss 2.92378e-17
C9667 clock_46 vss 2.92378e-17
C9668 clock_51 vss 8.77133e-17
C9669 clock_48 vss 8.77133e-17
C9670 clock_50 vss 8.77133e-17
C9671 clock_51 vss 8.77133e-17
C9672 clock_50 vss 1.3157e-17
C9673 clock_49 vss 1.3157e-17
C9674 clock_52 vss 3.65472e-17
C9675 clock_51 vss 3.65472e-17
C9676 clock_53 vss 2.92378e-17
C9677 clock_52 vss 2.92378e-17
C9678 clock_54 vss 2.92378e-17
C9679 clock_53 vss 2.92378e-17
C9680 clock_55 vss 2.92378e-17
C9681 clock_54 vss 2.92378e-17
C9682 clock_56 vss 2.92378e-17
C9683 clock_55 vss 2.92378e-17
C9684 clock_57 vss 2.92378e-17
C9685 clock_56 vss 2.92378e-17
C9686 clock_58 vss 2.92378e-17
C9687 clock_57 vss 2.92378e-17

R164_1 p17_logic_ck_2 p17_logic_ck_9 0.001
R164_2 p17_logic_ck_7 p17_logic_ck_159 0.001
R164_3 p17_logic_ck_5 p17_logic_ck_159 0.001
R164_4 p17_logic_ck_6 p17_logic_ck_159 0.001
R164_5 p17_logic_ck_137 p17_logic_ck_80 0.001
R164_6 p17_logic_ck_136 p17_logic_ck_56 0.001
R164_7 p17_logic_ck_135 p17_logic_ck_32 0.001
R164_8 p17_logic_ck_135 p17_logic_ck_33 0.001
R164_9 p17_logic_ck_136 p17_logic_ck_57 0.001
R164_10 p17_logic_ck_137 p17_logic_ck_81 0.001
R164_11 p17_logic_ck_138 p17_logic_ck_104 0.001
R164_12 p17_logic_ck_138 p17_logic_ck_105 0.001
R164_13 p17_logic_ck_79 p17_logic_ck_59 0.001
R164_14 p17_logic_ck_78 p17_logic_ck_59 0.001
R164_15 p17_logic_ck_77 p17_logic_ck_59 0.001
R164_16 p17_logic_ck_55 p17_logic_ck_35 0.001
R164_17 p17_logic_ck_54 p17_logic_ck_35 0.001
R164_18 p17_logic_ck_53 p17_logic_ck_35 0.001
R164_19 p17_logic_ck_31 p17_logic_ck_11 0.001
R164_20 p17_logic_ck_30 p17_logic_ck_11 0.001
R164_21 p17_logic_ck_29 p17_logic_ck_11 0.001
R164_22 p17_logic_ck_102 p17_logic_ck_83 0.001
R164_23 p17_logic_ck_103 p17_logic_ck_83 0.001
R164_24 p17_logic_ck_101 p17_logic_ck_83 0.001
R164_25 p17_logic_ck_76 p17_logic_ck_59 0.001
R164_26 p17_logic_ck_52 p17_logic_ck_35 0.001
R164_27 p17_logic_ck_28 p17_logic_ck_11 0.001
R164_28 p17_logic_ck_100 p17_logic_ck_83 0.001
R164_29 p17_logic_ck_75 p17_logic_ck_60 0.001
R164_30 p17_logic_ck_51 p17_logic_ck_36 0.001
R164_31 p17_logic_ck_27 p17_logic_ck_12 0.001
R164_32 p17_logic_ck_99 p17_logic_ck_84 0.001
R164_33 p17_logic_ck_73 p17_logic_ck_60 0.001
R164_34 p17_logic_ck_72 p17_logic_ck_60 0.001
R164_35 p17_logic_ck_71 p17_logic_ck_60 0.001
R164_36 p17_logic_ck_74 p17_logic_ck_60 0.001
R164_37 p17_logic_ck_48 p17_logic_ck_36 0.001
R164_38 p17_logic_ck_49 p17_logic_ck_36 0.001
R164_39 p17_logic_ck_47 p17_logic_ck_36 0.001
R164_40 p17_logic_ck_50 p17_logic_ck_36 0.001
R164_41 p17_logic_ck_25 p17_logic_ck_12 0.001
R164_42 p17_logic_ck_24 p17_logic_ck_12 0.001
R164_43 p17_logic_ck_23 p17_logic_ck_12 0.001
R164_44 p17_logic_ck_26 p17_logic_ck_12 0.001
R164_45 p17_logic_ck_95 p17_logic_ck_84 0.001
R164_46 p17_logic_ck_96 p17_logic_ck_84 0.001
R164_47 p17_logic_ck_97 p17_logic_ck_84 0.001
R164_48 p17_logic_ck_98 p17_logic_ck_84 0.001
R164_49 p17_logic_ck_70 p17_logic_ck_60 0.001
R164_50 p17_logic_ck_69 p17_logic_ck_60 0.001
R164_51 p17_logic_ck_68 p17_logic_ck_60 0.001
R164_52 p17_logic_ck_67 p17_logic_ck_60 0.001
R164_53 p17_logic_ck_45 p17_logic_ck_36 0.001
R164_54 p17_logic_ck_46 p17_logic_ck_36 0.001
R164_55 p17_logic_ck_43 p17_logic_ck_36 0.001
R164_56 p17_logic_ck_44 p17_logic_ck_36 0.001
R164_57 p17_logic_ck_22 p17_logic_ck_12 0.001
R164_58 p17_logic_ck_21 p17_logic_ck_12 0.001
R164_59 p17_logic_ck_20 p17_logic_ck_12 0.001
R164_60 p17_logic_ck_19 p17_logic_ck_12 0.001
R164_61 p17_logic_ck_93 p17_logic_ck_84 0.001
R164_62 p17_logic_ck_94 p17_logic_ck_84 0.001
R164_63 p17_logic_ck_91 p17_logic_ck_84 0.001
R164_64 p17_logic_ck_92 p17_logic_ck_84 0.001
R164_65 p17_logic_ck_64 p17_logic_ck_60 0.001
R164_66 p17_logic_ck_63 p17_logic_ck_60 0.001
R164_67 p17_logic_ck_62 p17_logic_ck_60 0.001
R164_68 p17_logic_ck_65 p17_logic_ck_60 0.001
R164_69 p17_logic_ck_66 p17_logic_ck_60 0.001
R164_70 p17_logic_ck_39 p17_logic_ck_36 0.001
R164_71 p17_logic_ck_40 p17_logic_ck_36 0.001
R164_72 p17_logic_ck_41 p17_logic_ck_36 0.001
R164_73 p17_logic_ck_38 p17_logic_ck_36 0.001
R164_74 p17_logic_ck_42 p17_logic_ck_36 0.001
R164_75 p17_logic_ck_14 p17_logic_ck_12 0.001
R164_76 p17_logic_ck_17 p17_logic_ck_12 0.001
R164_77 p17_logic_ck_16 p17_logic_ck_12 0.001
R164_78 p17_logic_ck_15 p17_logic_ck_12 0.001
R164_79 p17_logic_ck_18 p17_logic_ck_12 0.001
R164_80 p17_logic_ck_86 p17_logic_ck_84 0.001
R164_81 p17_logic_ck_87 p17_logic_ck_84 0.001
R164_82 p17_logic_ck_88 p17_logic_ck_84 0.001
R164_83 p17_logic_ck_89 p17_logic_ck_84 0.001
R164_84 p17_logic_ck_90 p17_logic_ck_84 0.001
R164_85 p17_logic_ck_109 p17_logic_ck_108 0.054
R164_86 p17_logic_ck_107 p17_logic_ck_111 0.756
R164_87 p17_logic_ck_108 p17_logic_ck_107 0.001
R164_88 p17_logic_ck_112 p17_logic_ck_109 0.054
R164_89 p17_logic_ck_110 p17_logic_ck_115 0.756
R164_90 p17_logic_ck_111 p17_logic_ck_110 0.001
R164_91 p17_logic_ck_113 p17_logic_ck_112 0.001
R164_92 p17_logic_ck_116 p17_logic_ck_113 0.756
R164_93 p17_logic_ck_114 p17_logic_ck_119 0.756
R164_94 p17_logic_ck_115 p17_logic_ck_114 0.001
R164_95 p17_logic_ck_117 p17_logic_ck_116 0.001
R164_96 p17_logic_ck_120 p17_logic_ck_117 0.756
R164_97 p17_logic_ck_118 p17_logic_ck_123 0.756
R164_98 p17_logic_ck_119 p17_logic_ck_118 0.001
R164_99 p17_logic_ck_121 p17_logic_ck_120 0.001
R164_100 p17_logic_ck_124 p17_logic_ck_121 0.756
R164_101 p17_logic_ck_122 p17_logic_ck_127 0.756
R164_102 p17_logic_ck_123 p17_logic_ck_122 0.001
R164_103 p17_logic_ck_125 p17_logic_ck_124 0.001
R164_104 p17_logic_ck_128 p17_logic_ck_125 0.756
R164_105 p17_logic_ck_86 p17_logic_ck_85 0.001
R164_106 p17_logic_ck_87 p17_logic_ck_86 0.108
R164_107 p17_logic_ck_88 p17_logic_ck_87 0.108
R164_108 p17_logic_ck_89 p17_logic_ck_88 0.108
R164_109 p17_logic_ck_90 p17_logic_ck_89 0.108
R164_110 p17_logic_ck_91 p17_logic_ck_90 0.108
R164_111 p17_logic_ck_92 p17_logic_ck_91 0.108
R164_112 p17_logic_ck_93 p17_logic_ck_92 0.108
R164_113 p17_logic_ck_94 p17_logic_ck_93 0.108
R164_114 p17_logic_ck_95 p17_logic_ck_94 0.108
R164_115 p17_logic_ck_96 p17_logic_ck_95 0.108
R164_116 p17_logic_ck_97 p17_logic_ck_96 0.108
R164_117 p17_logic_ck_98 p17_logic_ck_97 0.108
R164_118 p17_logic_ck_99 p17_logic_ck_98 0.108
R164_119 p17_logic_ck_100 p17_logic_ck_99 0.864
R164_120 p17_logic_ck_101 p17_logic_ck_100 0.108
R164_121 p17_logic_ck_102 p17_logic_ck_101 0.108
R164_122 p17_logic_ck_103 p17_logic_ck_102 0.108
R164_123 p17_logic_ck_104 p17_logic_ck_103 0.108
R164_124 p17_logic_ck_105 p17_logic_ck_104 0.108
R164_125 p17_logic_ck_106 p17_logic_ck_105 0.001
R164_126 p17_logic_ck_14 p17_logic_ck_13 0.001
R164_127 p17_logic_ck_15 p17_logic_ck_14 0.108
R164_128 p17_logic_ck_16 p17_logic_ck_15 0.108
R164_129 p17_logic_ck_17 p17_logic_ck_16 0.108
R164_130 p17_logic_ck_18 p17_logic_ck_17 0.108
R164_131 p17_logic_ck_19 p17_logic_ck_18 0.108
R164_132 p17_logic_ck_20 p17_logic_ck_19 0.108
R164_133 p17_logic_ck_21 p17_logic_ck_20 0.108
R164_134 p17_logic_ck_22 p17_logic_ck_21 0.108
R164_135 p17_logic_ck_23 p17_logic_ck_22 0.108
R164_136 p17_logic_ck_24 p17_logic_ck_23 0.108
R164_137 p17_logic_ck_25 p17_logic_ck_24 0.108
R164_138 p17_logic_ck_26 p17_logic_ck_25 0.108
R164_139 p17_logic_ck_27 p17_logic_ck_26 0.108
R164_140 p17_logic_ck_28 p17_logic_ck_27 0.864
R164_141 p17_logic_ck_29 p17_logic_ck_28 0.108
R164_142 p17_logic_ck_30 p17_logic_ck_29 0.108
R164_143 p17_logic_ck_31 p17_logic_ck_30 0.108
R164_144 p17_logic_ck_32 p17_logic_ck_31 0.108
R164_145 p17_logic_ck_33 p17_logic_ck_32 0.108
R164_146 p17_logic_ck_34 p17_logic_ck_33 0.001
R164_147 p17_logic_ck_38 p17_logic_ck_37 0.001
R164_148 p17_logic_ck_39 p17_logic_ck_38 0.108
R164_149 p17_logic_ck_40 p17_logic_ck_39 0.108
R164_150 p17_logic_ck_41 p17_logic_ck_40 0.108
R164_151 p17_logic_ck_42 p17_logic_ck_41 0.108
R164_152 p17_logic_ck_43 p17_logic_ck_42 0.108
R164_153 p17_logic_ck_44 p17_logic_ck_43 0.108
R164_154 p17_logic_ck_45 p17_logic_ck_44 0.108
R164_155 p17_logic_ck_46 p17_logic_ck_45 0.108
R164_156 p17_logic_ck_47 p17_logic_ck_46 0.108
R164_157 p17_logic_ck_48 p17_logic_ck_47 0.108
R164_158 p17_logic_ck_49 p17_logic_ck_48 0.108
R164_159 p17_logic_ck_50 p17_logic_ck_49 0.108
R164_160 p17_logic_ck_51 p17_logic_ck_50 0.108
R164_161 p17_logic_ck_52 p17_logic_ck_51 0.864
R164_162 p17_logic_ck_53 p17_logic_ck_52 0.108
R164_163 p17_logic_ck_54 p17_logic_ck_53 0.108
R164_164 p17_logic_ck_55 p17_logic_ck_54 0.108
R164_165 p17_logic_ck_56 p17_logic_ck_55 0.108
R164_166 p17_logic_ck_57 p17_logic_ck_56 0.108
R164_167 p17_logic_ck_58 p17_logic_ck_57 0.001
R164_168 p17_logic_ck_62 p17_logic_ck_61 0.001
R164_169 p17_logic_ck_63 p17_logic_ck_62 0.108
R164_170 p17_logic_ck_64 p17_logic_ck_63 0.108
R164_171 p17_logic_ck_65 p17_logic_ck_64 0.108
R164_172 p17_logic_ck_66 p17_logic_ck_65 0.108
R164_173 p17_logic_ck_67 p17_logic_ck_66 0.108
R164_174 p17_logic_ck_68 p17_logic_ck_67 0.108
R164_175 p17_logic_ck_69 p17_logic_ck_68 0.108
R164_176 p17_logic_ck_70 p17_logic_ck_69 0.108
R164_177 p17_logic_ck_71 p17_logic_ck_70 0.108
R164_178 p17_logic_ck_72 p17_logic_ck_71 0.108
R164_179 p17_logic_ck_73 p17_logic_ck_72 0.108
R164_180 p17_logic_ck_74 p17_logic_ck_73 0.108
R164_181 p17_logic_ck_75 p17_logic_ck_74 0.108
R164_182 p17_logic_ck_76 p17_logic_ck_75 0.864
R164_183 p17_logic_ck_77 p17_logic_ck_76 0.108
R164_184 p17_logic_ck_78 p17_logic_ck_77 0.108
R164_185 p17_logic_ck_79 p17_logic_ck_78 0.108
R164_186 p17_logic_ck_80 p17_logic_ck_79 0.108
R164_187 p17_logic_ck_81 p17_logic_ck_80 0.108
R164_188 p17_logic_ck_82 p17_logic_ck_81 0.001
R164_189 p17_logic_ck_126 p17_logic_ck_130 0.108
R164_190 p17_logic_ck_127 p17_logic_ck_126 0.001
R164_191 p17_logic_ck_129 p17_logic_ck_128 0.001
R164_192 p17_logic_ck_131 p17_logic_ck_129 0.756
R164_193 p17_logic_ck_133 p17_logic_ck_130 0.432
R164_194 p17_logic_ck_132 p17_logic_ck_131 0.001
R164_195 p17_logic_ck_139 p17_logic_ck_132 0.054
R164_196 p17_logic_ck_134 p17_logic_ck_133 0.001
R164_197 p17_logic_ck_135 p17_logic_ck_134 0.432
R164_198 p17_logic_ck_136 p17_logic_ck_135 0.054
R164_199 p17_logic_ck_137 p17_logic_ck_136 0.054
R164_200 p17_logic_ck_138 p17_logic_ck_137 0.054
R164_201 p17_logic_ck_140 p17_logic_ck_138 0.108
R164_202 p17_logic_ck_139 p17_logic_ck_143 0.108
R164_203 p17_logic_ck_141 p17_logic_ck_140 0.001
R164_204 p17_logic_ck_144 p17_logic_ck_141 0.756
R164_205 p17_logic_ck_142 p17_logic_ck_147 0.756
R164_206 p17_logic_ck_143 p17_logic_ck_142 0.001
R164_207 p17_logic_ck_145 p17_logic_ck_144 0.001
R164_208 p17_logic_ck_148 p17_logic_ck_145 0.756
R164_209 p17_logic_ck_146 p17_logic_ck_151 0.756
R164_210 p17_logic_ck_147 p17_logic_ck_146 0.001
R164_211 p17_logic_ck_149 p17_logic_ck_148 0.001
R164_212 p17_logic_ck_152 p17_logic_ck_149 0.756
R164_213 p17_logic_ck_150 p17_logic_ck_155 0.756
R164_214 p17_logic_ck_151 p17_logic_ck_150 0.001
R164_215 p17_logic_ck_153 p17_logic_ck_152 0.001
R164_216 p17_logic_ck_156 p17_logic_ck_153 0.432
R164_217 p17_logic_ck_154 p17_logic_ck_161 0.756
R164_218 p17_logic_ck_155 p17_logic_ck_154 0.001
R164_219 p17_logic_ck_157 p17_logic_ck_156 0.054
R164_220 p17_logic_ck_158 p17_logic_ck_157 0.001
R164_221 p17_logic_ck_159 p17_logic_ck_158 0.594
R164_222 p17_logic_ck_160 p17_logic_ck_159 0.162
R164_223 p17_logic_ck_161 p17_logic_ck_160 0.001
R164_224 p17_logic_ck_5 p17_logic_ck_4 0.001
R164_225 p17_logic_ck_6 p17_logic_ck_5 0.108
R164_226 p17_logic_ck_7 p17_logic_ck_6 0.108
R164_227 p17_logic_ck_10 p17_logic_ck_7 1.836
R164_228 p17_logic_ck_8 p17_logic_ck_10 0.001
R164_229 p17_logic_ck_10 p17_logic_ck_9 0.54
R164_230 p17_logic_ck_2 p17_logic_ck 144
R164_231 p17_logic_ck_3 p17_logic_ck_2 208.8

C9688 p17_logic_ck_109 vss 1.2636e-16
C9689 p17_logic_ck_108 vss 1.2636e-16
C9690 p17_logic_ck_107 vss 1.66212e-15
C9691 p17_logic_ck_111 vss 1.66212e-15
C9692 p17_logic_ck_108 vss 9.72e-18
C9693 p17_logic_ck_107 vss 9.72e-18
C9694 p17_logic_ck_112 vss 1.1664e-16
C9695 p17_logic_ck_109 vss 1.1664e-16
C9696 p17_logic_ck_110 vss 1.66212e-15
C9697 p17_logic_ck_115 vss 1.66212e-15
C9698 p17_logic_ck_111 vss 9.72e-18
C9699 p17_logic_ck_110 vss 9.72e-18
C9700 p17_logic_ck_113 vss 1.944e-17
C9701 p17_logic_ck_112 vss 1.944e-17
C9702 p17_logic_ck_116 vss 1.6524e-15
C9703 p17_logic_ck_113 vss 1.6524e-15
C9704 p17_logic_ck_114 vss 1.66212e-15
C9705 p17_logic_ck_119 vss 1.66212e-15
C9706 p17_logic_ck_115 vss 9.72e-18
C9707 p17_logic_ck_114 vss 9.72e-18
C9708 p17_logic_ck_117 vss 9.72e-18
C9709 p17_logic_ck_116 vss 9.72e-18
C9710 p17_logic_ck_120 vss 1.66212e-15
C9711 p17_logic_ck_117 vss 1.66212e-15
C9712 p17_logic_ck_118 vss 1.66212e-15
C9713 p17_logic_ck_123 vss 1.66212e-15
C9714 p17_logic_ck_119 vss 9.72e-18
C9715 p17_logic_ck_118 vss 9.72e-18
C9716 p17_logic_ck_121 vss 9.72e-18
C9717 p17_logic_ck_120 vss 9.72e-18
C9718 p17_logic_ck_124 vss 1.66212e-15
C9719 p17_logic_ck_121 vss 1.66212e-15
C9720 p17_logic_ck_122 vss 1.6524e-15
C9721 p17_logic_ck_127 vss 1.6524e-15
C9722 p17_logic_ck_123 vss 9.72e-18
C9723 p17_logic_ck_122 vss 9.72e-18
C9724 p17_logic_ck_125 vss 9.72e-18
C9725 p17_logic_ck_124 vss 9.72e-18
C9726 p17_logic_ck_128 vss 1.66212e-15
C9727 p17_logic_ck_125 vss 1.66212e-15
C9728 p17_logic_ck_86 vss 1.40901e-17
C9729 p17_logic_ck_85 vss 1.40901e-17
C9730 p17_logic_ck_87 vss 3.13114e-17
C9731 p17_logic_ck_86 vss 3.13114e-17
C9732 p17_logic_ck_88 vss 3.13114e-17
C9733 p17_logic_ck_87 vss 3.13114e-17
C9734 p17_logic_ck_89 vss 3.13114e-17
C9735 p17_logic_ck_88 vss 3.13114e-17
C9736 p17_logic_ck_90 vss 3.13114e-17
C9737 p17_logic_ck_89 vss 3.13114e-17
C9738 p17_logic_ck_91 vss 3.13114e-17
C9739 p17_logic_ck_90 vss 3.13114e-17
C9740 p17_logic_ck_92 vss 3.13114e-17
C9741 p17_logic_ck_91 vss 3.13114e-17
C9742 p17_logic_ck_93 vss 3.13114e-17
C9743 p17_logic_ck_92 vss 3.13114e-17
C9744 p17_logic_ck_94 vss 3.13114e-17
C9745 p17_logic_ck_93 vss 3.13114e-17
C9746 p17_logic_ck_95 vss 3.13114e-17
C9747 p17_logic_ck_94 vss 3.13114e-17
C9748 p17_logic_ck_96 vss 3.13114e-17
C9749 p17_logic_ck_95 vss 3.13114e-17
C9750 p17_logic_ck_97 vss 3.13114e-17
C9751 p17_logic_ck_96 vss 3.13114e-17
C9752 p17_logic_ck_98 vss 3.13114e-17
C9753 p17_logic_ck_97 vss 3.13114e-17
C9754 p17_logic_ck_99 vss 3.13114e-17
C9755 p17_logic_ck_98 vss 3.13114e-17
C9756 p17_logic_ck_100 vss 2.42663e-16
C9757 p17_logic_ck_99 vss 2.42663e-16
C9758 p17_logic_ck_101 vss 3.91392e-17
C9759 p17_logic_ck_100 vss 3.91392e-17
C9760 p17_logic_ck_102 vss 3.91392e-17
C9761 p17_logic_ck_101 vss 3.91392e-17
C9762 p17_logic_ck_103 vss 3.91392e-17
C9763 p17_logic_ck_102 vss 3.91392e-17
C9764 p17_logic_ck_104 vss 4.6967e-17
C9765 p17_logic_ck_103 vss 4.6967e-17
C9766 p17_logic_ck_105 vss 5.47949e-17
C9767 p17_logic_ck_104 vss 5.47949e-17
C9768 p17_logic_ck_106 vss 1.40901e-17
C9769 p17_logic_ck_105 vss 1.40901e-17
C9770 p17_logic_ck_14 vss 1.40901e-17
C9771 p17_logic_ck_13 vss 1.40901e-17
C9772 p17_logic_ck_15 vss 3.13114e-17
C9773 p17_logic_ck_14 vss 3.13114e-17
C9774 p17_logic_ck_16 vss 3.13114e-17
C9775 p17_logic_ck_15 vss 3.13114e-17
C9776 p17_logic_ck_17 vss 3.13114e-17
C9777 p17_logic_ck_16 vss 3.13114e-17
C9778 p17_logic_ck_18 vss 3.13114e-17
C9779 p17_logic_ck_17 vss 3.13114e-17
C9780 p17_logic_ck_19 vss 3.13114e-17
C9781 p17_logic_ck_18 vss 3.13114e-17
C9782 p17_logic_ck_20 vss 3.13114e-17
C9783 p17_logic_ck_19 vss 3.13114e-17
C9784 p17_logic_ck_21 vss 3.13114e-17
C9785 p17_logic_ck_20 vss 3.13114e-17
C9786 p17_logic_ck_22 vss 3.13114e-17
C9787 p17_logic_ck_21 vss 3.13114e-17
C9788 p17_logic_ck_23 vss 3.13114e-17
C9789 p17_logic_ck_22 vss 3.13114e-17
C9790 p17_logic_ck_24 vss 3.13114e-17
C9791 p17_logic_ck_23 vss 3.13114e-17
C9792 p17_logic_ck_25 vss 3.13114e-17
C9793 p17_logic_ck_24 vss 3.13114e-17
C9794 p17_logic_ck_26 vss 3.13114e-17
C9795 p17_logic_ck_25 vss 3.13114e-17
C9796 p17_logic_ck_27 vss 3.13114e-17
C9797 p17_logic_ck_26 vss 3.13114e-17
C9798 p17_logic_ck_28 vss 2.42663e-16
C9799 p17_logic_ck_27 vss 2.42663e-16
C9800 p17_logic_ck_29 vss 3.91392e-17
C9801 p17_logic_ck_28 vss 3.91392e-17
C9802 p17_logic_ck_30 vss 3.91392e-17
C9803 p17_logic_ck_29 vss 3.91392e-17
C9804 p17_logic_ck_31 vss 3.91392e-17
C9805 p17_logic_ck_30 vss 3.91392e-17
C9806 p17_logic_ck_32 vss 4.6967e-17
C9807 p17_logic_ck_31 vss 4.6967e-17
C9808 p17_logic_ck_33 vss 5.47949e-17
C9809 p17_logic_ck_32 vss 5.47949e-17
C9810 p17_logic_ck_34 vss 1.40901e-17
C9811 p17_logic_ck_33 vss 1.40901e-17
C9812 p17_logic_ck_38 vss 1.40901e-17
C9813 p17_logic_ck_37 vss 1.40901e-17
C9814 p17_logic_ck_39 vss 3.13114e-17
C9815 p17_logic_ck_38 vss 3.13114e-17
C9816 p17_logic_ck_40 vss 3.13114e-17
C9817 p17_logic_ck_39 vss 3.13114e-17
C9818 p17_logic_ck_41 vss 3.13114e-17
C9819 p17_logic_ck_40 vss 3.13114e-17
C9820 p17_logic_ck_42 vss 3.13114e-17
C9821 p17_logic_ck_41 vss 3.13114e-17
C9822 p17_logic_ck_43 vss 3.13114e-17
C9823 p17_logic_ck_42 vss 3.13114e-17
C9824 p17_logic_ck_44 vss 3.13114e-17
C9825 p17_logic_ck_43 vss 3.13114e-17
C9826 p17_logic_ck_45 vss 3.13114e-17
C9827 p17_logic_ck_44 vss 3.13114e-17
C9828 p17_logic_ck_46 vss 3.13114e-17
C9829 p17_logic_ck_45 vss 3.13114e-17
C9830 p17_logic_ck_47 vss 3.13114e-17
C9831 p17_logic_ck_46 vss 3.13114e-17
C9832 p17_logic_ck_48 vss 3.13114e-17
C9833 p17_logic_ck_47 vss 3.13114e-17
C9834 p17_logic_ck_49 vss 3.13114e-17
C9835 p17_logic_ck_48 vss 3.13114e-17
C9836 p17_logic_ck_50 vss 3.13114e-17
C9837 p17_logic_ck_49 vss 3.13114e-17
C9838 p17_logic_ck_51 vss 3.13114e-17
C9839 p17_logic_ck_50 vss 3.13114e-17
C9840 p17_logic_ck_52 vss 2.42663e-16
C9841 p17_logic_ck_51 vss 2.42663e-16
C9842 p17_logic_ck_53 vss 3.91392e-17
C9843 p17_logic_ck_52 vss 3.91392e-17
C9844 p17_logic_ck_54 vss 3.91392e-17
C9845 p17_logic_ck_53 vss 3.91392e-17
C9846 p17_logic_ck_55 vss 3.91392e-17
C9847 p17_logic_ck_54 vss 3.91392e-17
C9848 p17_logic_ck_56 vss 4.6967e-17
C9849 p17_logic_ck_55 vss 4.6967e-17
C9850 p17_logic_ck_57 vss 5.47949e-17
C9851 p17_logic_ck_56 vss 5.47949e-17
C9852 p17_logic_ck_58 vss 1.40901e-17
C9853 p17_logic_ck_57 vss 1.40901e-17
C9854 p17_logic_ck_62 vss 1.40901e-17
C9855 p17_logic_ck_61 vss 1.40901e-17
C9856 p17_logic_ck_63 vss 3.13114e-17
C9857 p17_logic_ck_62 vss 3.13114e-17
C9858 p17_logic_ck_64 vss 3.13114e-17
C9859 p17_logic_ck_63 vss 3.13114e-17
C9860 p17_logic_ck_65 vss 3.13114e-17
C9861 p17_logic_ck_64 vss 3.13114e-17
C9862 p17_logic_ck_66 vss 3.13114e-17
C9863 p17_logic_ck_65 vss 3.13114e-17
C9864 p17_logic_ck_67 vss 3.13114e-17
C9865 p17_logic_ck_66 vss 3.13114e-17
C9866 p17_logic_ck_68 vss 3.13114e-17
C9867 p17_logic_ck_67 vss 3.13114e-17
C9868 p17_logic_ck_69 vss 3.13114e-17
C9869 p17_logic_ck_68 vss 3.13114e-17
C9870 p17_logic_ck_70 vss 3.13114e-17
C9871 p17_logic_ck_69 vss 3.13114e-17
C9872 p17_logic_ck_71 vss 3.13114e-17
C9873 p17_logic_ck_70 vss 3.13114e-17
C9874 p17_logic_ck_72 vss 3.13114e-17
C9875 p17_logic_ck_71 vss 3.13114e-17
C9876 p17_logic_ck_73 vss 3.13114e-17
C9877 p17_logic_ck_72 vss 3.13114e-17
C9878 p17_logic_ck_74 vss 3.13114e-17
C9879 p17_logic_ck_73 vss 3.13114e-17
C9880 p17_logic_ck_75 vss 3.13114e-17
C9881 p17_logic_ck_74 vss 3.13114e-17
C9882 p17_logic_ck_76 vss 2.42663e-16
C9883 p17_logic_ck_75 vss 2.42663e-16
C9884 p17_logic_ck_77 vss 3.91392e-17
C9885 p17_logic_ck_76 vss 3.91392e-17
C9886 p17_logic_ck_78 vss 3.91392e-17
C9887 p17_logic_ck_77 vss 3.91392e-17
C9888 p17_logic_ck_79 vss 3.91392e-17
C9889 p17_logic_ck_78 vss 3.91392e-17
C9890 p17_logic_ck_80 vss 4.6967e-17
C9891 p17_logic_ck_79 vss 4.6967e-17
C9892 p17_logic_ck_81 vss 5.47949e-17
C9893 p17_logic_ck_80 vss 5.47949e-17
C9894 p17_logic_ck_82 vss 1.40901e-17
C9895 p17_logic_ck_81 vss 1.40901e-17
C9896 p17_logic_ck_126 vss 2.8188e-16
C9897 p17_logic_ck_130 vss 2.8188e-16
C9898 p17_logic_ck_127 vss 1.944e-17
C9899 p17_logic_ck_126 vss 1.944e-17
C9900 p17_logic_ck_129 vss 9.72e-18
C9901 p17_logic_ck_128 vss 9.72e-18
C9902 p17_logic_ck_131 vss 1.66212e-15
C9903 p17_logic_ck_129 vss 1.66212e-15
C9904 p17_logic_ck_133 vss 9.5256e-16
C9905 p17_logic_ck_130 vss 9.5256e-16
C9906 p17_logic_ck_132 vss 9.72e-18
C9907 p17_logic_ck_131 vss 9.72e-18
C9908 p17_logic_ck_139 vss 1.2636e-16
C9909 p17_logic_ck_132 vss 1.2636e-16
C9910 p17_logic_ck_134 vss 1.944e-17
C9911 p17_logic_ck_133 vss 1.944e-17
C9912 p17_logic_ck_135 vss 1.04004e-15
C9913 p17_logic_ck_134 vss 1.04004e-15
C9914 p17_logic_ck_136 vss 1.1664e-16
C9915 p17_logic_ck_135 vss 1.1664e-16
C9916 p17_logic_ck_137 vss 1.1664e-16
C9917 p17_logic_ck_136 vss 1.1664e-16
C9918 p17_logic_ck_138 vss 1.1664e-16
C9919 p17_logic_ck_137 vss 1.1664e-16
C9920 p17_logic_ck_140 vss 2.6244e-16
C9921 p17_logic_ck_138 vss 2.6244e-16
C9922 p17_logic_ck_139 vss 2.7216e-16
C9923 p17_logic_ck_143 vss 2.7216e-16
C9924 p17_logic_ck_141 vss 1.944e-17
C9925 p17_logic_ck_140 vss 1.944e-17
C9926 p17_logic_ck_144 vss 1.6524e-15
C9927 p17_logic_ck_141 vss 1.6524e-15
C9928 p17_logic_ck_142 vss 1.6524e-15
C9929 p17_logic_ck_147 vss 1.6524e-15
C9930 p17_logic_ck_143 vss 1.944e-17
C9931 p17_logic_ck_142 vss 1.944e-17
C9932 p17_logic_ck_145 vss 9.72e-18
C9933 p17_logic_ck_144 vss 9.72e-18
C9934 p17_logic_ck_148 vss 1.66212e-15
C9935 p17_logic_ck_145 vss 1.66212e-15
C9936 p17_logic_ck_146 vss 1.6524e-15
C9937 p17_logic_ck_151 vss 1.6524e-15
C9938 p17_logic_ck_147 vss 1.944e-17
C9939 p17_logic_ck_146 vss 1.944e-17
C9940 p17_logic_ck_149 vss 9.72e-18
C9941 p17_logic_ck_148 vss 9.72e-18
C9942 p17_logic_ck_152 vss 1.66212e-15
C9943 p17_logic_ck_149 vss 1.66212e-15
C9944 p17_logic_ck_150 vss 1.6524e-15
C9945 p17_logic_ck_155 vss 1.6524e-15
C9946 p17_logic_ck_151 vss 1.944e-17
C9947 p17_logic_ck_150 vss 1.944e-17
C9948 p17_logic_ck_153 vss 9.72e-18
C9949 p17_logic_ck_152 vss 9.72e-18
C9950 p17_logic_ck_156 vss 9.6228e-16
C9951 p17_logic_ck_153 vss 9.6228e-16
C9952 p17_logic_ck_154 vss 1.6524e-15
C9953 p17_logic_ck_161 vss 1.6524e-15
C9954 p17_logic_ck_155 vss 1.944e-17
C9955 p17_logic_ck_154 vss 1.944e-17
C9956 p17_logic_ck_157 vss 1.2636e-16
C9957 p17_logic_ck_156 vss 1.2636e-16
C9958 p17_logic_ck_158 vss 1.944e-17
C9959 p17_logic_ck_157 vss 1.944e-17
C9960 p17_logic_ck_159 vss 1.29276e-15
C9961 p17_logic_ck_158 vss 1.29276e-15
C9962 p17_logic_ck_160 vss 3.5964e-16
C9963 p17_logic_ck_159 vss 3.5964e-16
C9964 p17_logic_ck_161 vss 1.944e-17
C9965 p17_logic_ck_160 vss 1.944e-17
C9966 p17_logic_ck_5 vss 1.3157e-17
C9967 p17_logic_ck_4 vss 1.3157e-17
C9968 p17_logic_ck_6 vss 2.92378e-17
C9969 p17_logic_ck_5 vss 2.92378e-17
C9970 p17_logic_ck_7 vss 2.92378e-17
C9971 p17_logic_ck_6 vss 2.92378e-17
C9972 p17_logic_ck_10 vss 3.36234e-16
C9973 p17_logic_ck_7 vss 3.36234e-16
C9974 p17_logic_ck_8 vss 1.3157e-17
C9975 p17_logic_ck_10 vss 1.3157e-17
C9976 p17_logic_ck_10 vss 1.02332e-16
C9977 p17_logic_ck_9 vss 1.02332e-16
C9978 p17_logic_ck_2 vss 1.60405e-16
C9979 p17_logic_ck vss 1.60405e-16
C9980 p17_logic_ck_3 vss 2.30825e-16
C9981 p17_logic_ck_2 vss 2.30825e-16

R165_1 n6442_1 n6442_32 0.001
R165_2 n6442_1 n6442_33 0.001
R165_3 n6442_1 n6442_34 0.001
R165_4 n6442_1 n6442_31 0.001
R165_5 n6442_1 n6442_28 0.001
R165_6 n6442_1 n6442_29 0.001
R165_7 n6442_1 n6442_30 0.001
R165_8 n6442_1 n6442_25 0.001
R165_9 n6442_1 n6442_26 0.001
R165_10 n6442_1 n6442_27 0.001
R165_11 n6442_14 n6442_11 0.001
R165_12 n6442_18 n6442_13 0.001
R165_13 n6442_19 n6442_13 0.001
R165_14 n6442_15 n6442_13 0.001
R165_15 n6442_16 n6442_13 0.001
R165_16 n6442_17 n6442_13 0.001
R165_17 n6442_3 n6442_2 43.2
R165_18 n6442_12 n6442_3 43.2
R165_19 n6442_4 n6442_12 43.2
R165_20 n6442_5 n6442_4 43.2
R165_21 n6442_7 n6442_6 43.2
R165_22 n6442 n6442_7 43.2
R165_23 n6442_8 n6442 43.2
R165_24 n6442_9 n6442_8 43.2
R165_25 n6442_11 n6442 28.8
R165_26 n6442_12 n6442_11 36
R165_27 n6442_22 n6442_14 0.756
R165_28 n6442_16 n6442_15 0.108
R165_29 n6442_17 n6442_16 0.108
R165_30 n6442_18 n6442_17 0.108
R165_31 n6442_19 n6442_18 0.108
R165_32 n6442_20 n6442_19 0.108
R165_33 n6442_21 n6442_20 0.001
R165_34 n6442_22 n6442_21 0.108
R165_35 n6442_23 n6442_22 0.108
R165_36 n6442_24 n6442_23 0.001
R165_37 n6442_25 n6442_24 0.216
R165_38 n6442_26 n6442_25 0.108
R165_39 n6442_27 n6442_26 0.108
R165_40 n6442_28 n6442_27 0.108
R165_41 n6442_29 n6442_28 0.108
R165_42 n6442_30 n6442_29 0.108
R165_43 n6442_31 n6442_30 0.108
R165_44 n6442_32 n6442_31 0.108
R165_45 n6442_33 n6442_32 0.108
R165_46 n6442_34 n6442_33 0.108

C9982 n6442_3 vss 4.69476e-17
C9983 n6442_2 vss 4.69476e-17
C9984 n6442_12 vss 4.69476e-17
C9985 n6442_3 vss 4.69476e-17
C9986 n6442_4 vss 4.69476e-17
C9987 n6442_12 vss 4.69476e-17
C9988 n6442_5 vss 4.69476e-17
C9989 n6442_4 vss 4.69476e-17
C9990 n6442_7 vss 4.69476e-17
C9991 n6442_6 vss 4.69476e-17
C9992 n6442 vss 4.69476e-17
C9993 n6442_7 vss 4.69476e-17
C9994 n6442_8 vss 4.69476e-17
C9995 n6442 vss 4.69476e-17
C9996 n6442_9 vss 4.69476e-17
C9997 n6442_8 vss 4.69476e-17
C9998 n6442_11 vss 2.67361e-16
C9999 n6442 vss 2.67361e-16
C10000 n6442_12 vss 3.46579e-16
C10001 n6442_11 vss 3.46579e-16
C10002 n6442_22 vss 1.38879e-16
C10003 n6442_14 vss 1.38879e-16
C10004 n6442_16 vss 2.92378e-17
C10005 n6442_15 vss 2.92378e-17
C10006 n6442_17 vss 2.92378e-17
C10007 n6442_16 vss 2.92378e-17
C10008 n6442_18 vss 2.92378e-17
C10009 n6442_17 vss 2.92378e-17
C10010 n6442_19 vss 2.92378e-17
C10011 n6442_18 vss 2.92378e-17
C10012 n6442_20 vss 3.06996e-17
C10013 n6442_19 vss 3.06996e-17
C10014 n6442_21 vss 3.00465e-17
C10015 n6442_20 vss 3.00465e-17
C10016 n6442_22 vss 3.06996e-17
C10017 n6442_21 vss 3.06996e-17
C10018 n6442_23 vss 3.06996e-17
C10019 n6442_22 vss 3.06996e-17
C10020 n6442_24 vss 2.17002e-17
C10021 n6442_23 vss 2.17002e-17
C10022 n6442_25 vss 3.80091e-17
C10023 n6442_24 vss 3.80091e-17
C10024 n6442_26 vss 2.92378e-17
C10025 n6442_25 vss 2.92378e-17
C10026 n6442_27 vss 2.92378e-17
C10027 n6442_26 vss 2.92378e-17
C10028 n6442_28 vss 2.92378e-17
C10029 n6442_27 vss 2.92378e-17
C10030 n6442_29 vss 2.92378e-17
C10031 n6442_28 vss 2.92378e-17
C10032 n6442_30 vss 2.92378e-17
C10033 n6442_29 vss 2.92378e-17
C10034 n6442_31 vss 2.92378e-17
C10035 n6442_30 vss 2.92378e-17
C10036 n6442_32 vss 2.92378e-17
C10037 n6442_31 vss 2.92378e-17
C10038 n6442_33 vss 2.92378e-17
C10039 n6442_32 vss 2.92378e-17
C10040 n6442_34 vss 2.92378e-17
C10041 n6442_33 vss 2.92378e-17


.ends addaccu

