* glitcher

.subckt DLY4X1  VDD VSS A Y
mM0 VSS A 1 VSS TN L=1.8e-07 W=2.8e-07
mM1 3 1 VSS VSS TN L=7.2e-07 W=2.8e-07
mM2 VSS 3 4 VSS TN L=7.2e-07 W=2.8e-07
mM3 Y 4 VSS VSS TN L=1.8e-07 W=6e-07
mM4 VDD A 1 VDD TP L=1.8e-07 W=4.2e-07
mM5 3 1 VDD VDD TP L=7.2e-07 W=4.2e-07
mM6 VDD 3 4 VDD TP L=7.2e-07 W=4.2e-07
mM7 Y 4 VDD VDD TP L=1.8e-07 W=9e-07
.ends

.subckt INVX1  VDD VSS A Y
mM0 Y A VSS VSS TN L=3e-07 W=12e-07
mM1 Y A VDD VDD TP L=3e-07 W=18e-07
.ends

.subckt NOR2X1  VDD VSS A B Y
mM0 Y B VSS VSS TN L=1.8e-07 W=6e-07
mM1 VSS A Y VSS TN L=1.8e-07 W=6e-07
mM2 6 B VDD VDD TP L=1.8e-07 W=1.2e-06
mM3 Y A 6 VDD TP L=1.8e-07 W=1.2e-06
.ends

.subckt glitcher I O VDD VSS
XINV0 VDD VSS I S0 INVX1 
XINV2 VDD VSS S0 S1 INVX1 
XINV3 VDD VSS S1 S2 INVX1 
XINV4 VDD VSS S2 S3 INVX1 
XINV5 VDD VSS S3 S4 INVX1 
XINV6 VDD VSS S4 S5 INVX1 
XDLY0 VDD VSS I Idly DLY4X1
XINV7 VDD VSS Idly IdlyN INVX1
XNOR0 VDD VSS IdlyN S5 S6 NOR2X1 
XINV8 VDD VSS S6 O INVX1
.ends glitcher

