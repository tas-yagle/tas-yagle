* comb

.subckt INVX1  VDD VSS A Y
mM0 Y A VSS VSS TN L=3e-07 W=12e-07
mM1 Y A VDD VDD TP L=3e-07 W=18e-07
.ends

.subckt NOR2X1  VDD VSS A B Y
mM0 Y B VSS VSS TN L=1.8e-07 W=6e-07
mM1 VSS A Y VSS TN L=1.8e-07 W=6e-07
mM2 6 B VDD VDD TP L=1.8e-07 W=1.2e-06
mM3 Y A 6 VDD TP L=1.8e-07 W=1.2e-06
.ends

.subckt OR2X1  VDD VSS A B Y
mM0 5 A VSS VSS TN L=1.8e-07 W=3e-07
mM1 VSS B 5 VSS TN L=1.8e-07 W=3e-07
mM2 Y 5 VSS VSS TN L=1.8e-07 W=6e-07
mM3 7 A 5 VDD TP L=1.8e-07 W=5.6e-07
mM4 VDD B 7 VDD TP L=1.8e-07 W=5.6e-07
mM5 Y 5 VDD VDD TP L=1.8e-07 W=9e-07
.ends

.subckt MX2X1  VDD VSS A B S0 Y
mM0 VSS S0 3 VSS TN L=1.8e-07 W=3e-07
mM1 4 B VSS VSS TN L=1.8e-07 W=4.8e-07
mM2 7 S0 4 VSS TN L=1.8e-07 W=4.8e-07
mM3 5 3 7 VSS TN L=1.8e-07 W=4.8e-07
mM4 VSS A 5 VSS TN L=1.8e-07 W=4.8e-07
mM5 Y 7 VSS VSS TN L=1.8e-07 W=6e-07
mM6 VDD S0 3 VDD TP L=1.8e-07 W=4.2e-07
mM7 4 B VDD VDD TP L=1.8e-07 W=7.2e-07
mM8 7 3 4 VDD TP L=1.8e-07 W=7.2e-07
mM9 5 S0 7 VDD TP L=1.8e-07 W=7.2e-07
mM10 VDD A 5 VDD TP L=1.8e-07 W=7.2e-07
mM11 Y 7 VDD VDD TP L=1.8e-07 W=9e-07
.ends

.subckt comb I0 I1 I2 I3 SEL O VDD VSS
XNOR0 VDD VSS I0 I1 S0 NOR2X1 
XINV0 VDD VSS S0 S1 INVX1 
XINV1 VDD VSS I2 S2 INVX1 
XMUX0 VDD VSS S2 I3 SEL S3 MX2X1
XOR0 VDD VSS S1 S3 O OR2X1 
.ends comb

