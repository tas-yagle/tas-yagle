* Spice description of r256x8_1
* Spice driver version 700
* Date ( dd/mm/yyyy hh:mm:ss ): 20/09/2002 at 16:20:42

* INTERF adr[0] adr[1] adr[2] adr[3] adr[4] adr[5] adr[6] adr[7] ck[0] ck[1] 
* INTERF f[0] f[1] f[2] f[3] f[4] f[5] f[6] f[7] vdd vss 


.subckt r256x8_1 1332 1326 1327 1328 1320 1321 1322 1318 1234 1 1350 1347 
+ 1345 1343 1341 1339 1337 1335 1348 1351 
* NET 1 = ck[1] 
* NET 5 = rl/7.w1 
* NET 18 = rbl4/1/2.e0 
* NET 19 = rck.ckp 
* NET 25 = rl/7.e1 
* NET 26 = rl/7.tr_p 
* NET 27 = rl/7.w2 
* NET 28 = rl/7.w3 
* NET 29 = rl/7.w4 
* NET 98 = rbl4/1/2.e1 
* NET 99 = rbl4/1/2.e2 
* NET 100 = rbl4/1/2.e3 
* NET 106 = rl/6.e1 
* NET 107 = rl/6.tr_p 
* NET 108 = rl/6.w1 
* NET 109 = rl/6.w2 
* NET 110 = rl/6.w3 
* NET 111 = rl/6.w4 
* NET 224 = rbl4/1/2.e7 
* NET 225 = rbl4/1/2.e6 
* NET 226 = umf.e31 
* NET 227 = rbl4/1/2.e5 
* NET 232 = rl/5.w1 
* NET 233 = rl/5.w2 
* NET 234 = rl/5.w3 
* NET 311 = rbl4/1/2.e10 
* NET 312 = rbl4/1/2.e8 
* NET 313 = rbl4/1/2.e9 
* NET 318 = rl/5.e1 
* NET 319 = rl/5.tr_p 
* NET 320 = rl/5.w4 
* NET 321 = rl/4.w1 
* NET 322 = rl/4.w2 
* NET 459 = rbl4/1/2.e11 
* NET 460 = rbl4/1/2.e14 
* NET 461 = rbl4/1/2.e13 
* NET 462 = rbl4/1/2.e12 
* NET 467 = rl/4.e1 
* NET 468 = rl/4.tr_p 
* NET 469 = rl/4.w3 
* NET 470 = rl/4.w4 
* NET 471 = rl/3.w1 
* NET 472 = rl/3.w2 
* NET 557 = umf.e0 
* NET 558 = rbl4/1/2.e15 
* NET 559 = umf.e1 
* NET 573 = rl/3.e1 
* NET 574 = rl/3.tr_p 
* NET 575 = rl/3.w3 
* NET 576 = rl/3.w4 
* NET 577 = rl/2.w1 
* NET 578 = rl/2.w2 
* NET 691 = umf.e2 
* NET 692 = umf.e5 
* NET 693 = umf.e4 
* NET 694 = umf.e3 
* NET 716 = rl/2.e1 
* NET 717 = rl/2.tr_p 
* NET 718 = rl/2.w3 
* NET 719 = rl/2.w4 
* NET 720 = rl/1.w1 
* NET 817 = umf.e8 
* NET 818 = umf.e7 
* NET 819 = umf.e6 
* NET 835 = rl/1.e1 
* NET 836 = rl/1.tr_p 
* NET 837 = rl/1.w2 
* NET 838 = rl/1.w3 
* NET 839 = rl/1.w4 
* NET 840 = rl/0.w1 
* NET 961 = umf.e9 
* NET 978 = umf.e12 
* NET 979 = umf.e11 
* NET 980 = umf.e10 
* NET 999 = rck.ck_02 
* NET 1003 = rl/0.e1 
* NET 1004 = rl/0.tr_p 
* NET 1005 = rck.ck_03 
* NET 1006 = rl/0.w2 
* NET 1007 = rl/0.w3 
* NET 1008 = rl/0.w4 
* NET 1137 = umf.e14 
* NET 1138 = umf.e13 
* NET 1139 = umf.e15 
* NET 1152 = rw2.n1 
* NET 1153 = rw3.n1 
* NET 1154 = rw1.n1 
* NET 1155 = rw0.n1 
* NET 1156 = rc116.n2 
* NET 1167 = rp4/15.s3 
* NET 1168 = rmx4/15.bl0_p 
* NET 1169 = rp4/14.s2 
* NET 1170 = rp4/14.s1 
* NET 1171 = rp4/15.s2 
* NET 1172 = rp4/15.s1 
* NET 1173 = rp4/14.s3 
* NET 1174 = rmx4/14.bl0_p 
* NET 1175 = rp4/13.s3 
* NET 1176 = rmx4/13.bl0_p 
* NET 1177 = rp4/12.s2 
* NET 1178 = rp4/13.s2 
* NET 1179 = rp4/12.s3 
* NET 1180 = rp4/12.s1 
* NET 1181 = rp4/13.s1 
* NET 1182 = rp4/11.s3 
* NET 1183 = rmx4/11.bl0_p 
* NET 1184 = rp4/11.s2 
* NET 1185 = rp4/11.s1 
* NET 1186 = rmx4/12.bl0_p 
* NET 1187 = rp4/10.s2 
* NET 1188 = rp4/10.s3 
* NET 1189 = rp4/10.s1 
* NET 1190 = rmx4/10.bl0_p 
* NET 1191 = rp4/9.s3 
* NET 1192 = rmx4/9.bl0_p 
* NET 1193 = rp4/9.s2 
* NET 1194 = rp4/9.s1 
* NET 1195 = rmx4/7.bl0_p 
* NET 1196 = rp4/7.s3 
* NET 1197 = rp4/8.s3 
* NET 1198 = rmx4/8.bl0_p 
* NET 1199 = rp4/8.s2 
* NET 1200 = rp4/8.s1 
* NET 1201 = rp4/6.s2 
* NET 1202 = rp4/6.s1 
* NET 1203 = rp4/7.s2 
* NET 1204 = rp4/7.s1 
* NET 1205 = rp4/5.s3 
* NET 1206 = rmx4/5.bl0_p 
* NET 1207 = rp4/6.s3 
* NET 1208 = rmx4/6.bl0_p 
* NET 1209 = rp4/4.s2 
* NET 1210 = rp4/4.s1 
* NET 1211 = rp4/5.s2 
* NET 1212 = rp4/5.s1 
* NET 1213 = rp4/3.s2 
* NET 1214 = rp4/3.s3 
* NET 1215 = rp4/3.s1 
* NET 1216 = rmx4/3.bl0_p 
* NET 1217 = rp4/4.s3 
* NET 1218 = rmx4/4.bl0_p 
* NET 1219 = rp4/2.s2 
* NET 1220 = rp4/2.s3 
* NET 1221 = rp4/2.s1 
* NET 1222 = rmx4/2.bl0_p 
* NET 1223 = rp4/1.s2 
* NET 1224 = rp4/1.s3 
* NET 1225 = rp4/1.s1 
* NET 1226 = rmx4/1.bl0_p 
* NET 1227 = x0.w2 
* NET 1228 = x0.w1 
* NET 1229 = x0.w0 
* NET 1230 = rp4/0.s2 
* NET 1231 = rp4/0.s3 
* NET 1232 = rp4/0.s1 
* NET 1233 = rmx4/0.bl0_p 
* NET 1234 = ck[0] 
* NET 1241 = rw1.inv 
* NET 1244 = x2.ck_11 
* NET 1246 = x1.w3 
* NET 1247 = rmx4/15.bit_p 
* NET 1248 = rmx4/14.bit_p 
* NET 1249 = rmx4/13.bit_p 
* NET 1250 = rmx4/12.bit_p 
* NET 1251 = rmx4/11.bit_p 
* NET 1252 = rmx4/10.bit_p 
* NET 1253 = rmx4/9.bit_p 
* NET 1254 = rmx4/8.bit_p 
* NET 1255 = rmx4/7.bit_p 
* NET 1256 = rmx4/6.bit_p 
* NET 1257 = rmx4/5.bit_p 
* NET 1258 = rmx4/4.bit_p 
* NET 1259 = rmx4/3.bit_p 
* NET 1260 = rmx4/2.bit_p 
* NET 1261 = rmx4/1.bit_p 
* NET 1262 = x1.ck_13 
* NET 1263 = rmx4/0.bit_p 
* NET 1266 = x2.n3b 
* NET 1268 = rmx2/7.i1 
* NET 1270 = rmx2/7.i0 
* NET 1272 = rmx2/7.s_p 
* NET 1276 = rmx2/6.s_p 
* NET 1278 = rmx2/5.i1 
* NET 1281 = rmx2/5.i0 
* NET 1282 = rmx2/5.s_p 
* NET 1284 = rmx2/3.i1 
* NET 1289 = rmx2/4.s_p 
* NET 1290 = rmx2/3.i0 
* NET 1292 = rmx2/3.s_p 
* NET 1297 = rmx2/1.i1 
* NET 1298 = rmx2/2.s_p 
* NET 1301 = rmx2/1.i0 
* NET 1302 = rmx2/1.s_p 
* NET 1305 = bf.e1 
* NET 1306 = bf.e0 
* NET 1308 = rmx2/0.s_p 
* NET 1318 = adr[7] 
* NET 1319 = rli/0.f 
* NET 1320 = adr[4] 
* NET 1321 = adr[5] 
* NET 1322 = adr[6] 
* NET 1323 = rw3.e1 
* NET 1324 = rli/2.f 
* NET 1325 = rli/1.f 
* NET 1326 = adr[1] 
* NET 1327 = adr[2] 
* NET 1328 = adr[3] 
* NET 1329 = x1.s5 
* NET 1330 = x2.s0 
* NET 1331 = rw3.e3 
* NET 1332 = adr[0] 
* NET 1333 = x0.s7 
* NET 1334 = rob/7.vss1 
* NET 1335 = f[7] 
* NET 1336 = rob/6.vss1 
* NET 1337 = f[6] 
* NET 1338 = rob/5.vss1 
* NET 1339 = f[5] 
* NET 1340 = rob/4.vss1 
* NET 1341 = f[4] 
* NET 1342 = rob/3.vss1 
* NET 1343 = f[3] 
* NET 1344 = rob/2.vss1 
* NET 1345 = f[2] 
* NET 1346 = rob/1.vss1 
* NET 1347 = f[1] 
* NET 1348 = vdd 
* NET 1349 = rob/0.vss1 
* NET 1350 = f[0] 
* NET 1351 = vss 
Mtr_02885 2 1 1348 1348 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02884 999 2 1348 1348 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02883 1348 2 999 1348 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02882 999 2 1348 1348 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02881 1348 999 1005 1348 tp L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02880 1348 1005 3 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02879 1348 3 4 1348 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02878 19 4 1348 1348 tp L=1U W=54U AS=108P AD=108P PS=112U PD=112U 
Mtr_02877 23 1318 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02876 1348 23 21 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02875 23 1321 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02874 20 1351 25 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02873 21 999 20 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02872 1348 1322 23 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02871 26 1005 1348 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02870 1348 5 18 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02869 98 27 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02868 98 27 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02867 1348 18 5 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02866 27 98 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02865 1348 1005 5 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02864 27 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02863 1348 28 99 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02862 100 29 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02861 1348 28 99 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02860 100 29 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02859 1348 1005 28 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02858 29 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02857 29 100 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02856 1348 99 28 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02855 1348 5 18 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02854 105 1318 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02853 1348 105 102 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02852 105 1324 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02851 101 1351 106 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02850 102 999 101 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02849 1348 1322 105 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02848 107 1005 1348 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02847 1348 108 226 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02846 227 109 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02845 227 109 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02844 1348 226 108 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02843 109 227 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02842 1348 1005 108 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02841 109 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02840 1348 110 225 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02839 224 111 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02838 1348 110 225 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02837 224 111 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02836 1348 1005 110 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02835 111 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02834 111 224 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02833 1348 225 110 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02832 1348 108 226 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02831 317 1318 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02830 1348 317 229 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02829 317 1321 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02828 228 1351 318 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02827 229 999 228 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02826 1348 1325 317 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02825 319 1005 1348 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02824 1348 232 312 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02823 313 233 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02822 313 233 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02821 1348 312 232 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02820 233 313 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02819 1348 1005 232 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02818 233 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02817 1348 234 311 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02816 459 320 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02815 1348 234 311 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02814 459 320 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02813 1348 1005 234 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02812 320 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02811 320 459 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02810 1348 311 234 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02809 1348 232 312 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02808 465 1318 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02807 1348 465 315 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02806 465 1324 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02805 314 1351 467 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02804 315 999 314 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02803 1348 1325 465 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02802 468 1005 1348 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02801 1348 321 462 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02800 461 322 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02799 461 322 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02798 1348 462 321 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02797 322 461 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02796 1348 1005 321 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02795 322 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02794 1348 469 460 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02793 558 470 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02792 1348 469 460 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02791 558 470 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02790 1348 1005 469 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02789 470 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02788 470 558 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02787 1348 460 469 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02786 1348 321 462 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02785 570 1319 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02784 1348 570 464 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02783 570 1321 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02782 463 1351 573 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02781 464 999 463 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02780 1348 1322 570 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02779 574 1005 1348 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02778 1348 471 557 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02777 559 472 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02776 559 472 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02775 1348 557 471 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02774 472 559 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02773 1348 1005 471 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02772 472 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02771 1348 575 691 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02770 694 576 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02769 1348 575 691 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02768 694 576 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02767 1348 1005 575 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02766 576 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02765 576 694 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02764 1348 691 575 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02763 1348 471 557 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02762 713 1319 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02761 1348 713 568 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02760 713 1324 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02759 569 1351 716 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02758 568 999 569 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02757 1348 1322 713 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02756 717 1005 1348 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02755 1348 577 693 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02754 692 578 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02753 692 578 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02752 1348 693 577 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02751 578 692 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02750 1348 1005 577 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02749 578 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02748 1348 718 819 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02747 818 719 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02746 1348 718 819 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02745 818 719 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02744 1348 1005 718 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02743 719 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02742 719 818 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02741 1348 819 718 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02740 1348 577 693 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02739 832 1319 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02738 1348 832 711 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02737 832 1321 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02736 712 1351 835 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02735 711 999 712 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02734 1348 1325 832 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02733 836 1005 1348 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02732 1348 720 817 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02731 961 837 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02730 961 837 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02729 1348 817 720 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02728 837 961 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02727 1348 1005 720 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02726 837 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02725 1348 838 980 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02724 979 839 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02723 1348 838 980 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02722 979 839 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02721 1348 1005 838 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02720 839 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02719 839 979 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02718 1348 980 838 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02717 1348 720 817 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02716 1002 1319 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02715 1348 1002 998 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02714 1002 1324 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02713 997 1351 1003 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02712 998 999 997 1348 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02711 1348 1325 1002 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02710 1004 1005 1348 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02709 1348 840 978 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02708 1138 1006 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02707 1138 1006 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02706 1348 978 840 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02705 1006 1138 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02704 1348 1005 840 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02703 1006 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02702 1348 1007 1137 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02701 1139 1008 1348 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02700 1348 1007 1137 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02699 1139 1008 1348 1348 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02698 1348 1005 1007 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02697 1008 1005 1348 1348 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02696 1008 1139 1348 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02695 1348 1137 1007 1348 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02694 1348 840 978 1348 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02693 1244 1234 1348 1348 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02692 1348 1236 1153 1348 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02691 1153 1236 1348 1348 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02690 1236 1320 1348 1348 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02689 1348 1328 1236 1348 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02688 1348 1237 1152 1348 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02687 1152 1237 1348 1348 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02686 1348 1320 1237 1348 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02685 1237 1331 1348 1348 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02684 1348 1241 1154 1348 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02683 1154 1241 1348 1348 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02682 1241 1323 1348 1348 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02681 1348 1328 1241 1348 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02680 1348 1242 1155 1348 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02679 1155 1242 1348 1348 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02678 1348 1323 1242 1348 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02677 1242 1331 1348 1348 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02676 1348 1244 1156 1348 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02675 1262 1156 1348 1348 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02674 1348 1156 1262 1348 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02673 1262 1156 1348 1348 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02672 1348 1156 1262 1348 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02671 1348 1166 1229 1348 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02670 1228 1165 1348 1348 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02669 1348 1244 1165 1348 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02668 1165 1333 1348 1348 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02667 1348 1326 1165 1348 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02666 1166 1332 1348 1348 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02665 1348 1326 1166 1348 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02664 1348 1244 1166 1348 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02663 1348 1243 1227 1348 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02662 1246 1245 1348 1348 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02661 1243 1244 1348 1348 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02660 1243 1332 1348 1348 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02659 1245 1244 1348 1348 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02658 1348 1329 1245 1348 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02657 1245 1333 1348 1348 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02656 1348 1329 1243 1348 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02655 1348 1330 1266 1348 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02654 1266 1244 1348 1348 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02653 1348 1327 1267 1348 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02652 1267 1244 1348 1348 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02651 1306 1266 1348 1348 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02650 1348 1267 1305 1348 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02649 1247 1268 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02648 1348 1262 1247 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02647 1348 1247 1268 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02646 1248 1270 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02645 1348 1262 1248 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02644 1348 1248 1270 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02643 1249 1273 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02642 1348 1262 1249 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02641 1348 1249 1273 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02640 1250 1274 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02639 1348 1262 1250 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02638 1348 1250 1274 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02637 1251 1278 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02636 1348 1262 1251 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02635 1348 1251 1278 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02634 1252 1281 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02633 1348 1262 1252 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02632 1348 1252 1281 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02631 1253 1283 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02630 1348 1262 1253 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02629 1348 1253 1283 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02628 1254 1285 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02627 1348 1262 1254 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02626 1348 1254 1285 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02625 1255 1284 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02624 1348 1262 1255 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02623 1348 1255 1284 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02622 1256 1290 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02621 1348 1262 1256 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02620 1348 1256 1290 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02619 1257 1293 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02618 1348 1262 1257 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02617 1348 1257 1293 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02616 1258 1294 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02615 1348 1262 1258 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02614 1348 1258 1294 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02613 1259 1297 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02612 1348 1262 1259 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02611 1348 1259 1297 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02610 1260 1301 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02609 1348 1262 1260 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02608 1348 1260 1301 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02607 1261 1303 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02606 1348 1262 1261 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02605 1348 1261 1303 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02604 1263 1304 1348 1348 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02603 1348 1262 1263 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02602 1348 1263 1304 1348 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02601 1348 1318 1319 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02600 1319 1318 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02599 1319 1318 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02598 1348 1318 1319 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02597 1319 1318 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02596 1319 1318 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02595 1348 1322 1325 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02594 1325 1322 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02593 1325 1322 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02592 1348 1322 1325 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02591 1325 1322 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02590 1325 1322 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02589 1348 1321 1324 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02588 1324 1321 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02587 1324 1321 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02586 1348 1321 1324 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02585 1324 1321 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02584 1324 1321 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02583 1348 1320 1323 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02582 1323 1320 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02581 1323 1320 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02580 1348 1320 1323 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02579 1323 1320 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02578 1323 1320 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02577 1348 1328 1331 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02576 1331 1328 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02575 1331 1328 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02574 1348 1328 1331 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02573 1331 1328 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02572 1331 1328 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02571 1348 1327 1330 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02570 1330 1327 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02569 1330 1327 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02568 1348 1327 1330 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02567 1330 1327 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02566 1330 1327 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02565 1348 1326 1329 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02564 1329 1326 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02563 1329 1326 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02562 1348 1326 1329 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02561 1329 1326 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02560 1329 1326 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02559 1348 1332 1333 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02558 1333 1332 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02557 1333 1332 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02556 1348 1332 1333 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02555 1333 1332 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02554 1333 1332 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02553 1272 1262 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02552 1272 1310 1348 1348 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02551 1310 1272 1348 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02550 1348 1272 1310 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02549 1348 1334 1335 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02548 1335 1334 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02547 1348 1334 1335 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02546 1348 1334 1335 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02545 1335 1334 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02544 1348 1334 1335 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02543 1348 1310 1334 1348 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02542 1276 1262 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02541 1276 1311 1348 1348 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02540 1311 1276 1348 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02539 1348 1276 1311 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02538 1348 1336 1337 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02537 1337 1336 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02536 1348 1336 1337 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02535 1348 1336 1337 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02534 1337 1336 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02533 1348 1336 1337 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02532 1348 1311 1336 1348 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02531 1282 1262 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02530 1282 1312 1348 1348 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02529 1312 1282 1348 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02528 1348 1282 1312 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02527 1348 1338 1339 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02526 1339 1338 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02525 1348 1338 1339 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02524 1348 1338 1339 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02523 1339 1338 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02522 1348 1338 1339 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02521 1348 1312 1338 1348 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02520 1289 1262 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02519 1289 1313 1348 1348 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02518 1313 1289 1348 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02517 1348 1289 1313 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02516 1348 1340 1341 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02515 1341 1340 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02514 1348 1340 1341 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02513 1348 1340 1341 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02512 1341 1340 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02511 1348 1340 1341 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02510 1348 1313 1340 1348 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02509 1292 1262 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02508 1292 1314 1348 1348 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02507 1314 1292 1348 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02506 1348 1292 1314 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02505 1348 1342 1343 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02504 1343 1342 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02503 1348 1342 1343 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02502 1348 1342 1343 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02501 1343 1342 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02500 1348 1342 1343 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02499 1348 1314 1342 1348 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02498 1298 1262 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02497 1298 1315 1348 1348 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02496 1315 1298 1348 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02495 1348 1298 1315 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02494 1348 1344 1345 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02493 1345 1344 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02492 1348 1344 1345 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02491 1348 1344 1345 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02490 1345 1344 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02489 1348 1344 1345 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02488 1348 1315 1344 1348 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02487 1302 1262 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02486 1302 1316 1348 1348 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02485 1316 1302 1348 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02484 1348 1302 1316 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02483 1348 1346 1347 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02482 1347 1346 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02481 1348 1346 1347 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02480 1348 1346 1347 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02479 1347 1346 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02478 1348 1346 1347 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02477 1348 1316 1346 1348 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02476 1308 1262 1348 1348 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02475 1308 1317 1348 1348 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02474 1317 1308 1348 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02473 1348 1308 1317 1348 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02472 1348 1349 1350 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02471 1350 1349 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02470 1348 1349 1350 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02469 1348 1349 1350 1348 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02468 1350 1349 1348 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02467 1348 1349 1350 1348 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02466 1348 1317 1349 1348 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02465 2 1 1351 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02464 999 2 1351 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02463 1351 2 999 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02462 1351 1005 3 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02461 1005 999 1351 1351 tn L=1U W=18U AS=36P AD=36P PS=40U PD=40U 
Mtr_02460 1351 3 4 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02459 19 4 1351 1351 tn L=1U W=28U AS=56P AD=56P PS=60U PD=60U 
Mtr_02458 1351 1351 25 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02457 23 1321 22 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02456 22 1322 24 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02455 24 1318 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02454 1351 23 25 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02453 25 999 1351 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02452 26 1153 5 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02451 27 1152 26 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02450 26 1154 28 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02449 29 1155 26 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02448 1351 25 26 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02447 26 25 1351 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02446 1351 5 18 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02445 98 27 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02444 1351 28 99 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02443 100 29 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02442 1351 1351 106 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02441 105 1324 103 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02440 103 1322 104 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02439 104 1318 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02438 1351 105 106 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02437 106 999 1351 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02436 107 1153 108 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02435 109 1152 107 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02434 107 1154 110 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02433 111 1155 107 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02432 1351 106 107 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02431 107 106 1351 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02430 1351 108 226 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02429 227 109 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02428 1351 110 225 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02427 224 111 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02426 1351 1351 318 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02425 317 1321 231 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02424 231 1325 230 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02423 230 1318 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02422 1351 317 318 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02421 318 999 1351 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02420 319 1153 232 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02419 233 1152 319 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02418 319 1154 234 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02417 320 1155 319 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02416 1351 318 319 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02415 319 318 1351 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02414 1351 232 312 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02413 313 233 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02412 1351 234 311 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02411 459 320 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02410 1351 1351 467 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02409 465 1324 466 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02408 466 1325 316 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02407 316 1318 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02406 1351 465 467 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02405 467 999 1351 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02404 468 1153 321 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02403 322 1152 468 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02402 468 1154 469 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02401 470 1155 468 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02400 1351 467 468 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02399 468 467 1351 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02398 1351 321 462 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02397 461 322 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02396 1351 469 460 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02395 558 470 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02394 1351 1351 573 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02393 570 1321 571 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02392 571 1322 572 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02391 572 1319 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02390 1351 570 573 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02389 573 999 1351 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02388 574 1153 471 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02387 472 1152 574 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02386 574 1154 575 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02385 576 1155 574 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02384 1351 573 574 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02383 574 573 1351 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02382 1351 471 557 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02381 559 472 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02380 1351 575 691 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02379 694 576 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02378 1351 1351 716 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02377 713 1324 715 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02376 715 1322 714 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02375 714 1319 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02374 1351 713 716 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02373 716 999 1351 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02372 717 1153 577 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02371 578 1152 717 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02370 717 1154 718 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02369 719 1155 717 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02368 1351 716 717 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02367 717 716 1351 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02366 1351 577 693 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02365 692 578 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02364 1351 718 819 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02363 818 719 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02362 1351 1351 835 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02361 832 1321 833 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02360 833 1325 834 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02359 834 1319 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02358 1351 832 835 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02357 835 999 1351 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02356 836 1153 720 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02355 837 1152 836 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02354 836 1154 838 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02353 839 1155 836 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02352 1351 835 836 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02351 836 835 1351 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02350 1351 720 817 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02349 961 837 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02348 1351 838 980 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02347 979 839 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02346 1351 1351 1003 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02345 1002 1324 1000 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02344 1000 1325 1001 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02343 1001 1319 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02342 1351 1002 1003 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02341 1003 999 1351 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02340 1004 1153 840 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02339 1006 1152 1004 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02338 1004 1154 1007 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02337 1008 1155 1004 1351 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02336 1351 1003 1004 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02335 1004 1003 1351 1351 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02334 1351 840 978 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02333 1138 1006 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02332 1351 1007 1137 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02331 1139 1008 1351 1351 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02330 1351 1234 1244 1351 tn L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02329 1153 1236 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02328 1351 1236 1153 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02327 1236 1328 1235 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02326 1235 1320 1351 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02325 1152 1237 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02324 1351 1237 1152 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02323 1238 1331 1237 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02322 1351 1320 1238 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02321 1154 1241 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02320 1351 1241 1154 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02319 1240 1323 1351 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02318 1241 1328 1240 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02317 1351 1242 1155 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02316 1239 1331 1242 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02315 1351 1323 1239 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02314 1155 1242 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02313 1156 1244 1351 1351 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02312 1351 1156 1262 1351 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02311 1262 1156 1351 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02310 1163 1244 1165 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02309 1164 1333 1163 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02308 1351 1326 1164 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02307 1228 1165 1351 1351 tn L=1U W=26U AS=52P AD=52P PS=56U PD=56U 
Mtr_02306 1161 1244 1166 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02305 1162 1332 1161 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02304 1351 1326 1162 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02303 1351 1166 1229 1351 tn L=1U W=26U AS=52P AD=52P PS=56U PD=56U 
Mtr_02302 1159 1244 1351 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02301 1160 1329 1159 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02300 1243 1332 1160 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02299 1351 1243 1227 1351 tn L=1U W=26U AS=52P AD=52P PS=56U PD=56U 
Mtr_02298 1246 1245 1351 1351 tn L=1U W=26U AS=52P AD=52P PS=56U PD=56U 
Mtr_02297 1157 1244 1351 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02296 1158 1329 1157 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02295 1245 1333 1158 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02294 1266 1330 1264 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02293 1264 1244 1351 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02292 1306 1266 1351 1351 tn L=1U W=18U AS=36P AD=36P PS=40U PD=40U 
Mtr_02291 1351 1267 1305 1351 tn L=1U W=18U AS=36P AD=36P PS=40U PD=40U 
Mtr_02290 1267 1327 1265 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02289 1265 1244 1351 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02288 1168 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02287 1167 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02286 1171 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02285 1172 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02284 127 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02283 1171 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02282 1351 226 125 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02281 1351 226 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02280 40 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02279 1171 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02278 1351 99 41 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02277 1351 99 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02276 1351 18 9 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02275 1351 18 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02274 39 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02273 1171 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02272 115 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02271 1351 226 112 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02270 32 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02269 1351 99 30 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02268 31 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02267 1351 18 6 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02266 1168 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02265 1351 226 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02264 1168 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02263 1351 99 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02262 1168 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02261 1351 18 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02260 245 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02259 1171 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02258 1351 312 246 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02257 1351 312 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02256 1171 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02255 126 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02254 1351 225 124 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02253 1351 225 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02252 1351 225 114 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02251 113 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02250 1351 312 235 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02249 237 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02248 1351 225 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02247 1168 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02246 1351 312 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02245 1168 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02244 1351 311 244 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02243 1351 311 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02242 337 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02241 1171 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02240 1351 311 236 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02239 1351 311 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02238 323 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02237 1168 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02236 1351 462 338 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02235 1351 462 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02234 1351 462 326 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02233 1351 462 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02232 336 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02231 1171 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02230 325 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02229 1168 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02228 484 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02227 1351 460 335 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02226 1171 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02225 1351 460 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02224 475 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02223 1351 460 324 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02222 1351 460 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02221 1168 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02220 594 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02219 1171 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02218 1351 693 592 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02217 1351 693 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02216 593 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02215 1171 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02214 1351 691 590 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02213 1351 691 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02212 1351 557 483 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02211 1351 557 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02210 482 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02209 1171 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02208 582 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02207 1351 693 580 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02206 581 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02205 1351 691 579 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02204 473 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02203 1351 557 474 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02202 1168 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02201 1351 693 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02200 1168 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02199 1351 691 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02198 1168 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02197 1351 557 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02196 855 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02195 1171 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02194 1351 817 732 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02193 1351 817 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02192 1171 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02191 730 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02190 1351 819 731 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02189 1351 819 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02188 1351 819 721 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02187 723 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02186 1351 817 722 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02185 841 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02184 1351 819 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02183 1168 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02182 1351 817 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02181 1168 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02180 1351 980 856 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02179 1351 980 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02178 854 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02177 1171 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02176 1351 980 844 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02175 1351 980 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02174 843 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02173 1168 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02172 1351 978 853 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02171 1351 978 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02170 1351 978 842 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02169 1351 978 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02168 1019 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02167 1171 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02166 1009 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02165 1168 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02164 1020 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02163 1351 1137 1018 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02162 1171 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02161 1351 1137 1171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02160 1010 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02159 1351 1137 1011 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02158 1351 1137 1168 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02157 1168 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02156 1247 1229 1168 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02155 1351 1247 1268 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02154 1171 1227 1247 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02153 1247 1246 1172 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02152 1247 1228 1167 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02151 1174 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02150 1173 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02149 1169 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02148 1170 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02147 123 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02146 1169 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02145 1351 226 118 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02144 1351 226 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02143 35 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02142 1169 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02141 1351 99 37 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02140 1351 99 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02139 1351 18 8 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02138 1351 18 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02137 33 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02136 1169 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02135 119 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02134 1351 226 116 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02133 36 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02132 1351 99 38 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02131 34 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02130 1351 18 7 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02129 1174 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02128 1351 226 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02127 1174 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02126 1351 99 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02125 1174 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02124 1351 18 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02123 238 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02122 1169 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02121 1351 312 240 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02120 1351 312 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02119 1169 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02118 120 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02117 1351 225 122 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02116 1351 225 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02115 1351 225 117 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02114 121 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02113 1351 312 241 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02112 239 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02111 1351 225 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02110 1174 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02109 1351 312 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02108 1174 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02107 1351 311 242 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02106 1351 311 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02105 329 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02104 1169 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02103 1351 311 243 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02102 1351 311 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02101 330 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02100 1174 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02099 1351 462 327 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02098 1351 462 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02097 1351 462 328 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02096 1351 462 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02095 333 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02094 1169 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02093 334 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02092 1174 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02091 480 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02090 1351 460 331 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02089 1169 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02088 1351 460 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02087 481 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02086 1351 460 332 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02085 1351 460 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02084 1174 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02083 591 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02082 1169 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02081 1351 693 587 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02080 1351 693 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02079 589 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02078 1169 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02077 1351 691 584 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02076 1351 691 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02075 1351 557 477 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02074 1351 557 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02073 479 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02072 1169 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02071 586 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02070 1351 693 588 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02069 585 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02068 1351 691 583 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02067 476 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02066 1351 557 478 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02065 1174 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02064 1351 693 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02063 1174 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02062 1351 691 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02061 1174 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02060 1351 557 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02059 847 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02058 1169 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02057 1351 817 728 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02056 1351 817 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02055 1169 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02054 724 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02053 1351 819 726 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02052 1351 819 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02051 1351 819 727 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02050 725 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02049 1351 817 729 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02048 848 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02047 1351 819 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02046 1174 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02045 1351 817 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02044 1174 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02043 1351 980 845 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02042 1351 980 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02041 851 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02040 1169 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02039 1351 980 846 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02038 1351 980 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02037 852 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02036 1174 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02035 1351 978 849 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02034 1351 978 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02033 1351 978 850 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02032 1351 978 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02031 1016 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02030 1169 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02029 1012 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02028 1174 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02027 1017 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02026 1351 1137 1014 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02025 1169 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02024 1351 1137 1169 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02023 1013 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02022 1351 1137 1015 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02021 1351 1137 1174 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02020 1174 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02019 1248 1229 1174 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02018 1351 1248 1270 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02017 1169 1227 1248 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02016 1248 1246 1170 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02015 1248 1228 1173 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02014 1176 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02013 1175 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02012 1178 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02011 1181 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02010 143 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02009 130 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02008 1351 226 141 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02007 1351 226 129 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02006 52 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02005 43 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02004 1351 99 53 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02003 1351 99 44 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02002 1351 18 13 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02001 1351 18 10 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02000 51 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01999 42 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01998 1175 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01997 1351 226 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01996 1175 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01995 1351 99 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01994 1175 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01993 1351 18 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01992 1176 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01991 1351 226 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01990 1176 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01989 1351 99 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01988 1176 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01987 1351 18 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01986 257 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01985 248 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01984 1351 312 258 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01983 1351 312 249 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01982 131 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01981 142 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01980 1351 225 140 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01979 1351 225 128 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01978 1351 225 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01977 1175 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01976 1351 312 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01975 1175 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01974 1351 225 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01973 1176 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01972 1351 312 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01971 1176 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01970 1351 311 256 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01969 1351 311 247 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01968 353 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01967 341 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01966 1351 311 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01965 1351 311 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01964 1175 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01963 1176 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01962 1351 462 354 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01961 1351 462 340 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01960 1351 462 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01959 1351 462 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01958 352 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01957 339 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01956 1175 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01955 1176 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01954 496 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01953 1351 460 351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01952 487 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01951 1351 460 342 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01950 1175 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01949 1351 460 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01948 1351 460 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01947 1176 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01946 610 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01945 597 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01944 1351 693 608 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01943 1351 693 598 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01942 609 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01941 596 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01940 1351 691 605 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01939 1351 691 595 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01938 1351 557 495 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01937 1351 557 485 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01936 494 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01935 486 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01934 1175 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01933 1351 693 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01932 1175 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01931 1351 691 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01930 1175 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01929 1351 557 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01928 1176 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01927 1351 693 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01926 1176 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01925 1351 691 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01924 1176 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01923 1351 557 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01922 871 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01921 859 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01920 1351 817 744 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01919 1351 817 733 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01918 734 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01917 742 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01916 1351 819 743 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01915 1351 819 735 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01914 1351 819 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01913 1175 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01912 1351 817 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01911 1175 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01910 1351 819 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01909 1176 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01908 1351 817 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01907 1176 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01906 1351 980 872 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01905 1351 980 858 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01904 870 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01903 857 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01902 1351 980 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01901 1351 980 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01900 1175 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01899 1176 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01898 1351 978 869 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01897 1351 978 860 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01896 1351 978 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01895 1351 978 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01894 1031 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01893 1021 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01892 1175 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01891 1176 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01890 1032 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01889 1351 1137 1030 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01888 1022 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01887 1351 1137 1023 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01886 1175 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01885 1351 1137 1175 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01884 1351 1137 1176 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01883 1176 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01882 1249 1229 1176 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01881 1351 1249 1273 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01880 1178 1227 1249 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01879 1249 1246 1181 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01878 1249 1228 1175 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01877 1186 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01876 1179 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01875 1177 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01874 1180 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01873 138 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01872 139 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01871 1351 226 133 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01870 1351 226 132 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01869 47 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01868 48 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01867 1351 99 49 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01866 1351 99 50 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01865 1351 18 11 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01864 1351 18 12 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01863 45 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01862 46 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01861 1179 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01860 1351 226 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01859 1179 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01858 1351 99 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01857 1179 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01856 1351 18 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01855 1186 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01854 1351 226 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01853 1186 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01852 1351 99 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01851 1186 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01850 1351 18 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01849 250 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01848 251 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01847 1351 312 252 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01846 1351 312 253 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01845 135 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01844 134 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01843 1351 225 136 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01842 1351 225 137 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01841 1351 225 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01840 1179 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01839 1351 312 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01838 1179 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01837 1351 225 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01836 1186 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01835 1351 312 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01834 1186 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01833 1351 311 254 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01832 1351 311 255 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01831 345 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01830 346 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01829 1351 311 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01828 1351 311 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01827 1179 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01826 1186 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01825 1351 462 343 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01824 1351 462 344 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01823 1351 462 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01822 1351 462 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01821 349 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01820 350 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01819 1179 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01818 1186 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01817 492 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01816 1351 460 347 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01815 493 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01814 1351 460 348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01813 1179 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01812 1351 460 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01811 1351 460 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01810 1186 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01809 606 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01808 607 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01807 1351 693 601 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01806 1351 693 602 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01805 603 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01804 604 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01803 1351 691 600 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01802 1351 691 599 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01801 1351 557 488 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01800 1351 557 489 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01799 490 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01798 491 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01797 1179 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01796 1351 693 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01795 1179 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01794 1351 691 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01793 1179 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01792 1351 557 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01791 1186 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01790 1351 693 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01789 1186 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01788 1351 691 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01787 1186 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01786 1351 557 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01785 863 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01784 864 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01783 1351 817 740 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01782 1351 817 741 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01781 737 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01780 736 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01779 1351 819 738 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01778 1351 819 739 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01777 1351 819 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01776 1179 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01775 1351 817 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01774 1179 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01773 1351 819 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01772 1186 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01771 1351 817 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01770 1186 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01769 1351 980 861 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01768 1351 980 862 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01767 867 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01766 868 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01765 1351 980 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01764 1351 980 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01763 1179 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01762 1186 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01761 1351 978 865 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01760 1351 978 866 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01759 1351 978 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01758 1351 978 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01757 1026 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01756 1027 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01755 1179 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01754 1186 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01753 1028 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01752 1351 1137 1024 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01751 1029 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01750 1351 1137 1025 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01749 1179 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01748 1351 1137 1179 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01747 1351 1137 1186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01746 1186 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01745 1250 1229 1186 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01744 1351 1250 1274 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01743 1177 1227 1250 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01742 1250 1246 1180 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01741 1250 1228 1179 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01740 1183 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01739 1182 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01738 1184 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01737 1185 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01736 159 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01735 151 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01734 1351 226 150 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01733 1351 226 145 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01732 59 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01731 60 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01730 1351 99 63 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01729 1351 99 64 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01728 1351 18 16 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01727 1351 18 17 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01726 55 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01725 56 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01724 152 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01723 1351 226 146 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01722 61 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01721 1351 99 65 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01720 57 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01719 1351 18 14 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01718 153 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01717 1351 226 144 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01716 62 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01715 1351 99 54 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01714 58 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01713 1351 18 15 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01712 259 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01711 260 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01710 1351 312 263 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01709 1351 312 264 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01708 155 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01707 154 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01706 1351 225 158 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01705 1351 225 147 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01704 1351 225 148 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01703 156 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01702 1351 312 265 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01701 261 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01700 1351 225 149 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01699 157 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01698 1351 312 266 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01697 262 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01696 1351 311 267 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01695 1351 311 268 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01694 359 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01693 360 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01692 1351 311 269 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01691 1351 311 270 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01690 361 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01689 362 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01688 1351 462 355 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01687 1351 462 356 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01686 1351 462 357 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01685 1351 462 358 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01684 367 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01683 368 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01682 369 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01681 370 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01680 506 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01679 1351 460 363 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01678 507 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01677 1351 460 364 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01676 508 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01675 1351 460 365 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01674 1351 460 366 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01673 505 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01672 626 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01671 618 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01670 1351 693 621 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01669 1351 693 622 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01668 625 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01667 615 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01666 1351 691 614 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01665 1351 691 613 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01664 1351 557 500 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01663 1351 557 501 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01662 504 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01661 497 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01660 619 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01659 1351 693 623 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01658 616 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01657 1351 691 612 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01656 498 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01655 1351 557 502 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01654 620 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01653 1351 693 624 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01652 617 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01651 1351 691 611 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01650 499 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01649 1351 557 503 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01648 877 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01647 878 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01646 1351 817 753 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01645 1351 817 754 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01644 746 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01643 745 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01642 1351 819 749 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01641 1351 819 750 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01640 1351 819 751 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01639 747 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01638 1351 817 755 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01637 879 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01636 1351 819 752 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01635 748 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01634 1351 817 756 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01633 880 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01632 1351 980 873 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01631 1351 980 874 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01630 885 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01629 886 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01628 1351 980 875 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01627 1351 980 876 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01626 887 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01625 888 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01624 1351 978 881 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01623 1351 978 882 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01622 1351 978 883 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01621 1351 978 884 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01620 1037 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01619 1034 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01618 1035 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01617 1036 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01616 1038 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01615 1351 1137 1042 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01614 1039 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01613 1351 1137 1043 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01612 1040 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01611 1351 1137 1044 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01610 1351 1137 1033 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01609 1041 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01608 1251 1229 1183 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01607 1351 1251 1278 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01606 1184 1227 1251 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01605 1251 1246 1185 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01604 1251 1228 1182 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01603 1190 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01602 1188 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01601 1187 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01600 1189 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01599 1189 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01598 1187 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01597 1351 226 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01596 1351 226 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01595 1189 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01594 1187 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01593 1351 99 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01592 1351 99 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01591 1351 18 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01590 1351 18 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01589 1189 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01588 1187 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01587 1188 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01586 1351 226 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01585 1188 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01584 1351 99 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01583 1188 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01582 1351 18 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01581 1190 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01580 1351 226 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01579 1190 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01578 1351 99 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01577 1190 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01576 1351 18 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01575 1189 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01574 1187 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01573 1351 312 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01572 1351 312 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01571 1187 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01570 1189 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01569 1351 225 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01568 1351 225 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01567 1351 225 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01566 1188 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01565 1351 312 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01564 1188 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01563 1351 225 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01562 1190 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01561 1351 312 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01560 1190 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01559 1351 311 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01558 1351 311 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01557 1189 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01556 1187 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01555 1351 311 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01554 1351 311 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01553 1188 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01552 1190 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01551 1351 462 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01550 1351 462 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01549 1351 462 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01548 1351 462 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01547 1189 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01546 1187 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01545 1188 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01544 1190 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01543 1189 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01542 1351 460 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01541 1187 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01540 1351 460 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01539 1188 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01538 1351 460 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01537 1351 460 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01536 1190 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01535 1189 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01534 1187 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01533 1351 693 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01532 1351 693 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01531 1189 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01530 1187 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01529 1351 691 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01528 1351 691 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01527 1351 557 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01526 1351 557 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01525 1189 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01524 1187 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01523 1188 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01522 1351 693 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01521 1188 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01520 1351 691 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01519 1188 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01518 1351 557 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01517 1190 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01516 1351 693 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01515 1190 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01514 1351 691 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01513 1190 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01512 1351 557 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01511 1189 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01510 1187 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01509 1351 817 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01508 1351 817 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01507 1187 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01506 1189 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01505 1351 819 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01504 1351 819 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01503 1351 819 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01502 1188 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01501 1351 817 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01500 1188 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01499 1351 819 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01498 1190 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01497 1351 817 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01496 1190 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01495 1351 980 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01494 1351 980 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01493 1189 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01492 1187 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01491 1351 980 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01490 1351 980 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01489 1188 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01488 1190 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01487 1351 978 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01486 1351 978 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01485 1351 978 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01484 1351 978 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01483 1189 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01482 1187 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01481 1188 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01480 1190 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01479 1189 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01478 1351 1137 1189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01477 1187 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01476 1351 1137 1187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01475 1188 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01474 1351 1137 1188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01473 1351 1137 1190 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01472 1190 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01471 1252 1229 1190 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01470 1351 1252 1281 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01469 1187 1227 1252 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01468 1252 1246 1189 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01467 1252 1228 1188 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01466 1192 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01465 1191 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01464 1193 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01463 1194 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01462 160 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01461 161 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01460 1351 226 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01459 1351 226 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01458 73 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01457 69 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01456 1351 99 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01455 1351 99 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01454 1351 18 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01453 1351 18 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01452 72 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01451 66 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01450 162 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01449 1351 226 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01448 70 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01447 1351 99 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01446 67 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01445 1351 18 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01444 163 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01443 1351 226 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01442 71 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01441 1351 99 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01440 68 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01439 1351 18 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01438 273 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01437 274 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01436 1351 312 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01435 1351 312 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01434 165 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01433 164 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01432 1351 225 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01431 1351 225 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01430 1351 225 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01429 166 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01428 1351 312 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01427 271 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01426 1351 225 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01425 167 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01424 1351 312 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01423 272 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01422 1351 311 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01421 1351 311 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01420 373 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01419 374 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01418 1351 311 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01417 1351 311 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01416 371 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01415 372 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01414 1351 462 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01413 1351 462 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01412 1351 462 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01411 1351 462 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01410 375 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01409 376 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01408 377 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01407 378 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01406 513 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01405 1351 460 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01404 514 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01403 1351 460 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01402 515 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01401 1351 460 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01400 1351 460 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01399 516 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01398 631 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01397 632 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01396 1351 693 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01395 1351 693 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01394 627 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01393 628 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01392 1351 691 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01391 1351 691 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01390 1351 557 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01389 1351 557 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01388 510 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01387 511 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01386 633 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01385 1351 693 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01384 629 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01383 1351 691 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01382 512 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01381 1351 557 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01380 634 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01379 1351 693 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01378 630 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01377 1351 691 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01376 509 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01375 1351 557 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01374 891 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01373 892 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01372 1351 817 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01371 1351 817 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01370 760 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01369 759 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01368 1351 819 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01367 1351 819 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01366 1351 819 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01365 757 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01364 1351 817 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01363 889 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01362 1351 819 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01361 758 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01360 1351 817 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01359 890 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01358 1351 980 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01357 1351 980 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01356 893 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01355 894 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01354 1351 980 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01353 1351 980 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01352 895 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01351 896 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01350 1351 978 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01349 1351 978 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01348 1351 978 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01347 1351 978 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01346 1048 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01345 1045 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01344 1046 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01343 1047 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01342 1049 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01341 1351 1137 1194 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01340 1050 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01339 1351 1137 1193 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01338 1051 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01337 1351 1137 1191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01336 1351 1137 1192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01335 1052 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01334 1253 1229 1192 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01333 1351 1253 1283 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01332 1193 1227 1253 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01331 1253 1246 1194 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01330 1253 1228 1191 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01329 1198 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01328 1197 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01327 1199 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01326 1200 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01325 176 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01324 177 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01323 1351 226 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01322 1351 226 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01321 82 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01320 83 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01319 1351 99 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01318 1351 99 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01317 1351 18 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01316 1351 18 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01315 78 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01314 79 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01313 178 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01312 1351 226 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01311 84 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01310 1351 99 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01309 80 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01308 1351 18 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01307 179 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01306 1351 226 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01305 85 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01304 1351 99 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01303 81 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01302 1351 18 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01301 277 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01300 278 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01299 1351 312 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01298 1351 312 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01297 173 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01296 172 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01295 1351 225 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01294 1351 225 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01293 1351 225 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01292 174 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01291 1351 312 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01290 279 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01289 1351 225 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01288 175 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01287 1351 312 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01286 280 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01285 1351 311 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01284 1351 311 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01283 383 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01282 384 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01281 1351 311 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01280 1351 311 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01279 385 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01278 386 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01277 1351 462 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01276 1351 462 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01275 1351 462 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01274 1351 462 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01273 387 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01272 388 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01271 389 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01270 390 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01269 525 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01268 1351 460 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01267 526 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01266 1351 460 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01265 524 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01264 1351 460 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01263 1351 460 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01262 523 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01261 643 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01260 644 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01259 1351 693 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01258 1351 693 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01257 639 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01256 640 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01255 1351 691 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01254 1351 691 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01253 1351 557 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01252 1351 557 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01251 522 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01250 519 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01249 645 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01248 1351 693 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01247 641 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01246 1351 691 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01245 520 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01244 1351 557 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01243 646 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01242 1351 693 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01241 642 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01240 1351 691 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01239 521 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01238 1351 557 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01237 901 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01236 902 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01235 1351 817 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01234 1351 817 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01233 766 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01232 765 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01231 1351 819 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01230 1351 819 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01229 1351 819 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01228 767 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01227 1351 817 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01226 903 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01225 1351 819 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01224 768 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01223 1351 817 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01222 904 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01221 1351 980 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01220 1351 980 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01219 905 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01218 906 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01217 1351 980 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01216 1351 980 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01215 907 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01214 908 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01213 1351 978 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01212 1351 978 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01211 1351 978 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01210 1351 978 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01209 1059 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01208 1060 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01207 1057 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01206 1058 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01205 1061 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01204 1351 1137 1200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01203 1062 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01202 1351 1137 1199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01201 1063 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01200 1351 1137 1197 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01199 1351 1137 1198 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01198 1064 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01197 1254 1229 1198 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01196 1351 1254 1285 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01195 1199 1227 1254 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01194 1254 1246 1200 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01193 1254 1228 1197 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01192 1195 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01191 1196 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01190 1203 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01189 1204 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01188 1204 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01187 1203 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01186 1351 226 1204 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01185 1351 226 1203 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01184 91 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01183 92 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01182 1351 99 93 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01181 1351 99 90 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01180 1351 18 1204 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01179 1351 18 1203 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01178 1204 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01177 1203 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01176 1196 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01175 1351 226 1196 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01174 76 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01173 1351 99 74 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01172 1196 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01171 1351 18 1196 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01170 1195 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01169 1351 226 1195 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01168 77 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01167 1351 99 75 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01166 1195 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01165 1351 18 1195 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01164 1204 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01163 1203 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01162 1351 312 1204 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01161 1351 312 1203 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01160 185 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01159 184 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01158 1351 225 186 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01157 1351 225 187 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01156 1351 225 170 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01155 168 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01154 1351 312 1196 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01153 1196 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01152 1351 225 171 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01151 169 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01150 1351 312 1195 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01149 1195 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01148 1351 311 283 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01147 1351 311 284 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01146 395 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01145 396 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01144 1351 311 275 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01143 1351 311 276 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01142 379 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01141 380 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01140 1351 462 1204 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01139 1351 462 1203 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01138 1351 462 1196 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01137 1351 462 1195 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01136 1204 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01135 1203 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01134 1196 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01133 1195 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01132 530 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01131 1351 460 397 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01130 529 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01129 1351 460 398 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01128 518 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01127 1351 460 381 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01126 1351 460 382 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01125 517 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01124 1204 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01123 1203 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01122 1351 693 1204 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01121 1351 693 1203 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01120 654 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01119 653 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01118 1351 691 651 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01117 1351 691 652 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01116 1351 557 1204 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01115 1351 557 1203 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01114 1204 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01113 1203 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01112 1196 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01111 1351 693 1196 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01110 637 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01109 1351 691 636 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01108 1196 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01107 1351 557 1196 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01106 1195 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01105 1351 693 1195 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01104 638 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01103 1351 691 635 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01102 1195 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01101 1351 557 1195 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01100 1204 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01099 1203 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01098 1351 817 1204 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01097 1351 817 1203 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01096 774 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01095 773 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01094 1351 819 775 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01093 1351 819 776 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01092 1351 819 762 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01091 763 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01090 1351 817 1196 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01089 1196 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01088 1351 819 761 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01087 764 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01086 1351 817 1195 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01085 1195 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01084 1351 980 915 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01083 1351 980 916 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01082 913 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01081 914 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01080 1351 980 899 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01079 1351 980 900 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01078 897 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01077 898 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01076 1351 978 1204 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01075 1351 978 1203 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01074 1351 978 1196 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01073 1351 978 1195 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01072 1204 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01071 1203 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01070 1196 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01069 1195 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01068 1069 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01067 1351 1137 1071 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01066 1070 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01065 1351 1137 1072 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01064 1055 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01063 1351 1137 1053 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01062 1351 1137 1054 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01061 1056 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01060 1255 1229 1195 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01059 1351 1255 1284 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01058 1203 1227 1255 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01057 1255 1246 1204 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01056 1255 1228 1196 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01055 1208 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01054 1207 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01053 1201 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01052 1202 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01051 1202 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01050 1201 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01049 1351 226 1202 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01048 1351 226 1201 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01047 86 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01046 87 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01045 1351 99 88 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01044 1351 99 89 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01043 1351 18 1202 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01042 1351 18 1201 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01041 1202 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01040 1201 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01039 1207 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01038 1351 226 1207 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01037 94 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01036 1351 99 96 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01035 1207 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01034 1351 18 1207 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01033 1208 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01032 1351 226 1208 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01031 95 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01030 1351 99 97 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01029 1208 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01028 1351 18 1208 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01027 1202 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01026 1201 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01025 1351 312 1202 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01024 1351 312 1201 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01023 183 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01022 182 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01021 1351 225 180 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01020 1351 225 181 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01019 1351 225 199 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01018 197 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01017 1351 312 1207 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01016 1207 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01015 1351 225 196 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01014 198 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01013 1351 312 1208 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01012 1208 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01011 1351 311 281 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01010 1351 311 282 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01009 391 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01008 392 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01007 1351 311 285 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01006 1351 311 286 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01005 408 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01004 405 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01003 1351 462 1202 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01002 1351 462 1201 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01001 1351 462 1207 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01000 1351 462 1208 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00999 1202 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00998 1201 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00997 1207 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00996 1208 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00995 527 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00994 1351 460 393 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00993 528 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00992 1351 460 394 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00991 533 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00990 1351 460 406 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00989 1351 460 407 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00988 534 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00987 1202 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00986 1201 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00985 1351 693 1202 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00984 1351 693 1201 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00983 649 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00982 650 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00981 1351 691 647 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00980 1351 691 648 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00979 1351 557 1202 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00978 1351 557 1201 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00977 1202 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00976 1201 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00975 1207 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00974 1351 693 1207 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00973 661 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00972 1351 691 660 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00971 1207 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00970 1351 557 1207 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00969 1208 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00968 1351 693 1208 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00967 662 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00966 1351 691 658 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00965 1208 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00964 1351 557 1208 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00963 1202 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00962 1201 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00961 1351 817 1202 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00960 1351 817 1201 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00959 770 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00958 769 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00957 1351 819 771 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00956 1351 819 772 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00955 1351 819 784 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00954 781 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00953 1351 817 1207 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00952 1207 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00951 1351 819 783 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00950 782 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00949 1351 817 1208 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00948 1208 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00947 1351 980 909 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00946 1351 980 910 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00945 911 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00944 912 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00943 1351 980 922 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00942 1351 980 919 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00941 920 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00940 921 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00939 1351 978 1202 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00938 1351 978 1201 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00937 1351 978 1207 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00936 1351 978 1208 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00935 1202 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00934 1201 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00933 1207 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00932 1208 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00931 1065 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00930 1351 1137 1067 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00929 1066 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00928 1351 1137 1068 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00927 1080 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00926 1351 1137 1082 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00925 1351 1137 1079 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00924 1081 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00923 1256 1229 1208 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00922 1351 1256 1290 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00921 1201 1227 1256 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00920 1256 1246 1202 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00919 1256 1228 1207 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00918 1206 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00917 1205 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00916 1211 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00915 1212 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00914 217 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00913 218 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00912 1351 226 216 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00911 1351 226 212 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00910 1212 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00909 1211 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00908 1351 99 1212 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00907 1351 99 1211 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00906 1351 18 1212 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00905 1351 18 1211 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00904 1212 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00903 1211 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00902 193 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00901 1351 226 188 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00900 1205 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00899 1351 99 1205 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00898 1205 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00897 1351 18 1205 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00896 194 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00895 1351 226 189 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00894 1206 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00893 1351 99 1206 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00892 1206 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00891 1351 18 1206 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00890 1212 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00889 1211 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00888 1351 312 1212 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00887 1351 312 1211 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00886 213 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00885 219 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00884 1351 225 214 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00883 1351 225 215 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00882 1351 225 191 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00881 195 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00880 1351 312 1205 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00879 1205 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00878 1351 225 192 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00877 190 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00876 1351 312 1206 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00875 1206 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00874 1351 311 1212 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00873 1351 311 1211 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00872 1212 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00871 1211 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00870 1351 311 1205 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00869 1351 311 1206 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00868 1205 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00867 1206 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00866 1351 462 423 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00865 1351 462 418 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00864 1351 462 400 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00863 1351 462 401 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00862 421 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00861 422 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00860 404 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00859 399 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00858 538 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00857 1351 460 419 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00856 539 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00855 1351 460 420 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00854 532 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00853 1351 460 402 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00852 1351 460 403 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00851 531 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00850 672 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00849 669 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00848 1351 693 670 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00847 1351 693 671 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00846 1212 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00845 1211 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00844 1351 691 1212 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00843 1351 691 1211 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00842 1351 557 1212 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00841 1351 557 1211 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00840 1212 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00839 1211 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00838 659 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00837 1351 693 656 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00836 1205 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00835 1351 691 1205 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00834 1205 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00833 1351 557 1205 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00832 655 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00831 1351 693 657 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00830 1206 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00829 1351 691 1206 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00828 1206 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00827 1351 557 1206 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00826 1212 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00825 1211 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00824 1351 817 1212 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00823 1351 817 1211 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00822 792 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00821 791 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00820 1351 819 793 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00819 1351 819 794 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00818 1351 819 778 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00817 780 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00816 1351 817 1205 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00815 1205 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00814 1351 819 779 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00813 777 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00812 1351 817 1206 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00811 1206 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00810 1351 980 1212 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00809 1351 980 1211 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00808 1212 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00807 1211 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00806 1351 980 1205 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00805 1351 980 1206 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00804 1205 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00803 1206 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00802 1351 978 926 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00801 1351 978 927 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00800 1351 978 917 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00799 1351 978 918 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00798 1096 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00797 1095 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00796 1073 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00795 1074 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00794 1097 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00793 1351 1137 1093 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00792 1092 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00791 1351 1137 1094 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00790 1075 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00789 1351 1137 1077 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00788 1351 1137 1078 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00787 1076 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00786 1257 1229 1206 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00785 1351 1257 1293 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00784 1211 1227 1257 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00783 1257 1246 1212 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00782 1257 1228 1205 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00781 1218 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00780 1217 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00779 1209 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00778 1210 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00777 211 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00776 203 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00775 1351 226 201 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00774 1351 226 202 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00773 1210 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00772 1209 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00771 1351 99 1210 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00770 1351 99 1209 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00769 1351 18 1210 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00768 1351 18 1209 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00767 1210 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00766 1209 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00765 204 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00764 1351 226 200 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00763 1217 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00762 1351 99 1217 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00761 1217 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00760 1351 18 1217 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00759 223 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00758 1351 226 220 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00757 1218 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00756 1351 99 1218 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00755 1218 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00754 1351 18 1218 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00753 1210 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00752 1209 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00751 1351 312 1210 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00750 1351 312 1209 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00749 206 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00748 205 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00747 1351 225 208 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00746 1351 225 209 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00745 1351 225 210 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00744 207 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00743 1351 312 1217 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00742 1217 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00741 1351 225 222 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00740 221 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00739 1351 312 1218 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00738 1218 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00737 1351 311 1210 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00736 1351 311 1209 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00735 1210 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00734 1209 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00733 1351 311 1217 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00732 1351 311 1218 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00731 1217 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00730 1218 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00729 1351 462 414 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00728 1351 462 415 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00727 1351 462 416 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00726 1351 462 442 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00725 411 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00724 412 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00723 413 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00722 441 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00721 536 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00720 1351 460 417 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00719 537 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00718 1351 460 409 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00717 535 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00716 1351 460 410 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00715 1351 460 440 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00714 544 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00713 663 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00712 664 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00711 1351 693 666 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00710 1351 693 667 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00709 1210 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00708 1209 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00707 1351 691 1210 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00706 1351 691 1209 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00705 1351 557 1210 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00704 1351 557 1209 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00703 1210 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00702 1209 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00701 665 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00700 1351 693 668 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00699 1217 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00698 1351 691 1217 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00697 1217 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00696 1351 557 1217 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00695 673 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00694 1351 693 674 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00693 1218 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00692 1351 691 1218 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00691 1218 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00690 1351 557 1218 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00689 1210 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00688 1209 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00687 1351 817 1210 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00686 1351 817 1209 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00685 786 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00684 785 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00683 1351 819 788 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00682 1351 819 789 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00681 1351 819 790 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00680 787 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00679 1351 817 1217 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00678 1217 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00677 1351 819 799 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00676 800 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00675 1351 817 1218 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00674 1218 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00673 1351 980 1210 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00672 1351 980 1209 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00671 1210 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00670 1209 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00669 1351 980 1217 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00668 1351 980 1218 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00667 1217 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00666 1218 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00665 1351 978 923 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00664 1351 978 924 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00663 1351 978 925 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00662 1351 978 944 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00661 1088 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00660 1086 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00659 1087 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00658 1111 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00657 1089 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00656 1351 1137 1083 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00655 1090 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00654 1351 1137 1084 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00653 1091 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00652 1351 1137 1085 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00651 1351 1137 1112 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00650 1110 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00649 1258 1229 1218 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00648 1351 1258 1294 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00647 1209 1227 1258 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00646 1258 1246 1210 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00645 1258 1228 1217 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00644 1216 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00643 1214 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00642 1213 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00641 1215 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00640 1215 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00639 1213 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00638 1351 226 1215 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00637 1351 226 1213 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00636 1215 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00635 1213 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00634 1351 99 1215 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00633 1351 99 1213 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00632 1351 18 1215 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00631 1351 18 1213 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00630 1215 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00629 1213 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00628 1214 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00627 1351 226 1214 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00626 1214 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00625 1351 99 1214 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00624 1214 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00623 1351 18 1214 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00622 1216 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00621 1351 226 1216 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00620 1216 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00619 1351 99 1216 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00618 1216 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00617 1351 18 1216 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00616 295 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00615 296 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00614 1351 312 287 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00613 1351 312 288 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00612 1213 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00611 1215 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00610 1351 225 1215 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00609 1351 225 1213 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00608 1351 225 1214 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00607 1214 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00606 1351 312 289 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00605 297 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00604 1351 225 1216 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00603 1216 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00602 1351 312 290 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00601 298 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00600 1351 311 291 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00599 1351 311 292 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00598 430 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00597 427 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00596 1351 311 293 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00595 1351 311 294 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00594 428 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00593 429 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00592 1351 462 438 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00591 1351 462 424 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00590 1351 462 425 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00589 1351 462 426 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00588 434 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00587 435 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00586 436 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00585 437 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00584 541 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00583 1351 460 439 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00582 542 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00581 1351 460 431 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00580 543 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00579 1351 460 432 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00578 1351 460 433 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00577 540 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00576 1215 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00575 1213 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00574 1351 693 1215 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00573 1351 693 1213 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00572 1215 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00571 1213 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00570 1351 691 1215 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00569 1351 691 1213 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00568 1351 557 1215 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00567 1351 557 1213 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00566 1215 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00565 1213 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00564 1214 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00563 1351 693 1214 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00562 1214 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00561 1351 691 1214 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00560 1214 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00559 1351 557 1214 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00558 1216 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00557 1351 693 1216 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00556 1216 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00555 1351 691 1216 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00554 1216 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00553 1351 557 1216 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00552 930 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00551 931 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00550 1351 817 795 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00549 1351 817 796 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00548 1213 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00547 1215 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00546 1351 819 1215 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00545 1351 819 1213 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00544 1351 819 1214 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00543 1214 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00542 1351 817 797 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00541 932 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00540 1351 819 1216 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00539 1216 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00538 1351 817 798 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00537 929 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00536 1351 980 938 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00535 1351 980 939 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00534 934 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00533 935 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00532 1351 980 940 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00531 1351 980 928 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00530 936 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00529 937 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00528 1351 978 941 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00527 1351 978 942 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00526 1351 978 943 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00525 1351 978 933 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00524 1102 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00523 1103 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00522 1104 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00521 1105 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00520 1106 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00519 1351 1137 1098 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00518 1107 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00517 1351 1137 1099 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00516 1108 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00515 1351 1137 1100 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00514 1351 1137 1101 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00513 1109 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00512 1259 1229 1216 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00511 1351 1259 1297 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00510 1213 1227 1259 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00509 1259 1246 1215 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00508 1259 1228 1214 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00507 1222 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00506 1220 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00505 1219 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00504 1221 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00503 1221 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00502 1219 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00501 1351 226 1221 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00500 1351 226 1219 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00499 1221 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00498 1219 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00497 1351 99 1221 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00496 1351 99 1219 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00495 1351 18 1221 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00494 1351 18 1219 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00493 1221 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00492 1219 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00491 1220 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00490 1351 226 1220 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00489 1220 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00488 1351 99 1220 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00487 1220 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00486 1351 18 1220 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00485 1222 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00484 1351 226 1222 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00483 1222 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00482 1351 99 1222 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00481 1222 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00480 1351 18 1222 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00479 299 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00478 300 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00477 1351 312 303 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00476 1351 312 304 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00475 1219 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00474 1221 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00473 1351 225 1221 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00472 1351 225 1219 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00471 1351 225 1220 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00470 1220 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00469 1351 312 305 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00468 301 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00467 1351 225 1222 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00466 1222 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00465 1351 312 306 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00464 302 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00463 1351 311 307 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00462 1351 311 308 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00461 447 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00460 448 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00459 1351 311 309 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00458 1351 311 310 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00457 449 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00456 450 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00455 1351 462 443 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00454 1351 462 444 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00453 1351 462 445 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00452 1351 462 446 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00451 455 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00450 456 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00449 457 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00448 458 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00447 547 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00446 1351 460 451 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00445 548 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00444 1351 460 452 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00443 545 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00442 1351 460 453 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00441 1351 460 454 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00440 546 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00439 1221 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00438 1219 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00437 1351 693 1221 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00436 1351 693 1219 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00435 1221 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00434 1219 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00433 1351 691 1221 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00432 1351 691 1219 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00431 1351 557 1221 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00430 1351 557 1219 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00429 1221 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00428 1219 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00427 1220 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00426 1351 693 1220 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00425 1220 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00424 1351 691 1220 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00423 1220 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00422 1351 557 1220 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00421 1222 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00420 1351 693 1222 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00419 1222 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00418 1351 691 1222 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00417 1222 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00416 1351 557 1222 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00415 949 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00414 950 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00413 1351 817 801 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00412 1351 817 802 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00411 1219 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00410 1221 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00409 1351 819 1221 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00408 1351 819 1219 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00407 1351 819 1220 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00406 1220 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00405 1351 817 803 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00404 951 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00403 1351 819 1222 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00402 1222 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00401 1351 817 804 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00400 952 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00399 1351 980 945 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00398 1351 980 946 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00397 957 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00396 958 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00395 1351 980 947 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00394 1351 980 948 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00393 959 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00392 960 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00391 1351 978 953 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00390 1351 978 954 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00389 1351 978 955 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00388 1351 978 956 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00387 1117 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00386 1118 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00385 1119 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00384 1120 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00383 1121 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00382 1351 1137 1113 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00381 1122 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00380 1351 1137 1114 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00379 1123 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00378 1351 1137 1115 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00377 1351 1137 1116 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00376 1124 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00375 1260 1229 1222 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00374 1351 1260 1301 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00373 1219 1227 1260 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00372 1260 1246 1221 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00371 1260 1228 1220 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00370 1226 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00369 1224 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00368 1223 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00367 1225 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00366 1225 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00365 1223 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00364 1351 226 1225 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00363 1351 226 1223 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00362 1225 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00361 1223 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00360 1351 99 1225 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00359 1351 99 1223 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00358 1351 18 1225 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00357 1351 18 1223 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00356 1225 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00355 1223 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00354 1224 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00353 1351 226 1224 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00352 1224 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00351 1351 99 1224 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00350 1224 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00349 1351 18 1224 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00348 1226 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00347 1351 226 1226 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00346 1226 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00345 1351 99 1226 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00344 1226 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00343 1351 18 1226 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00342 1225 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00341 1223 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00340 1351 312 1225 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00339 1351 312 1223 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00338 1223 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00337 1225 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00336 1351 225 1225 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00335 1351 225 1223 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00334 1351 225 1224 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00333 1224 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00332 1351 312 1224 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00331 1224 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00330 1351 225 1226 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00329 1226 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00328 1351 312 1226 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00327 1226 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00326 1351 311 1225 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00325 1351 311 1223 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00324 1225 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00323 1223 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00322 1351 311 1224 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00321 1351 311 1226 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00320 1224 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00319 1226 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00318 1351 462 1225 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00317 1351 462 1223 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00316 1351 462 1224 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00315 1351 462 1226 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00314 1225 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00313 1223 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00312 1224 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00311 1226 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00310 1225 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00309 1351 460 1225 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00308 1223 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00307 1351 460 1223 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00306 1224 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00305 1351 460 1224 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00304 1351 460 1226 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00303 1226 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00302 683 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00301 684 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00300 1351 693 687 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00299 1351 693 688 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00298 679 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00297 680 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00296 1351 691 677 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00295 1351 691 678 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00294 1351 557 551 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00293 1351 557 552 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00292 555 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00291 556 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00290 685 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00289 1351 693 689 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00288 681 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00287 1351 691 676 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00286 549 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00285 1351 557 553 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00284 686 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00283 1351 693 690 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00282 682 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00281 1351 691 675 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00280 550 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00279 1351 557 554 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00278 962 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00277 963 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00276 1351 817 809 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00275 1351 817 810 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00274 814 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00273 813 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00272 1351 819 805 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00271 1351 819 806 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00270 1351 819 807 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00269 815 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00268 1351 817 811 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00267 964 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00266 1351 819 808 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00265 816 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00264 1351 817 812 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00263 965 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00262 1351 980 970 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00261 1351 980 971 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00260 966 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00259 967 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00258 1351 980 972 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00257 1351 980 973 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00256 968 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00255 969 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00254 1351 978 974 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00253 1351 978 975 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00252 1351 978 976 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00251 1351 978 977 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00250 1127 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00249 1128 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00248 1125 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00247 1126 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00246 1129 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00245 1351 1137 1133 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00244 1130 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00243 1351 1137 1134 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00242 1131 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00241 1351 1137 1135 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00240 1351 1137 1136 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00239 1132 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00238 1261 1229 1226 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00237 1351 1261 1303 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00236 1223 1227 1261 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00235 1261 1246 1225 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00234 1261 1228 1224 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00233 1233 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00232 1231 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00231 1230 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00230 1232 19 1348 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00229 1232 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00228 1230 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00227 1351 226 1232 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00226 1351 226 1230 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00225 1232 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00224 1230 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00223 1351 99 1232 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00222 1351 99 1230 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00221 1351 18 1232 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00220 1351 18 1230 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00219 1232 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00218 1230 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00217 1231 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00216 1351 226 1231 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00215 1231 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00214 1351 99 1231 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00213 1231 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00212 1351 18 1231 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00211 1233 227 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00210 1351 226 1233 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00209 1233 100 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00208 1351 99 1233 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00207 1233 98 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00206 1351 18 1233 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00205 1232 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00204 1230 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00203 1351 312 1232 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00202 1351 312 1230 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00201 1230 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00200 1232 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00199 1351 225 1232 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00198 1351 225 1230 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00197 1351 225 1231 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00196 1231 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00195 1351 312 1231 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00194 1231 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00193 1351 225 1233 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00192 1233 224 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00191 1351 312 1233 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00190 1233 313 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00189 1351 311 1232 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00188 1351 311 1230 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00187 1232 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00186 1230 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00185 1351 311 1231 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00184 1351 311 1233 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00183 1231 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00182 1233 459 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00181 1351 462 1232 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00180 1351 462 1230 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00179 1351 462 1231 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00178 1351 462 1233 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00177 1232 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00176 1230 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00175 1231 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00174 1233 461 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00173 1232 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00172 1351 460 1232 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00171 1230 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00170 1351 460 1230 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00169 1231 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00168 1351 460 1231 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00167 1351 460 1233 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00166 1233 558 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00165 707 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00164 708 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00163 1351 693 699 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00162 1351 693 700 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00161 703 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00160 704 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00159 1351 691 697 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00158 1351 691 698 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00157 1351 557 566 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00156 1351 557 567 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00155 562 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00154 563 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00153 709 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00152 1351 693 701 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00151 705 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00150 1351 691 696 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00149 564 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00148 1351 557 560 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00147 710 692 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00146 1351 693 702 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00145 706 694 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00144 1351 691 695 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00143 565 559 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00142 1351 557 561 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00141 985 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00140 986 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00139 1351 817 828 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00138 1351 817 829 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00137 821 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00136 820 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00135 1351 819 824 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00134 1351 819 825 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00133 1351 819 826 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00132 822 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00131 1351 817 830 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00130 987 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00129 1351 819 827 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00128 823 818 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00127 1351 817 831 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00126 988 961 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00125 1351 980 981 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00124 1351 980 982 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00123 993 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00122 994 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00121 1351 980 983 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00120 1351 980 984 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00119 995 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00118 996 979 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00117 1351 978 989 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00116 1351 978 990 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00115 1351 978 991 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00114 1351 978 992 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00113 1144 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00112 1145 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00111 1146 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00110 1147 1138 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00109 1148 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00108 1351 1137 1140 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00107 1149 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00106 1351 1137 1141 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00105 1150 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00104 1351 1137 1142 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00103 1351 1137 1143 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00102 1151 1139 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00101 1263 1229 1233 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00100 1351 1263 1304 1351 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00099 1230 1227 1263 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00098 1263 1246 1232 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00097 1263 1228 1231 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00096 1351 1318 1319 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00095 1319 1318 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00094 1319 1318 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00093 1351 1322 1325 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00092 1325 1322 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00091 1325 1322 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00090 1351 1321 1324 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00089 1324 1321 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00088 1324 1321 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00087 1351 1320 1323 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00086 1323 1320 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00085 1323 1320 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00084 1351 1328 1331 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00083 1331 1328 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00082 1331 1328 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00081 1351 1327 1330 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00080 1330 1327 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00079 1330 1327 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00078 1351 1326 1329 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00077 1329 1326 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00076 1329 1326 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00075 1351 1332 1333 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00074 1333 1332 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00073 1333 1332 1351 1351 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00072 1351 1270 1271 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00071 1271 1305 1272 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00070 1272 1306 1269 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00069 1269 1268 1351 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00068 1310 1272 1351 1351 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00067 1335 1334 1351 1351 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00066 1351 1334 1335 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00065 1351 1310 1334 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00064 1335 1334 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00063 1351 1274 1277 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00062 1277 1305 1276 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00061 1276 1306 1275 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00060 1275 1273 1351 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00059 1311 1276 1351 1351 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00058 1337 1336 1351 1351 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00057 1351 1336 1337 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00056 1351 1311 1336 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00055 1337 1336 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00054 1351 1281 1280 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00053 1280 1305 1282 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00052 1282 1306 1279 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00051 1279 1278 1351 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00050 1312 1282 1351 1351 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00049 1339 1338 1351 1351 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00048 1351 1338 1339 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00047 1351 1312 1338 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00046 1339 1338 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00045 1351 1285 1288 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00044 1288 1305 1289 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00043 1289 1306 1287 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00042 1287 1283 1351 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00041 1313 1289 1351 1351 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00040 1341 1340 1351 1351 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00039 1351 1340 1341 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00038 1351 1313 1340 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00037 1341 1340 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00036 1351 1290 1291 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00035 1291 1305 1292 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00034 1292 1306 1286 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00033 1286 1284 1351 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00032 1314 1292 1351 1351 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00031 1343 1342 1351 1351 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00030 1351 1342 1343 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00029 1351 1314 1342 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00028 1343 1342 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00027 1351 1294 1296 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00026 1296 1305 1298 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00025 1298 1306 1295 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00024 1295 1293 1351 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00023 1315 1298 1351 1351 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00022 1345 1344 1351 1351 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00021 1351 1344 1345 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00020 1351 1315 1344 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00019 1345 1344 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00018 1351 1301 1299 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00017 1299 1305 1302 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00016 1302 1306 1300 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00015 1300 1297 1351 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00014 1316 1302 1351 1351 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00013 1347 1346 1351 1351 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00012 1351 1346 1347 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 1351 1316 1346 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00010 1347 1346 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 1351 1304 1309 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00008 1309 1305 1308 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00007 1308 1306 1307 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00006 1307 1303 1351 1351 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00005 1317 1308 1351 1351 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00004 1350 1349 1351 1351 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00003 1351 1349 1350 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 1351 1317 1349 1351 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00001 1350 1349 1351 1351 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
.ends r256x8_1

