* Spice description of ram4x128
* Spice driver version 700
* Date ( dd/mm/yyyy hh:mm:ss ): 10/09/2002 at 18:56:47

* INTERF write vss vdd en dout[3] dout[2] dout[1] dout[0] ck adr[6] adr[5] 
* INTERF adr[4] adr[3] adr[2] adr[1] adr[0] 


.subckt ram4x128 1578 1579 1580 1581 1582 1583 1584 1585 1586 1587 1588 1589 
+ 1590 1591 1592 1593 
* net 1 = mbk_sig129 
* net 2 = mbk_sig135 
* net 3 = mbk_sig139 
* net 4 = mbk_sig140 
* net 5 = mbk_sig87 
* net 6 = mbk_sig104 
* net 7 = mbk_sig125 
* net 8 = mbk_sig1 
* net 9 = mbk_sig3 
* net 10 = mbk_sig132 
* net 11 = mbk_sig136 
* net 12 = mbk_sig142 
* net 13 = mbk_sig141 
* net 14 = mbk_sig90 
* net 15 = mbk_sig106 
* net 16 = mbk_sig126 
* net 17 = mbk_sig9 
* net 18 = mbk_sig10 
* net 19 = mbk_sig1591 
* net 20 = mbk_sig1589 
* net 21 = mbk_sig1577 
* net 22 = mbk_sig1575 
* net 23 = mbk_sig1544 
* net 24 = mbk_sig1576 
* net 25 = mbk_sig1543 
* net 26 = mbk_sig1542 
* net 27 = mbk_sig1512 
* net 28 = mbk_sig1511 
* net 29 = mbk_sig1573 
* net 30 = mbk_sig1541 
* net 31 = mbk_sig1486 
* net 32 = mbk_sig1487 
* net 33 = mbk_sig1466 
* net 34 = mbk_sig1465 
* net 35 = mbk_sig1443 
* net 36 = mbk_sig1440 
* net 37 = mbk_sig1441 
* net 38 = mbk_sig1442 
* net 39 = mbk_sig1463 
* net 40 = mbk_sig1437 
* net 41 = mbk_sig1407 
* net 42 = mbk_sig1408 
* net 43 = mbk_sig1377 
* net 44 = mbk_sig1376 
* net 45 = mbk_sig1353 
* net 46 = mbk_sig1352 
* net 47 = mbk_sig1329 
* net 48 = mbk_sig1328 
* net 49 = mbk_sig1374 
* net 50 = mbk_sig1349 
* net 51 = mbk_sig1307 
* net 52 = mbk_sig1304 
* net 53 = mbk_sig1305 
* net 54 = mbk_sig1306 
* net 55 = mbk_sig1272 
* net 56 = mbk_sig1273 
* net 57 = mbk_sig1240 
* net 58 = mbk_sig1241 
* net 59 = mbk_sig1302 
* net 60 = mbk_sig1271 
* net 61 = mbk_sig1217 
* net 62 = mbk_sig1216 
* net 63 = mbk_sig1196 
* net 64 = mbk_sig1195 
* net 65 = mbk_sig1165 
* net 66 = mbk_sig1162 
* net 67 = mbk_sig1163 
* net 68 = mbk_sig1164 
* net 69 = mbk_sig1193 
* net 70 = mbk_sig1159 
* net 71 = mbk_sig1128 
* net 72 = mbk_sig1129 
* net 73 = mbk_sig1106 
* net 74 = mbk_sig1107 
* net 75 = mbk_sig1083 
* net 76 = mbk_sig1082 
* net 77 = mbk_sig1058 
* net 78 = mbk_sig1059 
* net 79 = mbk_sig1104 
* net 80 = mbk_sig1079 
* net 81 = mbk_sig1027 
* net 82 = mbk_sig1057 
* net 83 = mbk_sig1026 
* net 84 = mbk_sig1025 
* net 85 = mbk_sig994 
* net 86 = mbk_sig993 
* net 87 = mbk_sig969 
* net 88 = mbk_sig970 
* net 89 = mbk_sig1023 
* net 90 = mbk_sig991 
* net 91 = mbk_sig947 
* net 92 = mbk_sig946 
* net 93 = mbk_sig925 
* net 94 = mbk_sig926 
* net 95 = mbk_sig893 
* net 96 = mbk_sig924 
* net 97 = mbk_sig892 
* net 98 = mbk_sig891 
* net 99 = mbk_sig922 
* net 100 = mbk_sig887 
* net 101 = mbk_sig856 
* net 102 = mbk_sig857 
* net 103 = mbk_sig836 
* net 104 = mbk_sig837 
* net 105 = mbk_sig813 
* net 106 = mbk_sig812 
* net 107 = mbk_sig788 
* net 108 = mbk_sig789 
* net 109 = mbk_sig834 
* net 110 = mbk_sig809 
* net 111 = mbk_sig786 
* net 112 = mbk_sig787 
* net 113 = mbk_sig755 
* net 114 = mbk_sig756 
* net 115 = mbk_sig723 
* net 116 = mbk_sig724 
* net 117 = mbk_sig699 
* net 118 = mbk_sig698 
* net 119 = mbk_sig753 
* net 120 = mbk_sig720 
* net 121 = mbk_sig677 
* net 122 = mbk_sig675 
* net 123 = mbk_sig644 
* net 124 = mbk_sig676 
* net 125 = mbk_sig643 
* net 126 = mbk_sig642 
* net 127 = mbk_sig612 
* net 128 = mbk_sig611 
* net 129 = mbk_sig673 
* net 130 = mbk_sig641 
* net 131 = mbk_sig586 
* net 132 = mbk_sig587 
* net 133 = mbk_sig566 
* net 134 = mbk_sig565 
* net 135 = mbk_sig543 
* net 136 = mbk_sig541 
* net 137 = mbk_sig542 
* net 138 = mbk_sig509 
* net 139 = mbk_sig563 
* net 140 = mbk_sig538 
* net 141 = mbk_sig507 
* net 142 = mbk_sig508 
* net 143 = mbk_sig477 
* net 144 = mbk_sig476 
* net 145 = mbk_sig454 
* net 146 = mbk_sig453 
* net 147 = mbk_sig429 
* net 148 = mbk_sig428 
* net 149 = mbk_sig474 
* net 150 = mbk_sig450 
* net 151 = mbk_sig406 
* net 152 = mbk_sig407 
* net 153 = mbk_sig404 
* net 154 = mbk_sig405 
* net 155 = mbk_sig372 
* net 156 = mbk_sig373 
* net 157 = mbk_sig341 
* net 158 = mbk_sig340 
* net 159 = mbk_sig402 
* net 160 = mbk_sig371 
* net 161 = mbk_sig317 
* net 162 = mbk_sig316 
* net 163 = mbk_sig296 
* net 164 = mbk_sig295 
* net 165 = mbk_sig273 
* net 166 = mbk_sig270 
* net 167 = mbk_sig271 
* net 168 = mbk_sig272 
* net 169 = mbk_sig293 
* net 170 = mbk_sig267 
* net 171 = mbk_sig237 
* net 172 = mbk_sig238 
* net 173 = mbk_sig206 
* net 174 = mbk_sig207 
* net 175 = mbk_sig183 
* net 176 = mbk_sig182 
* net 177 = mbk_sig159 
* net 178 = mbk_sig158 
* net 179 = mbk_sig204 
* net 180 = mbk_sig179 
* net 181 = mbk_sig77 
* net 182 = mbk_sig79 
* net 183 = mbk_sig92 
* net 184 = mbk_sig91 
* net 185 = mbk_sig48 
* net 186 = mbk_sig52 
* net 187 = mbk_sig44 
* net 188 = mbk_sig41 
* net 189 = mbk_sig18 
* net 190 = mbk_sig133 
* net 191 = mbk_sig137 
* net 192 = mbk_sig143 
* net 193 = mbk_sig144 
* net 194 = mbk_sig97 
* net 195 = mbk_sig112 
* net 196 = mbk_sig127 
* net 197 = mbk_sig31 
* net 198 = mbk_sig30 
* net 199 = mbk_sig134 
* net 200 = mbk_sig138 
* net 201 = mbk_sig145 
* net 202 = mbk_sig146 
* net 203 = mbk_sig99 
* net 204 = mbk_sig114 
* net 205 = mbk_sig128 
* net 206 = mbk_sig35 
* net 207 = mbk_sig37 
* net 208 = rbit_0_0.ram_63_1.m0_s 
* net 209 = rbit_0_0.ram_63_1.m1_s 
* net 210 = rbit_0_0.ram_63_0.m0_s 
* net 211 = rbit_0_0.ram_63_0.m1_s 
* net 212 = rbit_0_0.ram_62_1.m0_s 
* net 213 = rbit_0_0.ram_62_1.m1_s 
* net 214 = rbit_0_0.ram_62_0.m0_s 
* net 215 = rbit_0_0.ram_62_0.m1_s 
* net 216 = rbit_0_0.ram_61_1.m0_s 
* net 217 = rbit_0_0.ram_61_1.m1_s 
* net 218 = rbit_0_0.ram_61_0.m0_s 
* net 219 = rbit_0_0.ram_61_0.m1_s 
* net 220 = rbit_0_0.ram_60_1.m0_s 
* net 221 = rbit_0_0.ram_60_1.m1_s 
* net 222 = rbit_0_0.ram_60_0.m0_s 
* net 223 = rbit_0_0.ram_60_0.m1_s 
* net 224 = rbit_0_0.ram_59_1.m0_s 
* net 225 = rbit_0_0.ram_59_1.m1_s 
* net 226 = rbit_0_0.ram_59_0.m0_s 
* net 227 = rbit_0_0.ram_59_0.m1_s 
* net 228 = rbit_0_0.ram_58_1.m0_s 
* net 229 = rbit_0_0.ram_58_1.m1_s 
* net 230 = rbit_0_0.ram_58_0.m0_s 
* net 231 = rbit_0_0.ram_58_0.m1_s 
* net 232 = rbit_0_0.ram_57_1.m0_s 
* net 233 = rbit_0_0.ram_57_1.m1_s 
* net 234 = rbit_0_0.ram_57_0.m0_s 
* net 235 = rbit_0_0.ram_57_0.m1_s 
* net 236 = rbit_0_0.ram_56_1.m0_s 
* net 237 = rbit_0_0.ram_56_1.m1_s 
* net 238 = rbit_0_0.ram_56_0.m0_s 
* net 239 = rbit_0_0.ram_56_0.m1_s 
* net 240 = rbit_0_0.ram_55_1.m0_s 
* net 241 = rbit_0_0.ram_55_1.m1_s 
* net 242 = rbit_0_0.ram_55_0.m0_s 
* net 243 = rbit_0_0.ram_55_0.m1_s 
* net 244 = rbit_0_0.ram_54_1.m0_s 
* net 245 = rbit_0_0.ram_54_1.m1_s 
* net 246 = rbit_0_0.ram_54_0.m0_s 
* net 247 = rbit_0_0.ram_54_0.m1_s 
* net 248 = rbit_0_0.ram_53_1.m0_s 
* net 249 = rbit_0_0.ram_53_1.m1_s 
* net 250 = rbit_0_0.ram_53_0.m0_s 
* net 251 = rbit_0_0.ram_53_0.m1_s 
* net 252 = rbit_0_0.ram_52_1.m0_s 
* net 253 = rbit_0_0.ram_52_1.m1_s 
* net 254 = rbit_0_0.ram_52_0.m0_s 
* net 255 = rbit_0_0.ram_52_0.m1_s 
* net 256 = rbit_0_0.ram_51_1.m0_s 
* net 257 = rbit_0_0.ram_51_1.m1_s 
* net 258 = rbit_0_0.ram_51_0.m0_s 
* net 259 = rbit_0_0.ram_51_0.m1_s 
* net 260 = rbit_0_0.ram_50_1.m0_s 
* net 261 = rbit_0_0.ram_50_1.m1_s 
* net 262 = rbit_0_0.ram_50_0.m0_s 
* net 263 = rbit_0_0.ram_50_0.m1_s 
* net 264 = rbit_0_0.ram_49_1.m0_s 
* net 265 = rbit_0_0.ram_49_1.m1_s 
* net 266 = rbit_0_0.ram_49_0.m0_s 
* net 267 = rbit_0_0.ram_49_0.m1_s 
* net 268 = rbit_0_0.ram_48_1.m0_s 
* net 269 = rbit_0_0.ram_48_1.m1_s 
* net 270 = rbit_0_0.ram_48_0.m0_s 
* net 271 = rbit_0_0.ram_48_0.m1_s 
* net 272 = rbit_0_0.ram_47_1.m0_s 
* net 273 = rbit_0_0.ram_47_1.m1_s 
* net 274 = rbit_0_0.ram_47_0.m0_s 
* net 275 = rbit_0_0.ram_47_0.m1_s 
* net 276 = rbit_0_0.ram_46_1.m0_s 
* net 277 = rbit_0_0.ram_46_1.m1_s 
* net 278 = rbit_0_0.ram_46_0.m0_s 
* net 279 = rbit_0_0.ram_46_0.m1_s 
* net 280 = rbit_0_0.ram_45_1.m0_s 
* net 281 = rbit_0_0.ram_45_1.m1_s 
* net 282 = rbit_0_0.ram_45_0.m0_s 
* net 283 = rbit_0_0.ram_45_0.m1_s 
* net 284 = rbit_0_0.ram_44_1.m0_s 
* net 285 = rbit_0_0.ram_44_1.m1_s 
* net 286 = rbit_0_0.ram_44_0.m0_s 
* net 287 = rbit_0_0.ram_44_0.m1_s 
* net 288 = rbit_0_0.ram_43_1.m0_s 
* net 289 = rbit_0_0.ram_43_1.m1_s 
* net 290 = rbit_0_0.ram_43_0.m0_s 
* net 291 = rbit_0_0.ram_43_0.m1_s 
* net 292 = rbit_0_0.ram_42_1.m0_s 
* net 293 = rbit_0_0.ram_42_1.m1_s 
* net 294 = rbit_0_0.ram_42_0.m0_s 
* net 295 = rbit_0_0.ram_42_0.m1_s 
* net 296 = rbit_0_0.ram_41_1.m0_s 
* net 297 = rbit_0_0.ram_41_1.m1_s 
* net 298 = rbit_0_0.ram_41_0.m0_s 
* net 299 = rbit_0_0.ram_41_0.m1_s 
* net 300 = rbit_0_0.ram_40_1.m0_s 
* net 301 = rbit_0_0.ram_40_1.m1_s 
* net 302 = rbit_0_0.ram_40_0.m0_s 
* net 303 = rbit_0_0.ram_40_0.m1_s 
* net 304 = rbit_0_0.ram_39_1.m0_s 
* net 305 = rbit_0_0.ram_39_1.m1_s 
* net 306 = rbit_0_0.ram_39_0.m0_s 
* net 307 = rbit_0_0.ram_39_0.m1_s 
* net 308 = rbit_0_0.ram_38_1.m0_s 
* net 309 = rbit_0_0.ram_38_1.m1_s 
* net 310 = rbit_0_0.ram_38_0.m0_s 
* net 311 = rbit_0_0.ram_38_0.m1_s 
* net 312 = rbit_0_0.ram_37_1.m0_s 
* net 313 = rbit_0_0.ram_37_1.m1_s 
* net 314 = rbit_0_0.ram_37_0.m0_s 
* net 315 = rbit_0_0.ram_37_0.m1_s 
* net 316 = rbit_0_0.ram_36_1.m0_s 
* net 317 = rbit_0_0.ram_36_1.m1_s 
* net 318 = rbit_0_0.ram_36_0.m0_s 
* net 319 = rbit_0_0.ram_36_0.m1_s 
* net 320 = rbit_0_0.ram_35_1.m0_s 
* net 321 = rbit_0_0.ram_35_1.m1_s 
* net 322 = rbit_0_0.ram_35_0.m0_s 
* net 323 = rbit_0_0.ram_35_0.m1_s 
* net 324 = rbit_0_0.ram_34_1.m0_s 
* net 325 = rbit_0_0.ram_34_1.m1_s 
* net 326 = rbit_0_0.ram_34_0.m0_s 
* net 327 = rbit_0_0.ram_34_0.m1_s 
* net 328 = rbit_0_0.ram_33_1.m0_s 
* net 329 = rbit_0_0.ram_33_1.m1_s 
* net 330 = rbit_0_0.ram_33_0.m0_s 
* net 331 = rbit_0_0.ram_33_0.m1_s 
* net 332 = rbit_0_0.ram_32_1.m0_s 
* net 333 = rbit_0_0.ram_32_1.m1_s 
* net 334 = rbit_0_0.ram_32_0.m0_s 
* net 335 = rbit_0_0.ram_32_0.m1_s 
* net 336 = rbit_0_0.ram_31_1.m0_s 
* net 337 = rbit_0_0.ram_31_1.m1_s 
* net 338 = rbit_0_0.ram_31_0.m0_s 
* net 339 = rbit_0_0.ram_31_0.m1_s 
* net 340 = rbit_0_0.ram_30_1.m0_s 
* net 341 = rbit_0_0.ram_30_1.m1_s 
* net 342 = rbit_0_0.ram_30_0.m0_s 
* net 343 = rbit_0_0.ram_30_0.m1_s 
* net 344 = rbit_0_0.ram_29_1.m0_s 
* net 345 = rbit_0_0.ram_29_1.m1_s 
* net 346 = rbit_0_0.ram_29_0.m0_s 
* net 347 = rbit_0_0.ram_29_0.m1_s 
* net 348 = rbit_0_0.ram_28_1.m0_s 
* net 349 = rbit_0_0.ram_28_1.m1_s 
* net 350 = rbit_0_0.ram_28_0.m0_s 
* net 351 = rbit_0_0.ram_28_0.m1_s 
* net 352 = rbit_0_0.ram_27_1.m0_s 
* net 353 = rbit_0_0.ram_27_1.m1_s 
* net 354 = rbit_0_0.ram_27_0.m0_s 
* net 355 = rbit_0_0.ram_27_0.m1_s 
* net 356 = rbit_0_0.ram_26_1.m0_s 
* net 357 = rbit_0_0.ram_26_1.m1_s 
* net 358 = rbit_0_0.ram_26_0.m0_s 
* net 359 = rbit_0_0.ram_26_0.m1_s 
* net 360 = rbit_0_0.ram_25_1.m0_s 
* net 361 = rbit_0_0.ram_25_1.m1_s 
* net 362 = rbit_0_0.ram_25_0.m0_s 
* net 363 = rbit_0_0.ram_25_0.m1_s 
* net 364 = rbit_0_0.ram_24_1.m0_s 
* net 365 = rbit_0_0.ram_24_1.m1_s 
* net 366 = rbit_0_0.ram_24_0.m0_s 
* net 367 = rbit_0_0.ram_24_0.m1_s 
* net 368 = rbit_0_0.ram_23_1.m0_s 
* net 369 = rbit_0_0.ram_23_1.m1_s 
* net 370 = rbit_0_0.ram_23_0.m0_s 
* net 371 = rbit_0_0.ram_23_0.m1_s 
* net 372 = rbit_0_0.ram_22_1.m0_s 
* net 373 = rbit_0_0.ram_22_1.m1_s 
* net 374 = rbit_0_0.ram_22_0.m0_s 
* net 375 = rbit_0_0.ram_22_0.m1_s 
* net 376 = rbit_0_0.ram_21_1.m0_s 
* net 377 = rbit_0_0.ram_21_1.m1_s 
* net 378 = rbit_0_0.ram_21_0.m0_s 
* net 379 = rbit_0_0.ram_21_0.m1_s 
* net 380 = rbit_0_0.ram_20_1.m0_s 
* net 381 = rbit_0_0.ram_20_1.m1_s 
* net 382 = rbit_0_0.ram_20_0.m0_s 
* net 383 = rbit_0_0.ram_20_0.m1_s 
* net 384 = rbit_0_0.ram_19_1.m0_s 
* net 385 = rbit_0_0.ram_19_1.m1_s 
* net 386 = rbit_0_0.ram_19_0.m0_s 
* net 387 = rbit_0_0.ram_19_0.m1_s 
* net 388 = rbit_0_0.ram_18_1.m0_s 
* net 389 = rbit_0_0.ram_18_1.m1_s 
* net 390 = rbit_0_0.ram_18_0.m0_s 
* net 391 = rbit_0_0.ram_18_0.m1_s 
* net 392 = rbit_0_0.ram_17_1.m0_s 
* net 393 = rbit_0_0.ram_17_1.m1_s 
* net 394 = rbit_0_0.ram_17_0.m0_s 
* net 395 = rbit_0_0.ram_17_0.m1_s 
* net 396 = rbit_0_0.ram_16_1.m0_s 
* net 397 = rbit_0_0.ram_16_1.m1_s 
* net 398 = rbit_0_0.ram_16_0.m0_s 
* net 399 = rbit_0_0.ram_16_0.m1_s 
* net 400 = rbit_0_0.ram_15_1.m0_s 
* net 401 = rbit_0_0.ram_15_1.m1_s 
* net 402 = rbit_0_0.ram_15_0.m0_s 
* net 403 = rbit_0_0.ram_15_0.m1_s 
* net 404 = rbit_0_0.ram_14_1.m0_s 
* net 405 = rbit_0_0.ram_14_1.m1_s 
* net 406 = rbit_0_0.ram_14_0.m0_s 
* net 407 = rbit_0_0.ram_14_0.m1_s 
* net 408 = rbit_0_0.ram_13_1.m0_s 
* net 409 = rbit_0_0.ram_13_1.m1_s 
* net 410 = rbit_0_0.ram_13_0.m0_s 
* net 411 = rbit_0_0.ram_13_0.m1_s 
* net 412 = rbit_0_0.ram_12_1.m0_s 
* net 413 = rbit_0_0.ram_12_1.m1_s 
* net 414 = rbit_0_0.ram_12_0.m0_s 
* net 415 = rbit_0_0.ram_12_0.m1_s 
* net 416 = rbit_0_0.ram_11_1.m0_s 
* net 417 = rbit_0_0.ram_11_1.m1_s 
* net 418 = rbit_0_0.ram_11_0.m0_s 
* net 419 = rbit_0_0.ram_11_0.m1_s 
* net 420 = rbit_0_0.ram_10_1.m0_s 
* net 421 = rbit_0_0.ram_10_1.m1_s 
* net 422 = rbit_0_0.ram_10_0.m0_s 
* net 423 = rbit_0_0.ram_10_0.m1_s 
* net 424 = rbit_0_0.ram_9_1.m0_s 
* net 425 = rbit_0_0.ram_9_1.m1_s 
* net 426 = rbit_0_0.ram_9_0.m0_s 
* net 427 = rbit_0_0.ram_9_0.m1_s 
* net 428 = rbit_0_0.ram_8_1.m0_s 
* net 429 = rbit_0_0.ram_8_1.m1_s 
* net 430 = rbit_0_0.ram_8_0.m0_s 
* net 431 = rbit_0_0.ram_8_0.m1_s 
* net 432 = rbit_0_0.ram_7_1.m0_s 
* net 433 = rbit_0_0.ram_7_1.m1_s 
* net 434 = rbit_0_0.ram_7_0.m0_s 
* net 435 = rbit_0_0.ram_7_0.m1_s 
* net 436 = rbit_0_0.ram_6_1.m0_s 
* net 437 = rbit_0_0.ram_6_1.m1_s 
* net 438 = rbit_0_0.ram_6_0.m0_s 
* net 439 = rbit_0_0.ram_6_0.m1_s 
* net 440 = rbit_0_0.ram_5_1.m0_s 
* net 441 = rbit_0_0.ram_5_1.m1_s 
* net 442 = rbit_0_0.ram_5_0.m0_s 
* net 443 = rbit_0_0.ram_5_0.m1_s 
* net 444 = rbit_0_0.ram_4_1.m0_s 
* net 445 = rbit_0_0.ram_4_1.m1_s 
* net 446 = rbit_0_0.ram_4_0.m0_s 
* net 447 = rbit_0_0.ram_4_0.m1_s 
* net 448 = rbit_0_0.ram_3_1.m0_s 
* net 449 = rbit_0_0.ram_3_1.m1_s 
* net 450 = rbit_0_0.ram_3_0.m0_s 
* net 451 = rbit_0_0.ram_3_0.m1_s 
* net 452 = rbit_0_0.ram_2_1.m0_s 
* net 453 = rbit_0_0.ram_2_1.m1_s 
* net 454 = rbit_0_0.ram_2_0.m0_s 
* net 455 = rbit_0_0.ram_2_0.m1_s 
* net 456 = rbit_0_0.ram_1_1.m0_s 
* net 457 = rbit_0_0.ram_1_1.m1_s 
* net 458 = rbit_0_0.ram_1_0.m0_s 
* net 459 = rbit_0_0.ram_1_0.m1_s 
* net 460 = rbit_0_0.ram_0_1.m0_s 
* net 461 = rbit_0_0.ram_0_1.m1_s 
* net 462 = rbit_0_0.ram_0_0.m0_s 
* net 463 = rbit_0_0.ram_0_0.m1_s 
* net 464 = mbk_sig88 
* net 465 = mbk_sig72 
* net 466 = mbk_sig105 
* net 467 = mbk_sig71 
* net 468 = mbk_sig119 
* net 469 = mbk_sig4 
* net 470 = mbk_sig2 
* net 471 = mbk_sig45 
* net 472 = mbk_sig65 
* net 473 = mbk_sig61 
* net 474 = mbk_sig57 
* net 475 = rbit_1_0.ram_63_1.m0_s 
* net 476 = rbit_1_0.ram_63_1.m1_s 
* net 477 = rbit_1_0.ram_63_0.m0_s 
* net 478 = rbit_1_0.ram_63_0.m1_s 
* net 479 = rbit_1_0.ram_62_1.m0_s 
* net 480 = rbit_1_0.ram_62_1.m1_s 
* net 481 = rbit_1_0.ram_62_0.m0_s 
* net 482 = rbit_1_0.ram_62_0.m1_s 
* net 483 = rbit_1_0.ram_61_1.m0_s 
* net 484 = rbit_1_0.ram_61_1.m1_s 
* net 485 = rbit_1_0.ram_61_0.m0_s 
* net 486 = rbit_1_0.ram_61_0.m1_s 
* net 487 = rbit_1_0.ram_60_1.m0_s 
* net 488 = rbit_1_0.ram_60_1.m1_s 
* net 489 = rbit_1_0.ram_60_0.m0_s 
* net 490 = rbit_1_0.ram_60_0.m1_s 
* net 491 = rbit_1_0.ram_59_1.m0_s 
* net 492 = rbit_1_0.ram_59_1.m1_s 
* net 493 = rbit_1_0.ram_59_0.m0_s 
* net 494 = rbit_1_0.ram_59_0.m1_s 
* net 495 = rbit_1_0.ram_58_1.m0_s 
* net 496 = rbit_1_0.ram_58_1.m1_s 
* net 497 = rbit_1_0.ram_58_0.m0_s 
* net 498 = rbit_1_0.ram_58_0.m1_s 
* net 499 = rbit_1_0.ram_57_1.m0_s 
* net 500 = rbit_1_0.ram_57_1.m1_s 
* net 501 = rbit_1_0.ram_57_0.m0_s 
* net 502 = rbit_1_0.ram_57_0.m1_s 
* net 503 = rbit_1_0.ram_56_1.m0_s 
* net 504 = rbit_1_0.ram_56_1.m1_s 
* net 505 = rbit_1_0.ram_56_0.m0_s 
* net 506 = rbit_1_0.ram_56_0.m1_s 
* net 507 = rbit_1_0.ram_55_1.m0_s 
* net 508 = rbit_1_0.ram_55_1.m1_s 
* net 509 = rbit_1_0.ram_55_0.m0_s 
* net 510 = rbit_1_0.ram_55_0.m1_s 
* net 511 = rbit_1_0.ram_54_1.m0_s 
* net 512 = rbit_1_0.ram_54_1.m1_s 
* net 513 = rbit_1_0.ram_54_0.m0_s 
* net 514 = rbit_1_0.ram_54_0.m1_s 
* net 515 = rbit_1_0.ram_53_1.m0_s 
* net 516 = rbit_1_0.ram_53_1.m1_s 
* net 517 = rbit_1_0.ram_53_0.m0_s 
* net 518 = rbit_1_0.ram_53_0.m1_s 
* net 519 = rbit_1_0.ram_52_1.m0_s 
* net 520 = rbit_1_0.ram_52_1.m1_s 
* net 521 = rbit_1_0.ram_52_0.m0_s 
* net 522 = rbit_1_0.ram_52_0.m1_s 
* net 523 = rbit_1_0.ram_51_1.m0_s 
* net 524 = rbit_1_0.ram_51_1.m1_s 
* net 525 = rbit_1_0.ram_51_0.m0_s 
* net 526 = rbit_1_0.ram_51_0.m1_s 
* net 527 = rbit_1_0.ram_50_1.m0_s 
* net 528 = rbit_1_0.ram_50_1.m1_s 
* net 529 = rbit_1_0.ram_50_0.m0_s 
* net 530 = rbit_1_0.ram_50_0.m1_s 
* net 531 = rbit_1_0.ram_49_1.m0_s 
* net 532 = rbit_1_0.ram_49_1.m1_s 
* net 533 = rbit_1_0.ram_49_0.m0_s 
* net 534 = rbit_1_0.ram_49_0.m1_s 
* net 535 = rbit_1_0.ram_48_1.m0_s 
* net 536 = rbit_1_0.ram_48_1.m1_s 
* net 537 = rbit_1_0.ram_48_0.m0_s 
* net 538 = rbit_1_0.ram_48_0.m1_s 
* net 539 = rbit_1_0.ram_47_1.m0_s 
* net 540 = rbit_1_0.ram_47_1.m1_s 
* net 541 = rbit_1_0.ram_47_0.m0_s 
* net 542 = rbit_1_0.ram_47_0.m1_s 
* net 543 = rbit_1_0.ram_46_1.m0_s 
* net 544 = rbit_1_0.ram_46_1.m1_s 
* net 545 = rbit_1_0.ram_46_0.m0_s 
* net 546 = rbit_1_0.ram_46_0.m1_s 
* net 547 = rbit_1_0.ram_45_1.m0_s 
* net 548 = rbit_1_0.ram_45_1.m1_s 
* net 549 = rbit_1_0.ram_45_0.m0_s 
* net 550 = rbit_1_0.ram_45_0.m1_s 
* net 551 = rbit_1_0.ram_44_1.m0_s 
* net 552 = rbit_1_0.ram_44_1.m1_s 
* net 553 = rbit_1_0.ram_44_0.m0_s 
* net 554 = rbit_1_0.ram_44_0.m1_s 
* net 555 = rbit_1_0.ram_43_1.m0_s 
* net 556 = rbit_1_0.ram_43_1.m1_s 
* net 557 = rbit_1_0.ram_43_0.m0_s 
* net 558 = rbit_1_0.ram_43_0.m1_s 
* net 559 = rbit_1_0.ram_42_1.m0_s 
* net 560 = rbit_1_0.ram_42_1.m1_s 
* net 561 = rbit_1_0.ram_42_0.m0_s 
* net 562 = rbit_1_0.ram_42_0.m1_s 
* net 563 = rbit_1_0.ram_41_1.m0_s 
* net 564 = rbit_1_0.ram_41_1.m1_s 
* net 565 = rbit_1_0.ram_41_0.m0_s 
* net 566 = rbit_1_0.ram_41_0.m1_s 
* net 567 = rbit_1_0.ram_40_1.m0_s 
* net 568 = rbit_1_0.ram_40_1.m1_s 
* net 569 = rbit_1_0.ram_40_0.m0_s 
* net 570 = rbit_1_0.ram_40_0.m1_s 
* net 571 = rbit_1_0.ram_39_1.m0_s 
* net 572 = rbit_1_0.ram_39_1.m1_s 
* net 573 = rbit_1_0.ram_39_0.m0_s 
* net 574 = rbit_1_0.ram_39_0.m1_s 
* net 575 = rbit_1_0.ram_38_1.m0_s 
* net 576 = rbit_1_0.ram_38_1.m1_s 
* net 577 = rbit_1_0.ram_38_0.m0_s 
* net 578 = rbit_1_0.ram_38_0.m1_s 
* net 579 = rbit_1_0.ram_37_1.m0_s 
* net 580 = rbit_1_0.ram_37_1.m1_s 
* net 581 = rbit_1_0.ram_37_0.m0_s 
* net 582 = rbit_1_0.ram_37_0.m1_s 
* net 583 = rbit_1_0.ram_36_1.m0_s 
* net 584 = rbit_1_0.ram_36_1.m1_s 
* net 585 = rbit_1_0.ram_36_0.m0_s 
* net 586 = rbit_1_0.ram_36_0.m1_s 
* net 587 = rbit_1_0.ram_35_1.m0_s 
* net 588 = rbit_1_0.ram_35_1.m1_s 
* net 589 = rbit_1_0.ram_35_0.m0_s 
* net 590 = rbit_1_0.ram_35_0.m1_s 
* net 591 = rbit_1_0.ram_34_1.m0_s 
* net 592 = rbit_1_0.ram_34_1.m1_s 
* net 593 = rbit_1_0.ram_34_0.m0_s 
* net 594 = rbit_1_0.ram_34_0.m1_s 
* net 595 = rbit_1_0.ram_33_1.m0_s 
* net 596 = rbit_1_0.ram_33_1.m1_s 
* net 597 = rbit_1_0.ram_33_0.m0_s 
* net 598 = rbit_1_0.ram_33_0.m1_s 
* net 599 = rbit_1_0.ram_32_1.m0_s 
* net 600 = rbit_1_0.ram_32_1.m1_s 
* net 601 = rbit_1_0.ram_32_0.m0_s 
* net 602 = rbit_1_0.ram_32_0.m1_s 
* net 603 = rbit_1_0.ram_31_1.m0_s 
* net 604 = rbit_1_0.ram_31_1.m1_s 
* net 605 = rbit_1_0.ram_31_0.m0_s 
* net 606 = rbit_1_0.ram_31_0.m1_s 
* net 607 = rbit_1_0.ram_30_1.m0_s 
* net 608 = rbit_1_0.ram_30_1.m1_s 
* net 609 = rbit_1_0.ram_30_0.m0_s 
* net 610 = rbit_1_0.ram_30_0.m1_s 
* net 611 = rbit_1_0.ram_29_1.m0_s 
* net 612 = rbit_1_0.ram_29_1.m1_s 
* net 613 = rbit_1_0.ram_29_0.m0_s 
* net 614 = rbit_1_0.ram_29_0.m1_s 
* net 615 = rbit_1_0.ram_28_1.m0_s 
* net 616 = rbit_1_0.ram_28_1.m1_s 
* net 617 = rbit_1_0.ram_28_0.m0_s 
* net 618 = rbit_1_0.ram_28_0.m1_s 
* net 619 = rbit_1_0.ram_27_1.m0_s 
* net 620 = rbit_1_0.ram_27_1.m1_s 
* net 621 = rbit_1_0.ram_27_0.m0_s 
* net 622 = rbit_1_0.ram_27_0.m1_s 
* net 623 = rbit_1_0.ram_26_1.m0_s 
* net 624 = rbit_1_0.ram_26_1.m1_s 
* net 625 = rbit_1_0.ram_26_0.m0_s 
* net 626 = rbit_1_0.ram_26_0.m1_s 
* net 627 = rbit_1_0.ram_25_1.m0_s 
* net 628 = rbit_1_0.ram_25_1.m1_s 
* net 629 = rbit_1_0.ram_25_0.m0_s 
* net 630 = rbit_1_0.ram_25_0.m1_s 
* net 631 = rbit_1_0.ram_24_1.m0_s 
* net 632 = rbit_1_0.ram_24_1.m1_s 
* net 633 = rbit_1_0.ram_24_0.m0_s 
* net 634 = rbit_1_0.ram_24_0.m1_s 
* net 635 = rbit_1_0.ram_23_1.m0_s 
* net 636 = rbit_1_0.ram_23_1.m1_s 
* net 637 = rbit_1_0.ram_23_0.m0_s 
* net 638 = rbit_1_0.ram_23_0.m1_s 
* net 639 = rbit_1_0.ram_22_1.m0_s 
* net 640 = rbit_1_0.ram_22_1.m1_s 
* net 641 = rbit_1_0.ram_22_0.m0_s 
* net 642 = rbit_1_0.ram_22_0.m1_s 
* net 643 = rbit_1_0.ram_21_1.m0_s 
* net 644 = rbit_1_0.ram_21_1.m1_s 
* net 645 = rbit_1_0.ram_21_0.m0_s 
* net 646 = rbit_1_0.ram_21_0.m1_s 
* net 647 = rbit_1_0.ram_20_1.m0_s 
* net 648 = rbit_1_0.ram_20_1.m1_s 
* net 649 = rbit_1_0.ram_20_0.m0_s 
* net 650 = rbit_1_0.ram_20_0.m1_s 
* net 651 = rbit_1_0.ram_19_1.m0_s 
* net 652 = rbit_1_0.ram_19_1.m1_s 
* net 653 = rbit_1_0.ram_19_0.m0_s 
* net 654 = rbit_1_0.ram_19_0.m1_s 
* net 655 = rbit_1_0.ram_18_1.m0_s 
* net 656 = rbit_1_0.ram_18_1.m1_s 
* net 657 = rbit_1_0.ram_18_0.m0_s 
* net 658 = rbit_1_0.ram_18_0.m1_s 
* net 659 = rbit_1_0.ram_17_1.m0_s 
* net 660 = rbit_1_0.ram_17_1.m1_s 
* net 661 = rbit_1_0.ram_17_0.m0_s 
* net 662 = rbit_1_0.ram_17_0.m1_s 
* net 663 = rbit_1_0.ram_16_1.m0_s 
* net 664 = rbit_1_0.ram_16_1.m1_s 
* net 665 = rbit_1_0.ram_16_0.m0_s 
* net 666 = rbit_1_0.ram_16_0.m1_s 
* net 667 = rbit_1_0.ram_15_1.m0_s 
* net 668 = rbit_1_0.ram_15_1.m1_s 
* net 669 = rbit_1_0.ram_15_0.m0_s 
* net 670 = rbit_1_0.ram_15_0.m1_s 
* net 671 = rbit_1_0.ram_14_1.m0_s 
* net 672 = rbit_1_0.ram_14_1.m1_s 
* net 673 = rbit_1_0.ram_14_0.m0_s 
* net 674 = rbit_1_0.ram_14_0.m1_s 
* net 675 = rbit_1_0.ram_13_1.m0_s 
* net 676 = rbit_1_0.ram_13_1.m1_s 
* net 677 = rbit_1_0.ram_13_0.m0_s 
* net 678 = rbit_1_0.ram_13_0.m1_s 
* net 679 = rbit_1_0.ram_12_1.m0_s 
* net 680 = rbit_1_0.ram_12_1.m1_s 
* net 681 = rbit_1_0.ram_12_0.m0_s 
* net 682 = rbit_1_0.ram_12_0.m1_s 
* net 683 = rbit_1_0.ram_11_1.m0_s 
* net 684 = rbit_1_0.ram_11_1.m1_s 
* net 685 = rbit_1_0.ram_11_0.m0_s 
* net 686 = rbit_1_0.ram_11_0.m1_s 
* net 687 = rbit_1_0.ram_10_1.m0_s 
* net 688 = rbit_1_0.ram_10_1.m1_s 
* net 689 = rbit_1_0.ram_10_0.m0_s 
* net 690 = rbit_1_0.ram_10_0.m1_s 
* net 691 = rbit_1_0.ram_9_1.m0_s 
* net 692 = rbit_1_0.ram_9_1.m1_s 
* net 693 = rbit_1_0.ram_9_0.m0_s 
* net 694 = rbit_1_0.ram_9_0.m1_s 
* net 695 = rbit_1_0.ram_8_1.m0_s 
* net 696 = rbit_1_0.ram_8_1.m1_s 
* net 697 = rbit_1_0.ram_8_0.m0_s 
* net 698 = rbit_1_0.ram_8_0.m1_s 
* net 699 = rbit_1_0.ram_7_1.m0_s 
* net 700 = rbit_1_0.ram_7_1.m1_s 
* net 701 = rbit_1_0.ram_7_0.m0_s 
* net 702 = rbit_1_0.ram_7_0.m1_s 
* net 703 = rbit_1_0.ram_6_1.m0_s 
* net 704 = rbit_1_0.ram_6_1.m1_s 
* net 705 = rbit_1_0.ram_6_0.m0_s 
* net 706 = rbit_1_0.ram_6_0.m1_s 
* net 707 = rbit_1_0.ram_5_1.m0_s 
* net 708 = rbit_1_0.ram_5_1.m1_s 
* net 709 = rbit_1_0.ram_5_0.m0_s 
* net 710 = rbit_1_0.ram_5_0.m1_s 
* net 711 = rbit_1_0.ram_4_1.m0_s 
* net 712 = rbit_1_0.ram_4_1.m1_s 
* net 713 = rbit_1_0.ram_4_0.m0_s 
* net 714 = rbit_1_0.ram_4_0.m1_s 
* net 715 = rbit_1_0.ram_3_1.m0_s 
* net 716 = rbit_1_0.ram_3_1.m1_s 
* net 717 = rbit_1_0.ram_3_0.m0_s 
* net 718 = rbit_1_0.ram_3_0.m1_s 
* net 719 = rbit_1_0.ram_2_1.m0_s 
* net 720 = rbit_1_0.ram_2_1.m1_s 
* net 721 = rbit_1_0.ram_2_0.m0_s 
* net 722 = rbit_1_0.ram_2_0.m1_s 
* net 723 = rbit_1_0.ram_1_1.m0_s 
* net 724 = rbit_1_0.ram_1_1.m1_s 
* net 725 = rbit_1_0.ram_1_0.m0_s 
* net 726 = rbit_1_0.ram_1_0.m1_s 
* net 727 = rbit_1_0.ram_0_1.m0_s 
* net 728 = rbit_1_0.ram_0_1.m1_s 
* net 729 = rbit_1_0.ram_0_0.m0_s 
* net 730 = rbit_1_0.ram_0_0.m1_s 
* net 731 = mbk_sig89 
* net 732 = mbk_sig73 
* net 733 = mbk_sig107 
* net 734 = mbk_sig74 
* net 735 = mbk_sig120 
* net 736 = mbk_sig11 
* net 737 = mbk_sig8 
* net 738 = mbk_sig46 
* net 739 = mbk_sig66 
* net 740 = mbk_sig62 
* net 741 = mbk_sig58 
* net 742 = mbk_sig1592 
* net 743 = mbk_sig1587 
* net 744 = mbk_sig1590 
* net 745 = mbk_sig1593 
* net 746 = mbk_sig1588 
* net 747 = mbk_sig1508 
* net 748 = mbk_sig1574 
* net 749 = mbk_sig1507 
* net 750 = decod.decd_15.wld[3] 
* net 751 = decod.decd_15.wld[2] 
* net 752 = decod.decd_15.wld[1] 
* net 753 = decod.decd_15.cd 
* net 754 = decod.decd_15.wld[0] 
* net 755 = decod.decg_15.wlg[2] 
* net 756 = mbk_sig1540 
* net 757 = decod.decg_15.wlg[1] 
* net 758 = mbk_sig1510 
* net 759 = decod.decg_15.wlg[0] 
* net 760 = mbk_sig1506 
* net 761 = decod.decg_15.wlg[3] 
* net 762 = mbk_sig1572 
* net 763 = mbk_sig1439 
* net 764 = mbk_sig1464 
* net 765 = mbk_sig1438 
* net 766 = decod.decd_14.wld[3] 
* net 767 = decod.decd_14.wld[2] 
* net 768 = decod.decd_14.wld[1] 
* net 769 = decod.decd_14.cd 
* net 770 = decod.decd_14.wld[0] 
* net 771 = decod.decg_14.wlg[2] 
* net 772 = mbk_sig1462 
* net 773 = decod.decg_14.wlg[1] 
* net 774 = mbk_sig1436 
* net 775 = decod.decg_14.wlg[0] 
* net 776 = mbk_sig1405 
* net 777 = decod.decg_14.wlg[3] 
* net 778 = mbk_sig1485 
* net 779 = mbk_sig1351 
* net 780 = mbk_sig1375 
* net 781 = mbk_sig1350 
* net 782 = decod.decd_13.wld[3] 
* net 783 = decod.decd_13.wld[2] 
* net 784 = decod.decd_13.wld[1] 
* net 785 = decod.decd_13.cd 
* net 786 = decod.decd_13.wld[0] 
* net 787 = decod.decg_13.wlg[2] 
* net 788 = mbk_sig1372 
* net 789 = decod.decg_13.wlg[1] 
* net 790 = mbk_sig1348 
* net 791 = decod.decg_13.wlg[0] 
* net 792 = mbk_sig1326 
* net 793 = decod.decg_13.wlg[3] 
* net 794 = mbk_sig1373 
* net 795 = mbk_sig1238 
* net 796 = mbk_sig1303 
* net 797 = mbk_sig1237 
* net 798 = decod.decd_12.wld[3] 
* net 799 = decod.decd_12.wld[2] 
* net 800 = decod.decd_12.wld[1] 
* net 801 = decod.decd_12.cd 
* net 802 = decod.decd_12.wld[0] 
* net 803 = decod.decg_12.wlg[2] 
* net 804 = mbk_sig1270 
* net 805 = decod.decg_12.wlg[1] 
* net 806 = mbk_sig1269 
* net 807 = decod.decg_12.wlg[0] 
* net 808 = mbk_sig1236 
* net 809 = decod.decg_12.wlg[3] 
* net 810 = mbk_sig1301 
* net 811 = mbk_sig1161 
* net 812 = mbk_sig1194 
* net 813 = mbk_sig1160 
* net 814 = decod.decd_11.wld[3] 
* net 815 = decod.decd_11.wld[2] 
* net 816 = decod.decd_11.wld[1] 
* net 817 = decod.decd_11.cd 
* net 818 = decod.decd_11.wld[0] 
* net 819 = decod.decg_11.wlg[2] 
* net 820 = mbk_sig1192 
* net 821 = decod.decg_11.wlg[1] 
* net 822 = mbk_sig1157 
* net 823 = decod.decg_11.wlg[0] 
* net 824 = mbk_sig1158 
* net 825 = decod.decg_11.wlg[3] 
* net 826 = mbk_sig1215 
* net 827 = mbk_sig1081 
* net 828 = mbk_sig1105 
* net 829 = mbk_sig1080 
* net 830 = decod.decd_10.wld[3] 
* net 831 = decod.decd_10.wld[2] 
* net 832 = decod.decd_10.wld[1] 
* net 833 = decod.decd_10.cd 
* net 834 = decod.decd_10.wld[0] 
* net 835 = decod.decg_10.wlg[2] 
* net 836 = mbk_sig1102 
* net 837 = decod.decg_10.wlg[1] 
* net 838 = mbk_sig1078 
* net 839 = decod.decg_10.wlg[0] 
* net 840 = mbk_sig1055 
* net 841 = decod.decg_10.wlg[3] 
* net 842 = mbk_sig1103 
* net 843 = mbk_sig992 
* net 844 = mbk_sig1024 
* net 845 = mbk_sig967 
* net 846 = decod.decd_9.wld[3] 
* net 847 = decod.decd_9.wld[2] 
* net 848 = decod.decd_9.wld[1] 
* net 849 = decod.decd_9.cd 
* net 850 = decod.decd_9.wld[0] 
* net 851 = decod.decg_9.wlg[2] 
* net 852 = mbk_sig990 
* net 853 = decod.decg_9.wlg[1] 
* net 854 = mbk_sig989 
* net 855 = decod.decg_9.wlg[0] 
* net 856 = mbk_sig966 
* net 857 = decod.decg_9.wlg[3] 
* net 858 = mbk_sig1022 
* net 859 = mbk_sig889 
* net 860 = mbk_sig923 
* net 861 = mbk_sig888 
* net 862 = decod.decd_8.wld[3] 
* net 863 = decod.decd_8.wld[2] 
* net 864 = decod.decd_8.wld[1] 
* net 865 = decod.decd_8.cd 
* net 866 = decod.decd_8.wld[0] 
* net 867 = decod.decg_8.wlg[2] 
* net 868 = mbk_sig921 
* net 869 = decod.decg_8.wlg[1] 
* net 870 = mbk_sig886 
* net 871 = decod.decg_8.wlg[0] 
* net 872 = mbk_sig884 
* net 873 = decod.decg_8.wlg[3] 
* net 874 = mbk_sig945 
* net 875 = mbk_sig811 
* net 876 = mbk_sig835 
* net 877 = mbk_sig810 
* net 878 = decod.decd_7.wld[3] 
* net 879 = decod.decd_7.wld[2] 
* net 880 = decod.decd_7.wld[1] 
* net 881 = decod.decd_7.cd 
* net 882 = decod.decd_7.wld[0] 
* net 883 = decod.decg_7.wlg[2] 
* net 884 = mbk_sig832 
* net 885 = decod.decg_7.wlg[1] 
* net 886 = mbk_sig808 
* net 887 = decod.decg_7.wlg[0] 
* net 888 = mbk_sig784 
* net 889 = decod.decg_7.wlg[3] 
* net 890 = mbk_sig833 
* net 891 = mbk_sig722 
* net 892 = mbk_sig754 
* net 893 = mbk_sig721 
* net 894 = decod.decd_6.wld[3] 
* net 895 = decod.decd_6.wld[2] 
* net 896 = decod.decd_6.wld[1] 
* net 897 = decod.decd_6.cd 
* net 898 = decod.decd_6.wld[0] 
* net 899 = decod.decg_6.wlg[2] 
* net 900 = mbk_sig719 
* net 901 = decod.decg_6.wlg[1] 
* net 902 = mbk_sig718 
* net 903 = decod.decg_6.wlg[0] 
* net 904 = mbk_sig696 
* net 905 = decod.decg_6.wlg[3] 
* net 906 = mbk_sig752 
* net 907 = mbk_sig608 
* net 908 = mbk_sig674 
* net 909 = mbk_sig607 
* net 910 = decod.decd_5.wld[3] 
* net 911 = decod.decd_5.wld[2] 
* net 912 = decod.decd_5.wld[1] 
* net 913 = decod.decd_5.cd 
* net 914 = decod.decd_5.wld[0] 
* net 915 = decod.decg_5.wlg[2] 
* net 916 = mbk_sig640 
* net 917 = decod.decg_5.wlg[1] 
* net 918 = mbk_sig610 
* net 919 = decod.decg_5.wlg[0] 
* net 920 = mbk_sig606 
* net 921 = decod.decg_5.wlg[3] 
* net 922 = mbk_sig672 
* net 923 = mbk_sig540 
* net 924 = mbk_sig564 
* net 925 = mbk_sig539 
* net 926 = decod.decd_4.wld[3] 
* net 927 = decod.decd_4.wld[2] 
* net 928 = decod.decd_4.wld[1] 
* net 929 = decod.decd_4.cd 
* net 930 = decod.decd_4.wld[0] 
* net 931 = decod.decg_4.wlg[2] 
* net 932 = mbk_sig562 
* net 933 = decod.decg_4.wlg[1] 
* net 934 = mbk_sig537 
* net 935 = decod.decg_4.wlg[0] 
* net 936 = mbk_sig505 
* net 937 = decod.decg_4.wlg[3] 
* net 938 = mbk_sig585 
* net 939 = mbk_sig452 
* net 940 = mbk_sig475 
* net 941 = mbk_sig451 
* net 942 = decod.decd_3.wld[3] 
* net 943 = decod.decd_3.wld[2] 
* net 944 = decod.decd_3.wld[1] 
* net 945 = decod.decd_3.cd 
* net 946 = decod.decd_3.wld[0] 
* net 947 = decod.decg_3.wlg[2] 
* net 948 = mbk_sig449 
* net 949 = decod.decg_3.wlg[1] 
* net 950 = mbk_sig448 
* net 951 = decod.decg_3.wlg[0] 
* net 952 = mbk_sig426 
* net 953 = decod.decg_3.wlg[3] 
* net 954 = mbk_sig473 
* net 955 = mbk_sig338 
* net 956 = mbk_sig403 
* net 957 = mbk_sig337 
* net 958 = decod.decd_2.wld[3] 
* net 959 = decod.decd_2.wld[2] 
* net 960 = decod.decd_2.wld[1] 
* net 961 = decod.decd_2.cd 
* net 962 = decod.decd_2.wld[0] 
* net 963 = decod.decg_2.wlg[2] 
* net 964 = mbk_sig370 
* net 965 = decod.decg_2.wlg[1] 
* net 966 = mbk_sig369 
* net 967 = decod.decg_2.wlg[0] 
* net 968 = mbk_sig336 
* net 969 = decod.decg_2.wlg[3] 
* net 970 = mbk_sig401 
* net 971 = mbk_sig269 
* net 972 = mbk_sig294 
* net 973 = mbk_sig268 
* net 974 = decod.decd_1.wld[3] 
* net 975 = decod.decd_1.wld[2] 
* net 976 = decod.decd_1.wld[1] 
* net 977 = decod.decd_1.cd 
* net 978 = decod.decd_1.wld[0] 
* net 979 = decod.decg_1.wlg[2] 
* net 980 = mbk_sig292 
* net 981 = decod.decg_1.wlg[1] 
* net 982 = mbk_sig266 
* net 983 = decod.decg_1.wlg[0] 
* net 984 = mbk_sig235 
* net 985 = decod.decg_1.wlg[3] 
* net 986 = mbk_sig315 
* net 987 = mbk_sig181 
* net 988 = mbk_sig205 
* net 989 = mbk_sig180 
* net 990 = decod.decd_0.wld[3] 
* net 991 = decod.decd_0.wld[2] 
* net 992 = decod.decd_0.wld[1] 
* net 993 = decod.decd_0.cd 
* net 994 = decod.decd_0.wld[0] 
* net 995 = decod.decg_0.wlg[2] 
* net 996 = mbk_sig202 
* net 997 = decod.decg_0.wlg[1] 
* net 998 = mbk_sig178 
* net 999 = decod.decg_0.wlg[0] 
* net 1000 = mbk_sig156 
* net 1001 = decod.decg_0.wlg[3] 
* net 1002 = mbk_sig203 
* net 1003 = mbk_sig130 
* net 1004 = mbk_sig131 
* net 1005 = mbk_sig117 
* net 1006 = decod.adr_1.adr_n[7] 
* net 1007 = mbk_sig122 
* net 1008 = mbk_sig109 
* net 1009 = mbk_sig116 
* net 1010 = mbk_sig118 
* net 1011 = mbk_sig110 
* net 1012 = mbk_sig108 
* net 1013 = mbk_sig111 
* net 1014 = mbk_sig102 
* net 1015 = mbk_sig101 
* net 1016 = mbk_sig103 
* net 1017 = mbk_sig75 
* net 1018 = mbk_sig80 
* net 1019 = decod.decd_0.cp[3] 
* net 1020 = mbk_sig93 
* net 1021 = mbk_sig94 
* net 1022 = decod.decd_0.cp[1] 
* net 1023 = decod.decd_0.cp[2] 
* net 1024 = mbk_sig76 
* net 1025 = mbk_sig78 
* net 1026 = decod.decd_0.cp[0] 
* net 1027 = mbk_sig70 
* net 1028 = mbk_sig69 
* net 1029 = mbk_sig55 
* net 1030 = mbk_sig49 
* net 1031 = mbk_sig51 
* net 1032 = mbk_sig5 
* net 1033 = mbk_sig47 
* net 1034 = mbk_sig50 
* net 1035 = mbk_sig43 
* net 1036 = mbk_sig33 
* net 1037 = mbk_sig40 
* net 1038 = mbk_sig6 
* net 1039 = mbk_sig42 
* net 1040 = decod.compg.cmk[0] 
* net 1041 = mbk_sig15 
* net 1042 = rbit_0_1.ram_63_1.m0_s 
* net 1043 = rbit_0_1.ram_63_1.m1_s 
* net 1044 = rbit_0_1.ram_63_0.m0_s 
* net 1045 = rbit_0_1.ram_63_0.m1_s 
* net 1046 = rbit_0_1.ram_62_1.m0_s 
* net 1047 = rbit_0_1.ram_62_1.m1_s 
* net 1048 = rbit_0_1.ram_62_0.m0_s 
* net 1049 = rbit_0_1.ram_62_0.m1_s 
* net 1050 = rbit_0_1.ram_61_1.m0_s 
* net 1051 = rbit_0_1.ram_61_1.m1_s 
* net 1052 = rbit_0_1.ram_61_0.m0_s 
* net 1053 = rbit_0_1.ram_61_0.m1_s 
* net 1054 = rbit_0_1.ram_60_1.m0_s 
* net 1055 = rbit_0_1.ram_60_1.m1_s 
* net 1056 = rbit_0_1.ram_60_0.m0_s 
* net 1057 = rbit_0_1.ram_60_0.m1_s 
* net 1058 = rbit_0_1.ram_59_1.m0_s 
* net 1059 = rbit_0_1.ram_59_1.m1_s 
* net 1060 = rbit_0_1.ram_59_0.m0_s 
* net 1061 = rbit_0_1.ram_59_0.m1_s 
* net 1062 = rbit_0_1.ram_58_1.m0_s 
* net 1063 = rbit_0_1.ram_58_1.m1_s 
* net 1064 = rbit_0_1.ram_58_0.m0_s 
* net 1065 = rbit_0_1.ram_58_0.m1_s 
* net 1066 = rbit_0_1.ram_57_1.m0_s 
* net 1067 = rbit_0_1.ram_57_1.m1_s 
* net 1068 = rbit_0_1.ram_57_0.m0_s 
* net 1069 = rbit_0_1.ram_57_0.m1_s 
* net 1070 = rbit_0_1.ram_56_1.m0_s 
* net 1071 = rbit_0_1.ram_56_1.m1_s 
* net 1072 = rbit_0_1.ram_56_0.m0_s 
* net 1073 = rbit_0_1.ram_56_0.m1_s 
* net 1074 = rbit_0_1.ram_55_1.m0_s 
* net 1075 = rbit_0_1.ram_55_1.m1_s 
* net 1076 = rbit_0_1.ram_55_0.m0_s 
* net 1077 = rbit_0_1.ram_55_0.m1_s 
* net 1078 = rbit_0_1.ram_54_1.m0_s 
* net 1079 = rbit_0_1.ram_54_1.m1_s 
* net 1080 = rbit_0_1.ram_54_0.m0_s 
* net 1081 = rbit_0_1.ram_54_0.m1_s 
* net 1082 = rbit_0_1.ram_53_1.m0_s 
* net 1083 = rbit_0_1.ram_53_1.m1_s 
* net 1084 = rbit_0_1.ram_53_0.m0_s 
* net 1085 = rbit_0_1.ram_53_0.m1_s 
* net 1086 = rbit_0_1.ram_52_1.m0_s 
* net 1087 = rbit_0_1.ram_52_1.m1_s 
* net 1088 = rbit_0_1.ram_52_0.m0_s 
* net 1089 = rbit_0_1.ram_52_0.m1_s 
* net 1090 = rbit_0_1.ram_51_1.m0_s 
* net 1091 = rbit_0_1.ram_51_1.m1_s 
* net 1092 = rbit_0_1.ram_51_0.m0_s 
* net 1093 = rbit_0_1.ram_51_0.m1_s 
* net 1094 = rbit_0_1.ram_50_1.m0_s 
* net 1095 = rbit_0_1.ram_50_1.m1_s 
* net 1096 = rbit_0_1.ram_50_0.m0_s 
* net 1097 = rbit_0_1.ram_50_0.m1_s 
* net 1098 = rbit_0_1.ram_49_1.m0_s 
* net 1099 = rbit_0_1.ram_49_1.m1_s 
* net 1100 = rbit_0_1.ram_49_0.m0_s 
* net 1101 = rbit_0_1.ram_49_0.m1_s 
* net 1102 = rbit_0_1.ram_48_1.m0_s 
* net 1103 = rbit_0_1.ram_48_1.m1_s 
* net 1104 = rbit_0_1.ram_48_0.m0_s 
* net 1105 = rbit_0_1.ram_48_0.m1_s 
* net 1106 = rbit_0_1.ram_47_1.m0_s 
* net 1107 = rbit_0_1.ram_47_1.m1_s 
* net 1108 = rbit_0_1.ram_47_0.m0_s 
* net 1109 = rbit_0_1.ram_47_0.m1_s 
* net 1110 = rbit_0_1.ram_46_1.m0_s 
* net 1111 = rbit_0_1.ram_46_1.m1_s 
* net 1112 = rbit_0_1.ram_46_0.m0_s 
* net 1113 = rbit_0_1.ram_46_0.m1_s 
* net 1114 = rbit_0_1.ram_45_1.m0_s 
* net 1115 = rbit_0_1.ram_45_1.m1_s 
* net 1116 = rbit_0_1.ram_45_0.m0_s 
* net 1117 = rbit_0_1.ram_45_0.m1_s 
* net 1118 = rbit_0_1.ram_44_1.m0_s 
* net 1119 = rbit_0_1.ram_44_1.m1_s 
* net 1120 = rbit_0_1.ram_44_0.m0_s 
* net 1121 = rbit_0_1.ram_44_0.m1_s 
* net 1122 = rbit_0_1.ram_43_1.m0_s 
* net 1123 = rbit_0_1.ram_43_1.m1_s 
* net 1124 = rbit_0_1.ram_43_0.m0_s 
* net 1125 = rbit_0_1.ram_43_0.m1_s 
* net 1126 = rbit_0_1.ram_42_1.m0_s 
* net 1127 = rbit_0_1.ram_42_1.m1_s 
* net 1128 = rbit_0_1.ram_42_0.m0_s 
* net 1129 = rbit_0_1.ram_42_0.m1_s 
* net 1130 = rbit_0_1.ram_41_1.m0_s 
* net 1131 = rbit_0_1.ram_41_1.m1_s 
* net 1132 = rbit_0_1.ram_41_0.m0_s 
* net 1133 = rbit_0_1.ram_41_0.m1_s 
* net 1134 = rbit_0_1.ram_40_1.m0_s 
* net 1135 = rbit_0_1.ram_40_1.m1_s 
* net 1136 = rbit_0_1.ram_40_0.m0_s 
* net 1137 = rbit_0_1.ram_40_0.m1_s 
* net 1138 = rbit_0_1.ram_39_1.m0_s 
* net 1139 = rbit_0_1.ram_39_1.m1_s 
* net 1140 = rbit_0_1.ram_39_0.m0_s 
* net 1141 = rbit_0_1.ram_39_0.m1_s 
* net 1142 = rbit_0_1.ram_38_1.m0_s 
* net 1143 = rbit_0_1.ram_38_1.m1_s 
* net 1144 = rbit_0_1.ram_38_0.m0_s 
* net 1145 = rbit_0_1.ram_38_0.m1_s 
* net 1146 = rbit_0_1.ram_37_1.m0_s 
* net 1147 = rbit_0_1.ram_37_1.m1_s 
* net 1148 = rbit_0_1.ram_37_0.m0_s 
* net 1149 = rbit_0_1.ram_37_0.m1_s 
* net 1150 = rbit_0_1.ram_36_1.m0_s 
* net 1151 = rbit_0_1.ram_36_1.m1_s 
* net 1152 = rbit_0_1.ram_36_0.m0_s 
* net 1153 = rbit_0_1.ram_36_0.m1_s 
* net 1154 = rbit_0_1.ram_35_1.m0_s 
* net 1155 = rbit_0_1.ram_35_1.m1_s 
* net 1156 = rbit_0_1.ram_35_0.m0_s 
* net 1157 = rbit_0_1.ram_35_0.m1_s 
* net 1158 = rbit_0_1.ram_34_1.m0_s 
* net 1159 = rbit_0_1.ram_34_1.m1_s 
* net 1160 = rbit_0_1.ram_34_0.m0_s 
* net 1161 = rbit_0_1.ram_34_0.m1_s 
* net 1162 = rbit_0_1.ram_33_1.m0_s 
* net 1163 = rbit_0_1.ram_33_1.m1_s 
* net 1164 = rbit_0_1.ram_33_0.m0_s 
* net 1165 = rbit_0_1.ram_33_0.m1_s 
* net 1166 = rbit_0_1.ram_32_1.m0_s 
* net 1167 = rbit_0_1.ram_32_1.m1_s 
* net 1168 = rbit_0_1.ram_32_0.m0_s 
* net 1169 = rbit_0_1.ram_32_0.m1_s 
* net 1170 = rbit_0_1.ram_31_1.m0_s 
* net 1171 = rbit_0_1.ram_31_1.m1_s 
* net 1172 = rbit_0_1.ram_31_0.m0_s 
* net 1173 = rbit_0_1.ram_31_0.m1_s 
* net 1174 = rbit_0_1.ram_30_1.m0_s 
* net 1175 = rbit_0_1.ram_30_1.m1_s 
* net 1176 = rbit_0_1.ram_30_0.m0_s 
* net 1177 = rbit_0_1.ram_30_0.m1_s 
* net 1178 = rbit_0_1.ram_29_1.m0_s 
* net 1179 = rbit_0_1.ram_29_1.m1_s 
* net 1180 = rbit_0_1.ram_29_0.m0_s 
* net 1181 = rbit_0_1.ram_29_0.m1_s 
* net 1182 = rbit_0_1.ram_28_1.m0_s 
* net 1183 = rbit_0_1.ram_28_1.m1_s 
* net 1184 = rbit_0_1.ram_28_0.m0_s 
* net 1185 = rbit_0_1.ram_28_0.m1_s 
* net 1186 = rbit_0_1.ram_27_1.m0_s 
* net 1187 = rbit_0_1.ram_27_1.m1_s 
* net 1188 = rbit_0_1.ram_27_0.m0_s 
* net 1189 = rbit_0_1.ram_27_0.m1_s 
* net 1190 = rbit_0_1.ram_26_1.m0_s 
* net 1191 = rbit_0_1.ram_26_1.m1_s 
* net 1192 = rbit_0_1.ram_26_0.m0_s 
* net 1193 = rbit_0_1.ram_26_0.m1_s 
* net 1194 = rbit_0_1.ram_25_1.m0_s 
* net 1195 = rbit_0_1.ram_25_1.m1_s 
* net 1196 = rbit_0_1.ram_25_0.m0_s 
* net 1197 = rbit_0_1.ram_25_0.m1_s 
* net 1198 = rbit_0_1.ram_24_1.m0_s 
* net 1199 = rbit_0_1.ram_24_1.m1_s 
* net 1200 = rbit_0_1.ram_24_0.m0_s 
* net 1201 = rbit_0_1.ram_24_0.m1_s 
* net 1202 = rbit_0_1.ram_23_1.m0_s 
* net 1203 = rbit_0_1.ram_23_1.m1_s 
* net 1204 = rbit_0_1.ram_23_0.m0_s 
* net 1205 = rbit_0_1.ram_23_0.m1_s 
* net 1206 = rbit_0_1.ram_22_1.m0_s 
* net 1207 = rbit_0_1.ram_22_1.m1_s 
* net 1208 = rbit_0_1.ram_22_0.m0_s 
* net 1209 = rbit_0_1.ram_22_0.m1_s 
* net 1210 = rbit_0_1.ram_21_1.m0_s 
* net 1211 = rbit_0_1.ram_21_1.m1_s 
* net 1212 = rbit_0_1.ram_21_0.m0_s 
* net 1213 = rbit_0_1.ram_21_0.m1_s 
* net 1214 = rbit_0_1.ram_20_1.m0_s 
* net 1215 = rbit_0_1.ram_20_1.m1_s 
* net 1216 = rbit_0_1.ram_20_0.m0_s 
* net 1217 = rbit_0_1.ram_20_0.m1_s 
* net 1218 = rbit_0_1.ram_19_1.m0_s 
* net 1219 = rbit_0_1.ram_19_1.m1_s 
* net 1220 = rbit_0_1.ram_19_0.m0_s 
* net 1221 = rbit_0_1.ram_19_0.m1_s 
* net 1222 = rbit_0_1.ram_18_1.m0_s 
* net 1223 = rbit_0_1.ram_18_1.m1_s 
* net 1224 = rbit_0_1.ram_18_0.m0_s 
* net 1225 = rbit_0_1.ram_18_0.m1_s 
* net 1226 = rbit_0_1.ram_17_1.m0_s 
* net 1227 = rbit_0_1.ram_17_1.m1_s 
* net 1228 = rbit_0_1.ram_17_0.m0_s 
* net 1229 = rbit_0_1.ram_17_0.m1_s 
* net 1230 = rbit_0_1.ram_16_1.m0_s 
* net 1231 = rbit_0_1.ram_16_1.m1_s 
* net 1232 = rbit_0_1.ram_16_0.m0_s 
* net 1233 = rbit_0_1.ram_16_0.m1_s 
* net 1234 = rbit_0_1.ram_15_1.m0_s 
* net 1235 = rbit_0_1.ram_15_1.m1_s 
* net 1236 = rbit_0_1.ram_15_0.m0_s 
* net 1237 = rbit_0_1.ram_15_0.m1_s 
* net 1238 = rbit_0_1.ram_14_1.m0_s 
* net 1239 = rbit_0_1.ram_14_1.m1_s 
* net 1240 = rbit_0_1.ram_14_0.m0_s 
* net 1241 = rbit_0_1.ram_14_0.m1_s 
* net 1242 = rbit_0_1.ram_13_1.m0_s 
* net 1243 = rbit_0_1.ram_13_1.m1_s 
* net 1244 = rbit_0_1.ram_13_0.m0_s 
* net 1245 = rbit_0_1.ram_13_0.m1_s 
* net 1246 = rbit_0_1.ram_12_1.m0_s 
* net 1247 = rbit_0_1.ram_12_1.m1_s 
* net 1248 = rbit_0_1.ram_12_0.m0_s 
* net 1249 = rbit_0_1.ram_12_0.m1_s 
* net 1250 = rbit_0_1.ram_11_1.m0_s 
* net 1251 = rbit_0_1.ram_11_1.m1_s 
* net 1252 = rbit_0_1.ram_11_0.m0_s 
* net 1253 = rbit_0_1.ram_11_0.m1_s 
* net 1254 = rbit_0_1.ram_10_1.m0_s 
* net 1255 = rbit_0_1.ram_10_1.m1_s 
* net 1256 = rbit_0_1.ram_10_0.m0_s 
* net 1257 = rbit_0_1.ram_10_0.m1_s 
* net 1258 = rbit_0_1.ram_9_1.m0_s 
* net 1259 = rbit_0_1.ram_9_1.m1_s 
* net 1260 = rbit_0_1.ram_9_0.m0_s 
* net 1261 = rbit_0_1.ram_9_0.m1_s 
* net 1262 = rbit_0_1.ram_8_1.m0_s 
* net 1263 = rbit_0_1.ram_8_1.m1_s 
* net 1264 = rbit_0_1.ram_8_0.m0_s 
* net 1265 = rbit_0_1.ram_8_0.m1_s 
* net 1266 = rbit_0_1.ram_7_1.m0_s 
* net 1267 = rbit_0_1.ram_7_1.m1_s 
* net 1268 = rbit_0_1.ram_7_0.m0_s 
* net 1269 = rbit_0_1.ram_7_0.m1_s 
* net 1270 = rbit_0_1.ram_6_1.m0_s 
* net 1271 = rbit_0_1.ram_6_1.m1_s 
* net 1272 = rbit_0_1.ram_6_0.m0_s 
* net 1273 = rbit_0_1.ram_6_0.m1_s 
* net 1274 = rbit_0_1.ram_5_1.m0_s 
* net 1275 = rbit_0_1.ram_5_1.m1_s 
* net 1276 = rbit_0_1.ram_5_0.m0_s 
* net 1277 = rbit_0_1.ram_5_0.m1_s 
* net 1278 = rbit_0_1.ram_4_1.m0_s 
* net 1279 = rbit_0_1.ram_4_1.m1_s 
* net 1280 = rbit_0_1.ram_4_0.m0_s 
* net 1281 = rbit_0_1.ram_4_0.m1_s 
* net 1282 = rbit_0_1.ram_3_1.m0_s 
* net 1283 = rbit_0_1.ram_3_1.m1_s 
* net 1284 = rbit_0_1.ram_3_0.m0_s 
* net 1285 = rbit_0_1.ram_3_0.m1_s 
* net 1286 = rbit_0_1.ram_2_1.m0_s 
* net 1287 = rbit_0_1.ram_2_1.m1_s 
* net 1288 = rbit_0_1.ram_2_0.m0_s 
* net 1289 = rbit_0_1.ram_2_0.m1_s 
* net 1290 = rbit_0_1.ram_1_1.m0_s 
* net 1291 = rbit_0_1.ram_1_1.m1_s 
* net 1292 = rbit_0_1.ram_1_0.m0_s 
* net 1293 = rbit_0_1.ram_1_0.m1_s 
* net 1294 = rbit_0_1.ram_0_1.m0_s 
* net 1295 = rbit_0_1.ram_0_1.m1_s 
* net 1296 = rbit_0_1.ram_0_0.m0_s 
* net 1297 = rbit_0_1.ram_0_0.m1_s 
* net 1298 = mbk_sig98 
* net 1299 = mbk_sig84 
* net 1300 = mbk_sig113 
* net 1301 = mbk_sig83 
* net 1302 = mbk_sig123 
* net 1303 = mbk_sig29 
* net 1304 = mbk_sig32 
* net 1305 = mbk_sig53 
* net 1306 = mbk_sig67 
* net 1307 = mbk_sig63 
* net 1308 = mbk_sig59 
* net 1309 = rbit_1_1.ram_63_1.m0_s 
* net 1310 = rbit_1_1.ram_63_1.m1_s 
* net 1311 = rbit_1_1.ram_63_0.m0_s 
* net 1312 = rbit_1_1.ram_63_0.m1_s 
* net 1313 = rbit_1_1.ram_62_1.m0_s 
* net 1314 = rbit_1_1.ram_62_1.m1_s 
* net 1315 = rbit_1_1.ram_62_0.m0_s 
* net 1316 = rbit_1_1.ram_62_0.m1_s 
* net 1317 = rbit_1_1.ram_61_1.m0_s 
* net 1318 = rbit_1_1.ram_61_1.m1_s 
* net 1319 = rbit_1_1.ram_61_0.m0_s 
* net 1320 = rbit_1_1.ram_61_0.m1_s 
* net 1321 = rbit_1_1.ram_60_1.m0_s 
* net 1322 = rbit_1_1.ram_60_1.m1_s 
* net 1323 = rbit_1_1.ram_60_0.m0_s 
* net 1324 = rbit_1_1.ram_60_0.m1_s 
* net 1325 = rbit_1_1.ram_59_1.m0_s 
* net 1326 = rbit_1_1.ram_59_1.m1_s 
* net 1327 = rbit_1_1.ram_59_0.m0_s 
* net 1328 = rbit_1_1.ram_59_0.m1_s 
* net 1329 = rbit_1_1.ram_58_1.m0_s 
* net 1330 = rbit_1_1.ram_58_1.m1_s 
* net 1331 = rbit_1_1.ram_58_0.m0_s 
* net 1332 = rbit_1_1.ram_58_0.m1_s 
* net 1333 = rbit_1_1.ram_57_1.m0_s 
* net 1334 = rbit_1_1.ram_57_1.m1_s 
* net 1335 = rbit_1_1.ram_57_0.m0_s 
* net 1336 = rbit_1_1.ram_57_0.m1_s 
* net 1337 = rbit_1_1.ram_56_1.m0_s 
* net 1338 = rbit_1_1.ram_56_1.m1_s 
* net 1339 = rbit_1_1.ram_56_0.m0_s 
* net 1340 = rbit_1_1.ram_56_0.m1_s 
* net 1341 = rbit_1_1.ram_55_1.m0_s 
* net 1342 = rbit_1_1.ram_55_1.m1_s 
* net 1343 = rbit_1_1.ram_55_0.m0_s 
* net 1344 = rbit_1_1.ram_55_0.m1_s 
* net 1345 = rbit_1_1.ram_54_1.m0_s 
* net 1346 = rbit_1_1.ram_54_1.m1_s 
* net 1347 = rbit_1_1.ram_54_0.m0_s 
* net 1348 = rbit_1_1.ram_54_0.m1_s 
* net 1349 = rbit_1_1.ram_53_1.m0_s 
* net 1350 = rbit_1_1.ram_53_1.m1_s 
* net 1351 = rbit_1_1.ram_53_0.m0_s 
* net 1352 = rbit_1_1.ram_53_0.m1_s 
* net 1353 = rbit_1_1.ram_52_1.m0_s 
* net 1354 = rbit_1_1.ram_52_1.m1_s 
* net 1355 = rbit_1_1.ram_52_0.m0_s 
* net 1356 = rbit_1_1.ram_52_0.m1_s 
* net 1357 = rbit_1_1.ram_51_1.m0_s 
* net 1358 = rbit_1_1.ram_51_1.m1_s 
* net 1359 = rbit_1_1.ram_51_0.m0_s 
* net 1360 = rbit_1_1.ram_51_0.m1_s 
* net 1361 = rbit_1_1.ram_50_1.m0_s 
* net 1362 = rbit_1_1.ram_50_1.m1_s 
* net 1363 = rbit_1_1.ram_50_0.m0_s 
* net 1364 = rbit_1_1.ram_50_0.m1_s 
* net 1365 = rbit_1_1.ram_49_1.m0_s 
* net 1366 = rbit_1_1.ram_49_1.m1_s 
* net 1367 = rbit_1_1.ram_49_0.m0_s 
* net 1368 = rbit_1_1.ram_49_0.m1_s 
* net 1369 = rbit_1_1.ram_48_1.m0_s 
* net 1370 = rbit_1_1.ram_48_1.m1_s 
* net 1371 = rbit_1_1.ram_48_0.m0_s 
* net 1372 = rbit_1_1.ram_48_0.m1_s 
* net 1373 = rbit_1_1.ram_47_1.m0_s 
* net 1374 = rbit_1_1.ram_47_1.m1_s 
* net 1375 = rbit_1_1.ram_47_0.m0_s 
* net 1376 = rbit_1_1.ram_47_0.m1_s 
* net 1377 = rbit_1_1.ram_46_1.m0_s 
* net 1378 = rbit_1_1.ram_46_1.m1_s 
* net 1379 = rbit_1_1.ram_46_0.m0_s 
* net 1380 = rbit_1_1.ram_46_0.m1_s 
* net 1381 = rbit_1_1.ram_45_1.m0_s 
* net 1382 = rbit_1_1.ram_45_1.m1_s 
* net 1383 = rbit_1_1.ram_45_0.m0_s 
* net 1384 = rbit_1_1.ram_45_0.m1_s 
* net 1385 = rbit_1_1.ram_44_1.m0_s 
* net 1386 = rbit_1_1.ram_44_1.m1_s 
* net 1387 = rbit_1_1.ram_44_0.m0_s 
* net 1388 = rbit_1_1.ram_44_0.m1_s 
* net 1389 = rbit_1_1.ram_43_1.m0_s 
* net 1390 = rbit_1_1.ram_43_1.m1_s 
* net 1391 = rbit_1_1.ram_43_0.m0_s 
* net 1392 = rbit_1_1.ram_43_0.m1_s 
* net 1393 = rbit_1_1.ram_42_1.m0_s 
* net 1394 = rbit_1_1.ram_42_1.m1_s 
* net 1395 = rbit_1_1.ram_42_0.m0_s 
* net 1396 = rbit_1_1.ram_42_0.m1_s 
* net 1397 = rbit_1_1.ram_41_1.m0_s 
* net 1398 = rbit_1_1.ram_41_1.m1_s 
* net 1399 = rbit_1_1.ram_41_0.m0_s 
* net 1400 = rbit_1_1.ram_41_0.m1_s 
* net 1401 = rbit_1_1.ram_40_1.m0_s 
* net 1402 = rbit_1_1.ram_40_1.m1_s 
* net 1403 = rbit_1_1.ram_40_0.m0_s 
* net 1404 = rbit_1_1.ram_40_0.m1_s 
* net 1405 = rbit_1_1.ram_39_1.m0_s 
* net 1406 = rbit_1_1.ram_39_1.m1_s 
* net 1407 = rbit_1_1.ram_39_0.m0_s 
* net 1408 = rbit_1_1.ram_39_0.m1_s 
* net 1409 = rbit_1_1.ram_38_1.m0_s 
* net 1410 = rbit_1_1.ram_38_1.m1_s 
* net 1411 = rbit_1_1.ram_38_0.m0_s 
* net 1412 = rbit_1_1.ram_38_0.m1_s 
* net 1413 = rbit_1_1.ram_37_1.m0_s 
* net 1414 = rbit_1_1.ram_37_1.m1_s 
* net 1415 = rbit_1_1.ram_37_0.m0_s 
* net 1416 = rbit_1_1.ram_37_0.m1_s 
* net 1417 = rbit_1_1.ram_36_1.m0_s 
* net 1418 = rbit_1_1.ram_36_1.m1_s 
* net 1419 = rbit_1_1.ram_36_0.m0_s 
* net 1420 = rbit_1_1.ram_36_0.m1_s 
* net 1421 = rbit_1_1.ram_35_1.m0_s 
* net 1422 = rbit_1_1.ram_35_1.m1_s 
* net 1423 = rbit_1_1.ram_35_0.m0_s 
* net 1424 = rbit_1_1.ram_35_0.m1_s 
* net 1425 = rbit_1_1.ram_34_1.m0_s 
* net 1426 = rbit_1_1.ram_34_1.m1_s 
* net 1427 = rbit_1_1.ram_34_0.m0_s 
* net 1428 = rbit_1_1.ram_34_0.m1_s 
* net 1429 = rbit_1_1.ram_33_1.m0_s 
* net 1430 = rbit_1_1.ram_33_1.m1_s 
* net 1431 = rbit_1_1.ram_33_0.m0_s 
* net 1432 = rbit_1_1.ram_33_0.m1_s 
* net 1433 = rbit_1_1.ram_32_1.m0_s 
* net 1434 = rbit_1_1.ram_32_1.m1_s 
* net 1435 = rbit_1_1.ram_32_0.m0_s 
* net 1436 = rbit_1_1.ram_32_0.m1_s 
* net 1437 = rbit_1_1.ram_31_1.m0_s 
* net 1438 = rbit_1_1.ram_31_1.m1_s 
* net 1439 = rbit_1_1.ram_31_0.m0_s 
* net 1440 = rbit_1_1.ram_31_0.m1_s 
* net 1441 = rbit_1_1.ram_30_1.m0_s 
* net 1442 = rbit_1_1.ram_30_1.m1_s 
* net 1443 = rbit_1_1.ram_30_0.m0_s 
* net 1444 = rbit_1_1.ram_30_0.m1_s 
* net 1445 = rbit_1_1.ram_29_1.m0_s 
* net 1446 = rbit_1_1.ram_29_1.m1_s 
* net 1447 = rbit_1_1.ram_29_0.m0_s 
* net 1448 = rbit_1_1.ram_29_0.m1_s 
* net 1449 = rbit_1_1.ram_28_1.m0_s 
* net 1450 = rbit_1_1.ram_28_1.m1_s 
* net 1451 = rbit_1_1.ram_28_0.m0_s 
* net 1452 = rbit_1_1.ram_28_0.m1_s 
* net 1453 = rbit_1_1.ram_27_1.m0_s 
* net 1454 = rbit_1_1.ram_27_1.m1_s 
* net 1455 = rbit_1_1.ram_27_0.m0_s 
* net 1456 = rbit_1_1.ram_27_0.m1_s 
* net 1457 = rbit_1_1.ram_26_1.m0_s 
* net 1458 = rbit_1_1.ram_26_1.m1_s 
* net 1459 = rbit_1_1.ram_26_0.m0_s 
* net 1460 = rbit_1_1.ram_26_0.m1_s 
* net 1461 = rbit_1_1.ram_25_1.m0_s 
* net 1462 = rbit_1_1.ram_25_1.m1_s 
* net 1463 = rbit_1_1.ram_25_0.m0_s 
* net 1464 = rbit_1_1.ram_25_0.m1_s 
* net 1465 = rbit_1_1.ram_24_1.m0_s 
* net 1466 = rbit_1_1.ram_24_1.m1_s 
* net 1467 = rbit_1_1.ram_24_0.m0_s 
* net 1468 = rbit_1_1.ram_24_0.m1_s 
* net 1469 = rbit_1_1.ram_23_1.m0_s 
* net 1470 = rbit_1_1.ram_23_1.m1_s 
* net 1471 = rbit_1_1.ram_23_0.m0_s 
* net 1472 = rbit_1_1.ram_23_0.m1_s 
* net 1473 = rbit_1_1.ram_22_1.m0_s 
* net 1474 = rbit_1_1.ram_22_1.m1_s 
* net 1475 = rbit_1_1.ram_22_0.m0_s 
* net 1476 = rbit_1_1.ram_22_0.m1_s 
* net 1477 = rbit_1_1.ram_21_1.m0_s 
* net 1478 = rbit_1_1.ram_21_1.m1_s 
* net 1479 = rbit_1_1.ram_21_0.m0_s 
* net 1480 = rbit_1_1.ram_21_0.m1_s 
* net 1481 = rbit_1_1.ram_20_1.m0_s 
* net 1482 = rbit_1_1.ram_20_1.m1_s 
* net 1483 = rbit_1_1.ram_20_0.m0_s 
* net 1484 = rbit_1_1.ram_20_0.m1_s 
* net 1485 = rbit_1_1.ram_19_1.m0_s 
* net 1486 = rbit_1_1.ram_19_1.m1_s 
* net 1487 = rbit_1_1.ram_19_0.m0_s 
* net 1488 = rbit_1_1.ram_19_0.m1_s 
* net 1489 = rbit_1_1.ram_18_1.m0_s 
* net 1490 = rbit_1_1.ram_18_1.m1_s 
* net 1491 = rbit_1_1.ram_18_0.m0_s 
* net 1492 = rbit_1_1.ram_18_0.m1_s 
* net 1493 = rbit_1_1.ram_17_1.m0_s 
* net 1494 = rbit_1_1.ram_17_1.m1_s 
* net 1495 = rbit_1_1.ram_17_0.m0_s 
* net 1496 = rbit_1_1.ram_17_0.m1_s 
* net 1497 = rbit_1_1.ram_16_1.m0_s 
* net 1498 = rbit_1_1.ram_16_1.m1_s 
* net 1499 = rbit_1_1.ram_16_0.m0_s 
* net 1500 = rbit_1_1.ram_16_0.m1_s 
* net 1501 = rbit_1_1.ram_15_1.m0_s 
* net 1502 = rbit_1_1.ram_15_1.m1_s 
* net 1503 = rbit_1_1.ram_15_0.m0_s 
* net 1504 = rbit_1_1.ram_15_0.m1_s 
* net 1505 = rbit_1_1.ram_14_1.m0_s 
* net 1506 = rbit_1_1.ram_14_1.m1_s 
* net 1507 = rbit_1_1.ram_14_0.m0_s 
* net 1508 = rbit_1_1.ram_14_0.m1_s 
* net 1509 = rbit_1_1.ram_13_1.m0_s 
* net 1510 = rbit_1_1.ram_13_1.m1_s 
* net 1511 = rbit_1_1.ram_13_0.m0_s 
* net 1512 = rbit_1_1.ram_13_0.m1_s 
* net 1513 = rbit_1_1.ram_12_1.m0_s 
* net 1514 = rbit_1_1.ram_12_1.m1_s 
* net 1515 = rbit_1_1.ram_12_0.m0_s 
* net 1516 = rbit_1_1.ram_12_0.m1_s 
* net 1517 = rbit_1_1.ram_11_1.m0_s 
* net 1518 = rbit_1_1.ram_11_1.m1_s 
* net 1519 = rbit_1_1.ram_11_0.m0_s 
* net 1520 = rbit_1_1.ram_11_0.m1_s 
* net 1521 = rbit_1_1.ram_10_1.m0_s 
* net 1522 = rbit_1_1.ram_10_1.m1_s 
* net 1523 = rbit_1_1.ram_10_0.m0_s 
* net 1524 = rbit_1_1.ram_10_0.m1_s 
* net 1525 = rbit_1_1.ram_9_1.m0_s 
* net 1526 = rbit_1_1.ram_9_1.m1_s 
* net 1527 = rbit_1_1.ram_9_0.m0_s 
* net 1528 = rbit_1_1.ram_9_0.m1_s 
* net 1529 = rbit_1_1.ram_8_1.m0_s 
* net 1530 = rbit_1_1.ram_8_1.m1_s 
* net 1531 = rbit_1_1.ram_8_0.m0_s 
* net 1532 = rbit_1_1.ram_8_0.m1_s 
* net 1533 = rbit_1_1.ram_7_1.m0_s 
* net 1534 = rbit_1_1.ram_7_1.m1_s 
* net 1535 = rbit_1_1.ram_7_0.m0_s 
* net 1536 = rbit_1_1.ram_7_0.m1_s 
* net 1537 = rbit_1_1.ram_6_1.m0_s 
* net 1538 = rbit_1_1.ram_6_1.m1_s 
* net 1539 = rbit_1_1.ram_6_0.m0_s 
* net 1540 = rbit_1_1.ram_6_0.m1_s 
* net 1541 = rbit_1_1.ram_5_1.m0_s 
* net 1542 = rbit_1_1.ram_5_1.m1_s 
* net 1543 = rbit_1_1.ram_5_0.m0_s 
* net 1544 = rbit_1_1.ram_5_0.m1_s 
* net 1545 = rbit_1_1.ram_4_1.m0_s 
* net 1546 = rbit_1_1.ram_4_1.m1_s 
* net 1547 = rbit_1_1.ram_4_0.m0_s 
* net 1548 = rbit_1_1.ram_4_0.m1_s 
* net 1549 = rbit_1_1.ram_3_1.m0_s 
* net 1550 = rbit_1_1.ram_3_1.m1_s 
* net 1551 = rbit_1_1.ram_3_0.m0_s 
* net 1552 = rbit_1_1.ram_3_0.m1_s 
* net 1553 = rbit_1_1.ram_2_1.m0_s 
* net 1554 = rbit_1_1.ram_2_1.m1_s 
* net 1555 = rbit_1_1.ram_2_0.m0_s 
* net 1556 = rbit_1_1.ram_2_0.m1_s 
* net 1557 = rbit_1_1.ram_1_1.m0_s 
* net 1558 = rbit_1_1.ram_1_1.m1_s 
* net 1559 = rbit_1_1.ram_1_0.m0_s 
* net 1560 = rbit_1_1.ram_1_0.m1_s 
* net 1561 = rbit_1_1.ram_0_1.m0_s 
* net 1562 = rbit_1_1.ram_0_1.m1_s 
* net 1563 = rbit_1_1.ram_0_0.m0_s 
* net 1564 = rbit_1_1.ram_0_0.m1_s 
* net 1565 = mbk_sig100 
* net 1566 = mbk_sig86 
* net 1567 = mbk_sig115 
* net 1568 = mbk_sig85 
* net 1569 = mbk_sig124 
* net 1570 = mbk_sig38 
* net 1571 = mbk_sig36 
* net 1572 = mbk_sig54 
* net 1573 = mbk_sig56 
* net 1574 = mbk_sig68 
* net 1575 = mbk_sig64 
* net 1576 = mbk_sig28 
* net 1577 = mbk_sig60 
* net 1578 = write 
* net 1579 = vss 
* net 1580 = vdd 
* net 1581 = en 
* net 1582 = dout[3] 
* net 1583 = dout[2] 
* net 1584 = dout[1] 
* net 1585 = dout[0] 
* net 1586 = ck 
* net 1587 = adr[6] 
* net 1588 = adr[5] 
* net 1589 = adr[4] 
* net 1590 = adr[3] 
* net 1591 = adr[2] 
* net 1592 = adr[1] 
* net 1593 = adr[0] 
Mtr_00001 4 743 2 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00002 4 743 1580 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00003 2 743 1580 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00004 3 743 1 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00005 1580 743 3 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00006 1580 743 1 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00007 1579 209 208 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00008 209 208 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00009 4 761 208 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00010 2 761 209 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00011 1579 211 210 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00012 211 210 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00013 3 761 210 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00014 1 761 211 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00015 1579 213 212 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00016 213 212 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00017 4 755 212 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00018 2 755 213 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00019 1579 215 214 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00020 215 214 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00021 3 755 214 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00022 1 755 215 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00023 1579 217 216 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00024 217 216 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00025 4 757 216 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00026 2 757 217 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00027 1579 219 218 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00028 219 218 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00029 3 757 218 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00030 1 757 219 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00031 1579 221 220 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00032 221 220 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00033 4 759 220 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00034 2 759 221 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00035 1579 223 222 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00036 223 222 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00037 3 759 222 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00038 1 759 223 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00039 1579 225 224 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00040 225 224 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00041 4 777 224 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00042 2 777 225 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00043 1579 227 226 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00044 227 226 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00045 3 777 226 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00046 1 777 227 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00047 1579 229 228 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00048 229 228 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00049 4 771 228 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00050 2 771 229 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00051 1579 231 230 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00052 231 230 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00053 3 771 230 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00054 1 771 231 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00055 1579 233 232 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00056 233 232 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00057 4 773 232 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00058 2 773 233 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00059 1579 235 234 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00060 235 234 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00061 3 773 234 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00062 1 773 235 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00063 1579 237 236 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00064 237 236 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00065 4 775 236 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00066 2 775 237 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00067 1579 239 238 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00068 239 238 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00069 3 775 238 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00070 1 775 239 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00071 1579 241 240 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00072 241 240 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00073 4 793 240 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00074 2 793 241 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00075 1579 243 242 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00076 243 242 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00077 3 793 242 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00078 1 793 243 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00079 1579 245 244 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00080 245 244 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00081 4 787 244 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00082 2 787 245 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00083 1579 247 246 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00084 247 246 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00085 3 787 246 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00086 1 787 247 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00087 1579 249 248 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00088 249 248 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00089 4 789 248 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00090 2 789 249 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00091 1579 251 250 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00092 251 250 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00093 3 789 250 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00094 1 789 251 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00095 1579 253 252 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00096 253 252 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00097 4 791 252 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00098 2 791 253 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00099 1579 255 254 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00100 255 254 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00101 3 791 254 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00102 1 791 255 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00103 1579 257 256 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00104 257 256 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00105 4 809 256 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00106 2 809 257 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00107 1579 259 258 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00108 259 258 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00109 3 809 258 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00110 1 809 259 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00111 1579 261 260 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00112 261 260 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00113 4 803 260 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00114 2 803 261 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00115 1579 263 262 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00116 263 262 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00117 3 803 262 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00118 1 803 263 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00119 1579 265 264 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00120 265 264 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00121 4 805 264 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00122 2 805 265 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00123 1579 267 266 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00124 267 266 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00125 3 805 266 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00126 1 805 267 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00127 1579 269 268 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00128 269 268 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00129 4 807 268 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00130 2 807 269 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00131 1579 271 270 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00132 271 270 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00133 3 807 270 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00134 1 807 271 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00135 1579 273 272 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00136 273 272 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00137 4 825 272 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00138 2 825 273 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00139 1579 275 274 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00140 275 274 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00141 3 825 274 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00142 1 825 275 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00143 1579 277 276 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00144 277 276 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00145 4 819 276 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00146 2 819 277 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00147 1579 279 278 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00148 279 278 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00149 3 819 278 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00150 1 819 279 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00151 1579 281 280 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00152 281 280 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00153 4 821 280 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00154 2 821 281 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00155 1579 283 282 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00156 283 282 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00157 3 821 282 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00158 1 821 283 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00159 1579 285 284 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00160 285 284 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00161 4 823 284 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00162 2 823 285 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00163 1579 287 286 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00164 287 286 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00165 3 823 286 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00166 1 823 287 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00167 1579 289 288 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00168 289 288 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00169 4 841 288 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00170 2 841 289 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00171 1579 291 290 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00172 291 290 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00173 3 841 290 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00174 1 841 291 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00175 1579 293 292 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00176 293 292 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00177 4 835 292 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00178 2 835 293 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00179 1579 295 294 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00180 295 294 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00181 3 835 294 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00182 1 835 295 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00183 1579 297 296 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00184 297 296 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00185 4 837 296 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00186 2 837 297 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00187 1579 299 298 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00188 299 298 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00189 3 837 298 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00190 1 837 299 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00191 1579 301 300 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00192 301 300 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00193 4 839 300 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00194 2 839 301 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00195 1579 303 302 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00196 303 302 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00197 3 839 302 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00198 1 839 303 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00199 1579 305 304 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00200 305 304 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00201 4 857 304 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00202 2 857 305 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00203 1579 307 306 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00204 307 306 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00205 3 857 306 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00206 1 857 307 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00207 1579 309 308 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00208 309 308 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00209 4 851 308 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00210 2 851 309 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00211 1579 311 310 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00212 311 310 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00213 3 851 310 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00214 1 851 311 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00215 1579 313 312 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00216 313 312 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00217 4 853 312 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00218 2 853 313 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00219 1579 315 314 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00220 315 314 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00221 3 853 314 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00222 1 853 315 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00223 1579 317 316 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00224 317 316 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00225 4 855 316 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00226 2 855 317 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00227 1579 319 318 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00228 319 318 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00229 3 855 318 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00230 1 855 319 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00231 1579 321 320 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00232 321 320 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00233 4 873 320 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00234 2 873 321 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00235 1579 323 322 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00236 323 322 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00237 3 873 322 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00238 1 873 323 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00239 1579 325 324 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00240 325 324 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00241 4 867 324 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00242 2 867 325 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00243 1579 327 326 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00244 327 326 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00245 3 867 326 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00246 1 867 327 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00247 1579 329 328 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00248 329 328 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00249 4 869 328 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00250 2 869 329 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00251 1579 331 330 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00252 331 330 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00253 3 869 330 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00254 1 869 331 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00255 1579 333 332 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00256 333 332 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00257 4 871 332 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00258 2 871 333 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00259 1579 335 334 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00260 335 334 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00261 3 871 334 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00262 1 871 335 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00263 1579 337 336 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00264 337 336 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00265 4 889 336 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00266 2 889 337 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00267 1579 339 338 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00268 339 338 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00269 3 889 338 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00270 1 889 339 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00271 1579 341 340 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00272 341 340 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00273 4 883 340 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00274 2 883 341 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00275 1579 343 342 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00276 343 342 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00277 3 883 342 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00278 1 883 343 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00279 1579 345 344 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00280 345 344 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00281 4 885 344 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00282 2 885 345 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00283 1579 347 346 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00284 347 346 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00285 3 885 346 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00286 1 885 347 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00287 1579 349 348 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00288 349 348 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00289 4 887 348 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00290 2 887 349 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00291 1579 351 350 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00292 351 350 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00293 3 887 350 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00294 1 887 351 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00295 1579 353 352 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00296 353 352 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00297 4 905 352 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00298 2 905 353 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00299 1579 355 354 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00300 355 354 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00301 3 905 354 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00302 1 905 355 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00303 1579 357 356 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00304 357 356 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00305 4 899 356 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00306 2 899 357 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00307 1579 359 358 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00308 359 358 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00309 3 899 358 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00310 1 899 359 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00311 1579 361 360 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00312 361 360 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00313 4 901 360 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00314 2 901 361 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00315 1579 363 362 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00316 363 362 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00317 3 901 362 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00318 1 901 363 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00319 1579 365 364 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00320 365 364 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00321 4 903 364 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00322 2 903 365 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00323 1579 367 366 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00324 367 366 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00325 3 903 366 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00326 1 903 367 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00327 1579 369 368 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00328 369 368 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00329 4 921 368 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00330 2 921 369 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00331 1579 371 370 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00332 371 370 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00333 3 921 370 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00334 1 921 371 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00335 1579 373 372 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00336 373 372 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00337 4 915 372 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00338 2 915 373 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00339 1579 375 374 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00340 375 374 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00341 3 915 374 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00342 1 915 375 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00343 1579 377 376 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00344 377 376 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00345 4 917 376 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00346 2 917 377 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00347 1579 379 378 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00348 379 378 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00349 3 917 378 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00350 1 917 379 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00351 1579 381 380 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00352 381 380 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00353 4 919 380 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00354 2 919 381 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00355 1579 383 382 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00356 383 382 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00357 3 919 382 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00358 1 919 383 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00359 1579 385 384 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00360 385 384 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00361 4 937 384 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00362 2 937 385 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00363 1579 387 386 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00364 387 386 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00365 3 937 386 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00366 1 937 387 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00367 1579 389 388 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00368 389 388 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00369 4 931 388 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00370 2 931 389 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00371 1579 391 390 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00372 391 390 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00373 3 931 390 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00374 1 931 391 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00375 1579 393 392 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00376 393 392 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00377 4 933 392 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00378 2 933 393 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00379 1579 395 394 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00380 395 394 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00381 3 933 394 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00382 1 933 395 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00383 1579 397 396 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00384 397 396 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00385 4 935 396 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00386 2 935 397 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00387 1579 399 398 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00388 399 398 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00389 3 935 398 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00390 1 935 399 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00391 1579 401 400 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00392 401 400 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00393 4 953 400 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00394 2 953 401 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00395 1579 403 402 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00396 403 402 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00397 3 953 402 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00398 1 953 403 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00399 1579 405 404 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00400 405 404 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00401 4 947 404 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00402 2 947 405 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00403 1579 407 406 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00404 407 406 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00405 3 947 406 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00406 1 947 407 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00407 1579 409 408 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00408 409 408 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00409 4 949 408 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00410 2 949 409 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00411 1579 411 410 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00412 411 410 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00413 3 949 410 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00414 1 949 411 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00415 1579 413 412 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00416 413 412 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00417 4 951 412 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00418 2 951 413 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00419 1579 415 414 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00420 415 414 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00421 3 951 414 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00422 1 951 415 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00423 1579 417 416 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00424 417 416 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00425 4 969 416 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00426 2 969 417 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00427 1579 419 418 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00428 419 418 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00429 3 969 418 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00430 1 969 419 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00431 1579 421 420 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00432 421 420 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00433 4 963 420 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00434 2 963 421 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00435 1579 423 422 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00436 423 422 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00437 3 963 422 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00438 1 963 423 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00439 1579 425 424 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00440 425 424 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00441 4 965 424 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00442 2 965 425 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00443 1579 427 426 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00444 427 426 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00445 3 965 426 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00446 1 965 427 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00447 1579 429 428 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00448 429 428 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00449 4 967 428 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00450 2 967 429 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00451 1579 431 430 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00452 431 430 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00453 3 967 430 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00454 1 967 431 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00455 1579 433 432 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00456 433 432 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00457 4 985 432 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00458 2 985 433 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00459 1579 435 434 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00460 435 434 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00461 3 985 434 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00462 1 985 435 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00463 1579 437 436 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00464 437 436 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00465 4 979 436 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00466 2 979 437 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00467 1579 439 438 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00468 439 438 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00469 3 979 438 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00470 1 979 439 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00471 1579 441 440 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00472 441 440 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00473 4 981 440 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00474 2 981 441 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00475 1579 443 442 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00476 443 442 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00477 3 981 442 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00478 1 981 443 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00479 1579 445 444 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00480 445 444 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00481 4 983 444 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00482 2 983 445 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00483 1579 447 446 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00484 447 446 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00485 3 983 446 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00486 1 983 447 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00487 1579 449 448 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00488 449 448 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00489 4 1001 448 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00490 2 1001 449 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00491 1579 451 450 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00492 451 450 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00493 3 1001 450 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00494 1 1001 451 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00495 1579 453 452 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00496 453 452 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00497 4 995 452 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00498 2 995 453 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00499 1579 455 454 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00500 455 454 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00501 3 995 454 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00502 1 995 455 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00503 1579 457 456 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00504 457 456 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00505 4 997 456 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00506 2 997 457 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00507 1579 459 458 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00508 459 458 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00509 3 997 458 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00510 1 997 459 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00511 1579 461 460 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00512 461 460 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00513 4 999 460 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00514 2 999 461 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00515 1579 463 462 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00516 463 462 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00517 3 999 462 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00518 1 999 463 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00519 1 1003 8 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_00520 8 1004 2 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_00521 3 1003 9 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_00522 9 1004 4 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_00523 467 1038 465 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_00524 472 467 5 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00525 5 1029 1579 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00526 5 465 464 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00527 1579 1029 6 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00528 466 9 6 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00529 6 8 465 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00530 467 9 7 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00531 7 1029 1579 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00532 7 8 468 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00533 1580 1038 9 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_00534 9 1038 1580 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_00535 1580 1038 8 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_00536 8 1038 1580 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_00537 469 1032 9 1579 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_00538 8 1032 470 1579 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_00539 9 1038 8 1579 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_00540 1579 1585 469 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_00541 470 471 1579 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_00542 469 1585 1579 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_00543 1579 471 470 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_00544 1579 1585 471 1579 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00545 1585 473 1579 1579 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00546 1579 473 1585 1579 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00547 1579 1032 473 1579 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00548 473 472 1579 1579 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00549 473 1029 474 1579 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00550 13 743 11 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00551 13 743 1580 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00552 11 743 1580 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00553 12 743 10 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00554 1580 743 12 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00555 1580 743 10 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00556 1579 476 475 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00557 476 475 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00558 13 761 475 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00559 11 761 476 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00560 1579 478 477 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00561 478 477 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00562 12 761 477 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00563 10 761 478 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00564 1579 480 479 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00565 480 479 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00566 13 755 479 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00567 11 755 480 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00568 1579 482 481 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00569 482 481 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00570 12 755 481 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00571 10 755 482 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00572 1579 484 483 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00573 484 483 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00574 13 757 483 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00575 11 757 484 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00576 1579 486 485 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00577 486 485 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00578 12 757 485 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00579 10 757 486 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00580 1579 488 487 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00581 488 487 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00582 13 759 487 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00583 11 759 488 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00584 1579 490 489 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00585 490 489 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00586 12 759 489 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00587 10 759 490 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00588 1579 492 491 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00589 492 491 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00590 13 777 491 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00591 11 777 492 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00592 1579 494 493 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00593 494 493 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00594 12 777 493 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00595 10 777 494 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00596 1579 496 495 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00597 496 495 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00598 13 771 495 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00599 11 771 496 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00600 1579 498 497 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00601 498 497 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00602 12 771 497 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00603 10 771 498 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00604 1579 500 499 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00605 500 499 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00606 13 773 499 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00607 11 773 500 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00608 1579 502 501 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00609 502 501 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00610 12 773 501 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00611 10 773 502 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00612 1579 504 503 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00613 504 503 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00614 13 775 503 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00615 11 775 504 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00616 1579 506 505 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00617 506 505 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00618 12 775 505 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00619 10 775 506 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00620 1579 508 507 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00621 508 507 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00622 13 793 507 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00623 11 793 508 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00624 1579 510 509 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00625 510 509 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00626 12 793 509 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00627 10 793 510 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00628 1579 512 511 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00629 512 511 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00630 13 787 511 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00631 11 787 512 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00632 1579 514 513 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00633 514 513 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00634 12 787 513 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00635 10 787 514 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00636 1579 516 515 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00637 516 515 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00638 13 789 515 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00639 11 789 516 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00640 1579 518 517 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00641 518 517 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00642 12 789 517 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00643 10 789 518 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00644 1579 520 519 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00645 520 519 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00646 13 791 519 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00647 11 791 520 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00648 1579 522 521 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00649 522 521 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00650 12 791 521 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00651 10 791 522 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00652 1579 524 523 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00653 524 523 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00654 13 809 523 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00655 11 809 524 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00656 1579 526 525 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00657 526 525 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00658 12 809 525 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00659 10 809 526 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00660 1579 528 527 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00661 528 527 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00662 13 803 527 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00663 11 803 528 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00664 1579 530 529 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00665 530 529 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00666 12 803 529 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00667 10 803 530 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00668 1579 532 531 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00669 532 531 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00670 13 805 531 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00671 11 805 532 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00672 1579 534 533 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00673 534 533 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00674 12 805 533 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00675 10 805 534 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00676 1579 536 535 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00677 536 535 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00678 13 807 535 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00679 11 807 536 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00680 1579 538 537 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00681 538 537 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00682 12 807 537 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00683 10 807 538 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00684 1579 540 539 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00685 540 539 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00686 13 825 539 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00687 11 825 540 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00688 1579 542 541 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00689 542 541 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00690 12 825 541 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00691 10 825 542 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00692 1579 544 543 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00693 544 543 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00694 13 819 543 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00695 11 819 544 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00696 1579 546 545 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00697 546 545 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00698 12 819 545 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00699 10 819 546 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00700 1579 548 547 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00701 548 547 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00702 13 821 547 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00703 11 821 548 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00704 1579 550 549 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00705 550 549 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00706 12 821 549 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00707 10 821 550 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00708 1579 552 551 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00709 552 551 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00710 13 823 551 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00711 11 823 552 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00712 1579 554 553 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00713 554 553 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00714 12 823 553 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00715 10 823 554 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00716 1579 556 555 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00717 556 555 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00718 13 841 555 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00719 11 841 556 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00720 1579 558 557 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00721 558 557 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00722 12 841 557 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00723 10 841 558 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00724 1579 560 559 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00725 560 559 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00726 13 835 559 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00727 11 835 560 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00728 1579 562 561 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00729 562 561 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00730 12 835 561 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00731 10 835 562 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00732 1579 564 563 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00733 564 563 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00734 13 837 563 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00735 11 837 564 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00736 1579 566 565 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00737 566 565 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00738 12 837 565 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00739 10 837 566 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00740 1579 568 567 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00741 568 567 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00742 13 839 567 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00743 11 839 568 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00744 1579 570 569 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00745 570 569 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00746 12 839 569 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00747 10 839 570 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00748 1579 572 571 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00749 572 571 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00750 13 857 571 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00751 11 857 572 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00752 1579 574 573 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00753 574 573 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00754 12 857 573 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00755 10 857 574 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00756 1579 576 575 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00757 576 575 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00758 13 851 575 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00759 11 851 576 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00760 1579 578 577 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00761 578 577 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00762 12 851 577 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00763 10 851 578 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00764 1579 580 579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00765 580 579 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00766 13 853 579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00767 11 853 580 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00768 1579 582 581 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00769 582 581 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00770 12 853 581 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00771 10 853 582 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00772 1579 584 583 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00773 584 583 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00774 13 855 583 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00775 11 855 584 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00776 1579 586 585 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00777 586 585 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00778 12 855 585 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00779 10 855 586 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00780 1579 588 587 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00781 588 587 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00782 13 873 587 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00783 11 873 588 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00784 1579 590 589 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00785 590 589 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00786 12 873 589 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00787 10 873 590 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00788 1579 592 591 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00789 592 591 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00790 13 867 591 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00791 11 867 592 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00792 1579 594 593 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00793 594 593 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00794 12 867 593 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00795 10 867 594 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00796 1579 596 595 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00797 596 595 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00798 13 869 595 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00799 11 869 596 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00800 1579 598 597 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00801 598 597 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00802 12 869 597 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00803 10 869 598 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00804 1579 600 599 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00805 600 599 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00806 13 871 599 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00807 11 871 600 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00808 1579 602 601 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00809 602 601 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00810 12 871 601 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00811 10 871 602 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00812 1579 604 603 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00813 604 603 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00814 13 889 603 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00815 11 889 604 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00816 1579 606 605 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00817 606 605 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00818 12 889 605 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00819 10 889 606 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00820 1579 608 607 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00821 608 607 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00822 13 883 607 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00823 11 883 608 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00824 1579 610 609 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00825 610 609 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00826 12 883 609 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00827 10 883 610 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00828 1579 612 611 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00829 612 611 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00830 13 885 611 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00831 11 885 612 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00832 1579 614 613 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00833 614 613 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00834 12 885 613 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00835 10 885 614 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00836 1579 616 615 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00837 616 615 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00838 13 887 615 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00839 11 887 616 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00840 1579 618 617 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00841 618 617 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00842 12 887 617 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00843 10 887 618 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00844 1579 620 619 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00845 620 619 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00846 13 905 619 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00847 11 905 620 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00848 1579 622 621 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00849 622 621 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00850 12 905 621 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00851 10 905 622 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00852 1579 624 623 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00853 624 623 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00854 13 899 623 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00855 11 899 624 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00856 1579 626 625 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00857 626 625 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00858 12 899 625 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00859 10 899 626 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00860 1579 628 627 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00861 628 627 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00862 13 901 627 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00863 11 901 628 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00864 1579 630 629 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00865 630 629 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00866 12 901 629 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00867 10 901 630 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00868 1579 632 631 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00869 632 631 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00870 13 903 631 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00871 11 903 632 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00872 1579 634 633 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00873 634 633 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00874 12 903 633 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00875 10 903 634 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00876 1579 636 635 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00877 636 635 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00878 13 921 635 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00879 11 921 636 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00880 1579 638 637 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00881 638 637 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00882 12 921 637 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00883 10 921 638 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00884 1579 640 639 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00885 640 639 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00886 13 915 639 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00887 11 915 640 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00888 1579 642 641 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00889 642 641 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00890 12 915 641 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00891 10 915 642 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00892 1579 644 643 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00893 644 643 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00894 13 917 643 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00895 11 917 644 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00896 1579 646 645 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00897 646 645 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00898 12 917 645 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00899 10 917 646 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00900 1579 648 647 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00901 648 647 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00902 13 919 647 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00903 11 919 648 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00904 1579 650 649 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00905 650 649 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00906 12 919 649 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00907 10 919 650 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00908 1579 652 651 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00909 652 651 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00910 13 937 651 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00911 11 937 652 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00912 1579 654 653 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00913 654 653 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00914 12 937 653 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00915 10 937 654 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00916 1579 656 655 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00917 656 655 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00918 13 931 655 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00919 11 931 656 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00920 1579 658 657 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00921 658 657 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00922 12 931 657 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00923 10 931 658 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00924 1579 660 659 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00925 660 659 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00926 13 933 659 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00927 11 933 660 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00928 1579 662 661 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00929 662 661 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00930 12 933 661 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00931 10 933 662 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00932 1579 664 663 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00933 664 663 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00934 13 935 663 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00935 11 935 664 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00936 1579 666 665 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00937 666 665 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00938 12 935 665 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00939 10 935 666 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00940 1579 668 667 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00941 668 667 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00942 13 953 667 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00943 11 953 668 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00944 1579 670 669 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00945 670 669 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00946 12 953 669 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00947 10 953 670 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00948 1579 672 671 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00949 672 671 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00950 13 947 671 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00951 11 947 672 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00952 1579 674 673 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00953 674 673 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00954 12 947 673 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00955 10 947 674 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00956 1579 676 675 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00957 676 675 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00958 13 949 675 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00959 11 949 676 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00960 1579 678 677 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00961 678 677 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00962 12 949 677 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00963 10 949 678 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00964 1579 680 679 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00965 680 679 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00966 13 951 679 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00967 11 951 680 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00968 1579 682 681 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00969 682 681 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00970 12 951 681 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00971 10 951 682 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00972 1579 684 683 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00973 684 683 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00974 13 969 683 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00975 11 969 684 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00976 1579 686 685 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00977 686 685 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00978 12 969 685 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00979 10 969 686 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00980 1579 688 687 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00981 688 687 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00982 13 963 687 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00983 11 963 688 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00984 1579 690 689 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00985 690 689 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00986 12 963 689 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00987 10 963 690 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00988 1579 692 691 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00989 692 691 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00990 13 965 691 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00991 11 965 692 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00992 1579 694 693 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00993 694 693 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00994 12 965 693 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00995 10 965 694 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00996 1579 696 695 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00997 696 695 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00998 13 967 695 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00999 11 967 696 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01000 1579 698 697 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01001 698 697 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01002 12 967 697 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01003 10 967 698 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01004 1579 700 699 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01005 700 699 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01006 13 985 699 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01007 11 985 700 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01008 1579 702 701 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01009 702 701 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01010 12 985 701 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01011 10 985 702 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01012 1579 704 703 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01013 704 703 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01014 13 979 703 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01015 11 979 704 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01016 1579 706 705 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01017 706 705 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01018 12 979 705 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01019 10 979 706 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01020 1579 708 707 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01021 708 707 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01022 13 981 707 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01023 11 981 708 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01024 1579 710 709 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01025 710 709 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01026 12 981 709 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01027 10 981 710 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01028 1579 712 711 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01029 712 711 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01030 13 983 711 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01031 11 983 712 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01032 1579 714 713 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01033 714 713 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01034 12 983 713 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01035 10 983 714 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01036 1579 716 715 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01037 716 715 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01038 13 1001 715 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01039 11 1001 716 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01040 1579 718 717 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01041 718 717 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01042 12 1001 717 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01043 10 1001 718 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01044 1579 720 719 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01045 720 719 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01046 13 995 719 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01047 11 995 720 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01048 1579 722 721 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01049 722 721 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01050 12 995 721 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01051 10 995 722 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01052 1579 724 723 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01053 724 723 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01054 13 997 723 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01055 11 997 724 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01056 1579 726 725 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01057 726 725 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01058 12 997 725 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01059 10 997 726 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01060 1579 728 727 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01061 728 727 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01062 13 999 727 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01063 11 999 728 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01064 1579 730 729 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01065 730 729 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01066 12 999 729 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01067 10 999 730 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01068 10 1003 17 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01069 17 1004 11 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01070 12 1003 18 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01071 18 1004 13 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01072 734 1038 732 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01073 739 734 14 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01074 14 1029 1579 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01075 14 732 731 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01076 1579 1029 15 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01077 733 18 15 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01078 15 17 732 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01079 734 18 16 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01080 16 1029 1579 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01081 16 17 735 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01082 1580 1038 18 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01083 18 1038 1580 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01084 1580 1038 17 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01085 17 1038 1580 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01086 736 1032 18 1579 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_01087 17 1032 737 1579 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_01088 18 1038 17 1579 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_01089 1579 1584 736 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_01090 737 738 1579 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_01091 736 1584 1579 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_01092 1579 738 737 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_01093 1579 1584 738 1579 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01094 1584 740 1579 1579 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01095 1579 740 1584 1579 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01096 1579 1032 740 1579 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01097 740 739 1579 1579 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01098 740 1029 741 1579 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01099 742 744 1579 1579 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_01100 1579 744 742 1579 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_01101 742 744 1579 1579 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_01102 1579 744 742 1579 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_01103 743 746 1579 1579 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_01104 1579 746 743 1579 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_01105 743 746 1579 1579 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_01106 1579 746 743 1579 tn L=1U W=47U AS=94P AD=94P PS=98U PD=98U 
Mtr_01107 1579 1040 745 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01108 19 745 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01109 744 1041 19 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01110 20 745 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01111 746 1041 20 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01112 1579 762 750 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01113 754 760 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01114 1579 760 754 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01115 1579 758 752 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01116 752 758 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01117 1579 756 751 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01118 751 756 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01119 750 762 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01120 1579 747 753 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01121 753 749 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01122 21 1026 22 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01123 762 1040 21 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01124 22 753 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01125 23 1022 24 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01126 756 1040 23 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01127 24 753 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01128 25 1023 26 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01129 1579 753 25 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01130 26 1040 758 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01131 27 1040 760 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01132 1579 753 28 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01133 28 1019 27 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01134 29 1015 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01135 747 1012 29 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01136 1579 1006 30 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01137 30 1009 749 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01138 757 758 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01139 1579 758 757 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01140 759 760 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01141 1579 760 759 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01142 761 762 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01143 1579 762 761 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01144 755 756 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01145 1579 756 755 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01146 1579 778 766 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01147 770 776 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01148 1579 776 770 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01149 1579 774 768 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01150 768 774 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01151 1579 772 767 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01152 767 772 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01153 766 778 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01154 1579 763 769 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01155 769 765 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01156 31 1026 32 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01157 778 1040 31 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01158 32 769 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01159 33 1022 34 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01160 772 1040 33 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01161 34 769 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01162 35 1023 36 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01163 1579 769 35 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01164 36 1040 774 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01165 37 1040 776 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01166 1579 769 38 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01167 38 1019 37 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01168 39 1015 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01169 763 1012 39 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01170 1579 1005 40 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01171 40 1009 765 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01172 773 774 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01173 1579 774 773 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01174 775 776 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01175 1579 776 775 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01176 777 778 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01177 1579 778 777 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01178 771 772 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01179 1579 772 771 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01180 1579 794 782 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01181 786 792 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01182 1579 792 786 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01183 1579 790 784 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01184 784 790 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01185 1579 788 783 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01186 783 788 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01187 782 794 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01188 1579 779 785 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01189 785 781 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01190 41 1026 42 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01191 794 1040 41 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01192 42 785 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01193 43 1022 44 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01194 788 1040 43 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01195 44 785 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01196 45 1023 46 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01197 1579 785 45 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01198 46 1040 790 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01199 47 1040 792 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01200 1579 785 48 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01201 48 1019 47 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01202 49 1015 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01203 779 1012 49 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01204 1579 1006 50 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01205 50 1008 781 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01206 789 790 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01207 1579 790 789 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01208 791 792 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01209 1579 792 791 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01210 793 794 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01211 1579 794 793 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01212 787 788 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01213 1579 788 787 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01214 1579 810 798 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01215 802 808 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01216 1579 808 802 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01217 1579 806 800 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01218 800 806 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01219 1579 804 799 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01220 799 804 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01221 798 810 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01222 1579 795 801 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01223 801 797 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01224 51 1026 52 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01225 810 1040 51 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01226 52 801 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01227 53 1022 54 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01228 804 1040 53 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01229 54 801 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01230 55 1023 56 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01231 1579 801 55 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01232 56 1040 806 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01233 57 1040 808 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01234 1579 801 58 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01235 58 1019 57 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01236 59 1015 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01237 795 1012 59 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01238 1579 1005 60 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01239 60 1008 797 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01240 805 806 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01241 1579 806 805 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01242 807 808 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01243 1579 808 807 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01244 809 810 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01245 1579 810 809 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01246 803 804 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01247 1579 804 803 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01248 1579 826 814 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01249 818 824 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01250 1579 824 818 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01251 1579 822 816 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01252 816 822 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01253 1579 820 815 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01254 815 820 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01255 814 826 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01256 1579 811 817 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01257 817 813 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01258 61 1026 62 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01259 826 1040 61 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01260 62 817 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01261 63 1022 64 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01262 820 1040 63 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01263 64 817 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01264 65 1023 66 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01265 1579 817 65 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01266 66 1040 822 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01267 67 1040 824 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01268 1579 817 68 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01269 68 1019 67 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01270 69 1015 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01271 811 1011 69 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01272 1579 1006 70 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01273 70 1009 813 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01274 821 822 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01275 1579 822 821 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01276 823 824 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01277 1579 824 823 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01278 825 826 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01279 1579 826 825 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01280 819 820 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01281 1579 820 819 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01282 1579 842 830 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01283 834 840 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01284 1579 840 834 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01285 1579 838 832 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01286 832 838 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01287 1579 836 831 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01288 831 836 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01289 830 842 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01290 1579 827 833 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01291 833 829 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01292 71 1026 72 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01293 842 1040 71 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01294 72 833 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01295 73 1022 74 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01296 836 1040 73 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01297 74 833 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01298 75 1023 76 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01299 1579 833 75 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01300 76 1040 838 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01301 77 1040 840 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01302 1579 833 78 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01303 78 1019 77 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01304 79 1015 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01305 827 1011 79 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01306 1579 1005 80 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01307 80 1009 829 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01308 837 838 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01309 1579 838 837 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01310 839 840 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01311 1579 840 839 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01312 841 842 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01313 1579 842 841 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01314 835 836 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01315 1579 836 835 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01316 1579 858 846 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01317 850 856 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01318 1579 856 850 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01319 1579 854 848 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01320 848 854 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01321 1579 852 847 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01322 847 852 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01323 846 858 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01324 1579 843 849 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01325 849 845 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01326 81 1026 82 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01327 858 1040 81 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01328 82 849 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01329 83 1022 84 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01330 852 1040 83 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01331 84 849 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01332 85 1023 86 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01333 1579 849 85 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01334 86 1040 854 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01335 87 1040 856 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01336 1579 849 88 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01337 88 1019 87 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01338 89 1015 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01339 843 1011 89 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01340 1579 1006 90 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01341 90 1008 845 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01342 853 854 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01343 1579 854 853 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01344 855 856 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01345 1579 856 855 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01346 857 858 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01347 1579 858 857 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01348 851 852 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01349 1579 852 851 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01350 1579 874 862 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01351 866 872 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01352 1579 872 866 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01353 1579 870 864 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01354 864 870 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01355 1579 868 863 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01356 863 868 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01357 862 874 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01358 1579 859 865 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01359 865 861 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01360 91 1026 92 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01361 874 1040 91 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01362 92 865 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01363 93 1022 94 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01364 868 1040 93 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01365 94 865 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01366 95 1023 96 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01367 1579 865 95 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01368 96 1040 870 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01369 97 1040 872 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01370 1579 865 98 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01371 98 1019 97 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01372 99 1015 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01373 859 1011 99 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01374 1579 1005 100 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01375 100 1008 861 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01376 869 870 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01377 1579 870 869 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01378 871 872 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01379 1579 872 871 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01380 873 874 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01381 1579 874 873 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01382 867 868 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01383 1579 868 867 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01384 1579 890 878 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01385 882 888 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01386 1579 888 882 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01387 1579 886 880 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01388 880 886 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01389 1579 884 879 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01390 879 884 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01391 878 890 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01392 1579 875 881 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01393 881 877 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01394 101 1026 102 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01395 890 1040 101 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01396 102 881 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01397 103 1022 104 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01398 884 1040 103 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01399 104 881 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01400 105 1023 106 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01401 1579 881 105 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01402 106 1040 886 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01403 107 1040 888 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01404 1579 881 108 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01405 108 1019 107 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01406 109 1014 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01407 875 1012 109 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01408 1579 1006 110 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01409 110 1009 877 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01410 885 886 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01411 1579 886 885 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01412 887 888 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01413 1579 888 887 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01414 889 890 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01415 1579 890 889 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01416 883 884 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01417 1579 884 883 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01418 1579 906 894 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01419 898 904 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01420 1579 904 898 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01421 1579 902 896 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01422 896 902 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01423 1579 900 895 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01424 895 900 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01425 894 906 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01426 1579 891 897 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01427 897 893 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01428 111 1026 112 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01429 906 1040 111 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01430 112 897 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01431 113 1022 114 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01432 900 1040 113 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01433 114 897 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01434 115 1023 116 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01435 1579 897 115 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01436 116 1040 902 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01437 117 1040 904 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01438 1579 897 118 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01439 118 1019 117 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01440 119 1014 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01441 891 1012 119 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01442 1579 1005 120 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01443 120 1009 893 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01444 901 902 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01445 1579 902 901 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01446 903 904 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01447 1579 904 903 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01448 905 906 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01449 1579 906 905 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01450 899 900 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01451 1579 900 899 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01452 1579 922 910 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01453 914 920 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01454 1579 920 914 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01455 1579 918 912 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01456 912 918 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01457 1579 916 911 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01458 911 916 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01459 910 922 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01460 1579 907 913 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01461 913 909 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01462 121 1026 122 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01463 922 1040 121 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01464 122 913 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01465 123 1022 124 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01466 916 1040 123 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01467 124 913 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01468 125 1023 126 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01469 1579 913 125 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01470 126 1040 918 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01471 127 1040 920 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01472 1579 913 128 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01473 128 1019 127 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01474 129 1014 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01475 907 1012 129 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01476 1579 1006 130 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01477 130 1008 909 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01478 917 918 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01479 1579 918 917 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01480 919 920 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01481 1579 920 919 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01482 921 922 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01483 1579 922 921 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01484 915 916 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01485 1579 916 915 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01486 1579 938 926 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01487 930 936 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01488 1579 936 930 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01489 1579 934 928 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01490 928 934 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01491 1579 932 927 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01492 927 932 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01493 926 938 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01494 1579 923 929 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01495 929 925 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01496 131 1026 132 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01497 938 1040 131 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01498 132 929 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01499 133 1022 134 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01500 932 1040 133 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01501 134 929 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01502 135 1023 136 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01503 1579 929 135 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01504 136 1040 934 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01505 137 1040 936 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01506 1579 929 138 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01507 138 1019 137 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01508 139 1014 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01509 923 1012 139 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01510 1579 1005 140 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01511 140 1008 925 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01512 933 934 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01513 1579 934 933 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01514 935 936 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01515 1579 936 935 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01516 937 938 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01517 1579 938 937 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01518 931 932 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01519 1579 932 931 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01520 1579 954 942 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01521 946 952 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01522 1579 952 946 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01523 1579 950 944 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01524 944 950 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01525 1579 948 943 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01526 943 948 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01527 942 954 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01528 1579 939 945 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01529 945 941 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01530 141 1026 142 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01531 954 1040 141 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01532 142 945 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01533 143 1022 144 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01534 948 1040 143 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01535 144 945 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01536 145 1023 146 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01537 1579 945 145 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01538 146 1040 950 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01539 147 1040 952 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01540 1579 945 148 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01541 148 1019 147 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01542 149 1014 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01543 939 1011 149 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01544 1579 1006 150 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01545 150 1009 941 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01546 949 950 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01547 1579 950 949 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01548 951 952 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01549 1579 952 951 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01550 953 954 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01551 1579 954 953 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01552 947 948 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01553 1579 948 947 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01554 1579 970 958 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01555 962 968 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01556 1579 968 962 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01557 1579 966 960 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01558 960 966 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01559 1579 964 959 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01560 959 964 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01561 958 970 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01562 1579 955 961 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01563 961 957 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01564 151 1026 152 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01565 970 1040 151 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01566 152 961 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01567 153 1022 154 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01568 964 1040 153 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01569 154 961 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01570 155 1023 156 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01571 1579 961 155 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01572 156 1040 966 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01573 157 1040 968 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01574 1579 961 158 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01575 158 1019 157 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01576 159 1014 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01577 955 1011 159 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01578 1579 1005 160 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01579 160 1009 957 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01580 965 966 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01581 1579 966 965 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01582 967 968 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01583 1579 968 967 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01584 969 970 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01585 1579 970 969 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01586 963 964 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01587 1579 964 963 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01588 1579 986 974 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01589 978 984 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01590 1579 984 978 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01591 1579 982 976 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01592 976 982 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01593 1579 980 975 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01594 975 980 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01595 974 986 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01596 1579 971 977 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01597 977 973 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01598 161 1026 162 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01599 986 1040 161 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01600 162 977 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01601 163 1022 164 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01602 980 1040 163 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01603 164 977 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01604 165 1023 166 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01605 1579 977 165 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01606 166 1040 982 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01607 167 1040 984 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01608 1579 977 168 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01609 168 1019 167 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01610 169 1014 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01611 971 1011 169 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01612 1579 1006 170 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01613 170 1008 973 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01614 981 982 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01615 1579 982 981 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01616 983 984 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01617 1579 984 983 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01618 985 986 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01619 1579 986 985 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01620 979 980 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01621 1579 980 979 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01622 1579 1002 990 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01623 994 1000 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01624 1579 1000 994 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01625 1579 998 992 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01626 992 998 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01627 1579 996 991 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01628 991 996 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01629 990 1002 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01630 1579 987 993 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01631 993 989 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01632 171 1026 172 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01633 1002 1040 171 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01634 172 993 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01635 173 1022 174 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01636 996 1040 173 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01637 174 993 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01638 175 1023 176 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01639 1579 993 175 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01640 176 1040 998 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01641 177 1040 1000 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01642 1579 993 178 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01643 178 1019 177 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01644 179 1014 1579 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01645 987 1011 179 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01646 1579 1005 180 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01647 180 1008 989 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01648 997 998 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01649 1579 998 997 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01650 999 1000 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01651 1579 1000 999 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01652 1001 1002 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01653 1579 1002 1001 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01654 995 996 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01655 1579 996 995 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01656 1004 1028 1579 1579 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_01657 1579 1027 1003 1579 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_01658 1579 1007 1006 1579 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_01659 1005 1590 1579 1579 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_01660 1579 1590 1007 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01661 1579 1010 1009 1579 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_01662 1008 1589 1579 1579 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_01663 1579 1589 1010 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01664 1579 1013 1012 1579 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_01665 1011 1588 1579 1579 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_01666 1579 1588 1013 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01667 1579 1016 1015 1579 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_01668 1014 1587 1579 1579 tn L=1U W=30U AS=60P AD=60P PS=64U PD=64U 
Mtr_01669 1579 1587 1016 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_01670 1579 1592 1017 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01671 1579 1591 1018 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01672 1579 1592 181 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01673 181 1018 1024 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01674 1025 1592 182 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01675 182 1591 1579 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01676 1579 1017 183 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01677 183 1018 1020 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01678 1021 1017 184 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01679 184 1591 1579 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01680 1579 1020 1019 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01681 1022 1021 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01682 1579 1024 1023 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01683 1026 1025 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01684 1027 1028 1579 1579 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01685 1579 1593 1028 1579 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01686 1029 1030 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01687 1579 1030 1029 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01688 1030 1033 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01689 1573 1031 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01690 1579 1031 1573 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01691 1031 1034 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01692 1032 1033 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01693 1579 1033 1032 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01694 185 1040 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01695 1033 1578 185 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01696 1576 1034 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01697 1579 1034 1576 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01698 186 1040 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01699 1034 1578 186 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01700 1035 1039 187 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01701 187 1041 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01702 1579 1035 1036 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01703 1036 1035 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01704 1037 1039 188 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01705 188 1041 1579 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01706 1579 1037 1038 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01707 1038 1037 1579 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_01708 1579 1040 1039 1579 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01709 1040 1041 1579 1579 tn L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_01710 1579 1041 1040 1579 tn L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_01711 189 1586 1041 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01712 1579 1581 189 1579 tn L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_01713 193 742 191 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01714 193 742 1580 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01715 191 742 1580 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01716 192 742 190 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01717 1580 742 192 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01718 1580 742 190 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01719 1579 1043 1042 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01720 1043 1042 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01721 193 750 1042 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01722 191 750 1043 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01723 1579 1045 1044 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01724 1045 1044 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01725 192 750 1044 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01726 190 750 1045 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01727 1579 1047 1046 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01728 1047 1046 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01729 193 751 1046 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01730 191 751 1047 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01731 1579 1049 1048 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01732 1049 1048 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01733 192 751 1048 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01734 190 751 1049 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01735 1579 1051 1050 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01736 1051 1050 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01737 193 752 1050 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01738 191 752 1051 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01739 1579 1053 1052 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01740 1053 1052 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01741 192 752 1052 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01742 190 752 1053 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01743 1579 1055 1054 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01744 1055 1054 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01745 193 754 1054 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01746 191 754 1055 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01747 1579 1057 1056 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01748 1057 1056 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01749 192 754 1056 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01750 190 754 1057 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01751 1579 1059 1058 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01752 1059 1058 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01753 193 766 1058 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01754 191 766 1059 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01755 1579 1061 1060 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01756 1061 1060 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01757 192 766 1060 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01758 190 766 1061 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01759 1579 1063 1062 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01760 1063 1062 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01761 193 767 1062 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01762 191 767 1063 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01763 1579 1065 1064 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01764 1065 1064 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01765 192 767 1064 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01766 190 767 1065 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01767 1579 1067 1066 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01768 1067 1066 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01769 193 768 1066 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01770 191 768 1067 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01771 1579 1069 1068 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01772 1069 1068 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01773 192 768 1068 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01774 190 768 1069 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01775 1579 1071 1070 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01776 1071 1070 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01777 193 770 1070 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01778 191 770 1071 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01779 1579 1073 1072 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01780 1073 1072 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01781 192 770 1072 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01782 190 770 1073 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01783 1579 1075 1074 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01784 1075 1074 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01785 193 782 1074 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01786 191 782 1075 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01787 1579 1077 1076 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01788 1077 1076 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01789 192 782 1076 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01790 190 782 1077 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01791 1579 1079 1078 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01792 1079 1078 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01793 193 783 1078 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01794 191 783 1079 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01795 1579 1081 1080 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01796 1081 1080 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01797 192 783 1080 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01798 190 783 1081 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01799 1579 1083 1082 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01800 1083 1082 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01801 193 784 1082 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01802 191 784 1083 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01803 1579 1085 1084 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01804 1085 1084 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01805 192 784 1084 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01806 190 784 1085 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01807 1579 1087 1086 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01808 1087 1086 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01809 193 786 1086 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01810 191 786 1087 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01811 1579 1089 1088 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01812 1089 1088 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01813 192 786 1088 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01814 190 786 1089 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01815 1579 1091 1090 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01816 1091 1090 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01817 193 798 1090 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01818 191 798 1091 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01819 1579 1093 1092 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01820 1093 1092 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01821 192 798 1092 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01822 190 798 1093 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01823 1579 1095 1094 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01824 1095 1094 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01825 193 799 1094 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01826 191 799 1095 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01827 1579 1097 1096 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01828 1097 1096 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01829 192 799 1096 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01830 190 799 1097 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01831 1579 1099 1098 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01832 1099 1098 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01833 193 800 1098 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01834 191 800 1099 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01835 1579 1101 1100 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01836 1101 1100 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01837 192 800 1100 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01838 190 800 1101 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01839 1579 1103 1102 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01840 1103 1102 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01841 193 802 1102 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01842 191 802 1103 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01843 1579 1105 1104 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01844 1105 1104 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01845 192 802 1104 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01846 190 802 1105 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01847 1579 1107 1106 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01848 1107 1106 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01849 193 814 1106 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01850 191 814 1107 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01851 1579 1109 1108 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01852 1109 1108 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01853 192 814 1108 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01854 190 814 1109 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01855 1579 1111 1110 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01856 1111 1110 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01857 193 815 1110 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01858 191 815 1111 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01859 1579 1113 1112 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01860 1113 1112 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01861 192 815 1112 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01862 190 815 1113 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01863 1579 1115 1114 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01864 1115 1114 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01865 193 816 1114 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01866 191 816 1115 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01867 1579 1117 1116 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01868 1117 1116 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01869 192 816 1116 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01870 190 816 1117 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01871 1579 1119 1118 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01872 1119 1118 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01873 193 818 1118 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01874 191 818 1119 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01875 1579 1121 1120 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01876 1121 1120 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01877 192 818 1120 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01878 190 818 1121 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01879 1579 1123 1122 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01880 1123 1122 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01881 193 830 1122 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01882 191 830 1123 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01883 1579 1125 1124 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01884 1125 1124 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01885 192 830 1124 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01886 190 830 1125 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01887 1579 1127 1126 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01888 1127 1126 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01889 193 831 1126 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01890 191 831 1127 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01891 1579 1129 1128 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01892 1129 1128 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01893 192 831 1128 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01894 190 831 1129 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01895 1579 1131 1130 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01896 1131 1130 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01897 193 832 1130 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01898 191 832 1131 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01899 1579 1133 1132 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01900 1133 1132 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01901 192 832 1132 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01902 190 832 1133 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01903 1579 1135 1134 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01904 1135 1134 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01905 193 834 1134 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01906 191 834 1135 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01907 1579 1137 1136 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01908 1137 1136 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01909 192 834 1136 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01910 190 834 1137 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01911 1579 1139 1138 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01912 1139 1138 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01913 193 846 1138 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01914 191 846 1139 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01915 1579 1141 1140 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01916 1141 1140 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01917 192 846 1140 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01918 190 846 1141 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01919 1579 1143 1142 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01920 1143 1142 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01921 193 847 1142 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01922 191 847 1143 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01923 1579 1145 1144 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01924 1145 1144 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01925 192 847 1144 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01926 190 847 1145 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01927 1579 1147 1146 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01928 1147 1146 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01929 193 848 1146 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01930 191 848 1147 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01931 1579 1149 1148 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01932 1149 1148 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01933 192 848 1148 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01934 190 848 1149 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01935 1579 1151 1150 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01936 1151 1150 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01937 193 850 1150 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01938 191 850 1151 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01939 1579 1153 1152 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01940 1153 1152 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01941 192 850 1152 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01942 190 850 1153 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01943 1579 1155 1154 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01944 1155 1154 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01945 193 862 1154 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01946 191 862 1155 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01947 1579 1157 1156 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01948 1157 1156 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01949 192 862 1156 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01950 190 862 1157 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01951 1579 1159 1158 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01952 1159 1158 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01953 193 863 1158 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01954 191 863 1159 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01955 1579 1161 1160 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01956 1161 1160 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01957 192 863 1160 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01958 190 863 1161 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01959 1579 1163 1162 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01960 1163 1162 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01961 193 864 1162 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01962 191 864 1163 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01963 1579 1165 1164 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01964 1165 1164 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01965 192 864 1164 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01966 190 864 1165 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01967 1579 1167 1166 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01968 1167 1166 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01969 193 866 1166 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01970 191 866 1167 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01971 1579 1169 1168 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01972 1169 1168 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01973 192 866 1168 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01974 190 866 1169 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01975 1579 1171 1170 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01976 1171 1170 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01977 193 878 1170 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01978 191 878 1171 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01979 1579 1173 1172 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01980 1173 1172 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01981 192 878 1172 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01982 190 878 1173 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01983 1579 1175 1174 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01984 1175 1174 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01985 193 879 1174 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01986 191 879 1175 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01987 1579 1177 1176 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01988 1177 1176 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01989 192 879 1176 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01990 190 879 1177 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01991 1579 1179 1178 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01992 1179 1178 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01993 193 880 1178 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01994 191 880 1179 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01995 1579 1181 1180 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01996 1181 1180 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01997 192 880 1180 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01998 190 880 1181 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01999 1579 1183 1182 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02000 1183 1182 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02001 193 882 1182 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02002 191 882 1183 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02003 1579 1185 1184 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02004 1185 1184 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02005 192 882 1184 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02006 190 882 1185 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02007 1579 1187 1186 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02008 1187 1186 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02009 193 894 1186 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02010 191 894 1187 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02011 1579 1189 1188 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02012 1189 1188 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02013 192 894 1188 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02014 190 894 1189 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02015 1579 1191 1190 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02016 1191 1190 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02017 193 895 1190 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02018 191 895 1191 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02019 1579 1193 1192 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02020 1193 1192 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02021 192 895 1192 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02022 190 895 1193 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02023 1579 1195 1194 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02024 1195 1194 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02025 193 896 1194 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02026 191 896 1195 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02027 1579 1197 1196 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02028 1197 1196 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02029 192 896 1196 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02030 190 896 1197 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02031 1579 1199 1198 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02032 1199 1198 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02033 193 898 1198 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02034 191 898 1199 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02035 1579 1201 1200 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02036 1201 1200 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02037 192 898 1200 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02038 190 898 1201 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02039 1579 1203 1202 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02040 1203 1202 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02041 193 910 1202 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02042 191 910 1203 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02043 1579 1205 1204 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02044 1205 1204 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02045 192 910 1204 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02046 190 910 1205 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02047 1579 1207 1206 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02048 1207 1206 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02049 193 911 1206 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02050 191 911 1207 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02051 1579 1209 1208 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02052 1209 1208 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02053 192 911 1208 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02054 190 911 1209 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02055 1579 1211 1210 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02056 1211 1210 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02057 193 912 1210 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02058 191 912 1211 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02059 1579 1213 1212 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02060 1213 1212 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02061 192 912 1212 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02062 190 912 1213 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02063 1579 1215 1214 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02064 1215 1214 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02065 193 914 1214 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02066 191 914 1215 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02067 1579 1217 1216 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02068 1217 1216 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02069 192 914 1216 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02070 190 914 1217 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02071 1579 1219 1218 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02072 1219 1218 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02073 193 926 1218 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02074 191 926 1219 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02075 1579 1221 1220 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02076 1221 1220 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02077 192 926 1220 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02078 190 926 1221 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02079 1579 1223 1222 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02080 1223 1222 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02081 193 927 1222 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02082 191 927 1223 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02083 1579 1225 1224 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02084 1225 1224 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02085 192 927 1224 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02086 190 927 1225 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02087 1579 1227 1226 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02088 1227 1226 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02089 193 928 1226 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02090 191 928 1227 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02091 1579 1229 1228 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02092 1229 1228 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02093 192 928 1228 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02094 190 928 1229 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02095 1579 1231 1230 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02096 1231 1230 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02097 193 930 1230 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02098 191 930 1231 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02099 1579 1233 1232 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02100 1233 1232 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02101 192 930 1232 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02102 190 930 1233 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02103 1579 1235 1234 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02104 1235 1234 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02105 193 942 1234 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02106 191 942 1235 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02107 1579 1237 1236 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02108 1237 1236 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02109 192 942 1236 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02110 190 942 1237 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02111 1579 1239 1238 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02112 1239 1238 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02113 193 943 1238 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02114 191 943 1239 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02115 1579 1241 1240 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02116 1241 1240 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02117 192 943 1240 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02118 190 943 1241 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02119 1579 1243 1242 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02120 1243 1242 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02121 193 944 1242 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02122 191 944 1243 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02123 1579 1245 1244 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02124 1245 1244 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02125 192 944 1244 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02126 190 944 1245 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02127 1579 1247 1246 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02128 1247 1246 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02129 193 946 1246 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02130 191 946 1247 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02131 1579 1249 1248 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02132 1249 1248 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02133 192 946 1248 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02134 190 946 1249 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02135 1579 1251 1250 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02136 1251 1250 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02137 193 958 1250 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02138 191 958 1251 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02139 1579 1253 1252 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02140 1253 1252 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02141 192 958 1252 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02142 190 958 1253 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02143 1579 1255 1254 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02144 1255 1254 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02145 193 959 1254 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02146 191 959 1255 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02147 1579 1257 1256 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02148 1257 1256 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02149 192 959 1256 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02150 190 959 1257 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02151 1579 1259 1258 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02152 1259 1258 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02153 193 960 1258 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02154 191 960 1259 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02155 1579 1261 1260 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02156 1261 1260 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02157 192 960 1260 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02158 190 960 1261 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02159 1579 1263 1262 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02160 1263 1262 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02161 193 962 1262 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02162 191 962 1263 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02163 1579 1265 1264 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02164 1265 1264 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02165 192 962 1264 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02166 190 962 1265 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02167 1579 1267 1266 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02168 1267 1266 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02169 193 974 1266 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02170 191 974 1267 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02171 1579 1269 1268 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02172 1269 1268 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02173 192 974 1268 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02174 190 974 1269 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02175 1579 1271 1270 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02176 1271 1270 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02177 193 975 1270 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02178 191 975 1271 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02179 1579 1273 1272 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02180 1273 1272 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02181 192 975 1272 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02182 190 975 1273 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02183 1579 1275 1274 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02184 1275 1274 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02185 193 976 1274 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02186 191 976 1275 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02187 1579 1277 1276 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02188 1277 1276 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02189 192 976 1276 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02190 190 976 1277 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02191 1579 1279 1278 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02192 1279 1278 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02193 193 978 1278 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02194 191 978 1279 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02195 1579 1281 1280 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02196 1281 1280 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02197 192 978 1280 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02198 190 978 1281 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02199 1579 1283 1282 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02200 1283 1282 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02201 193 990 1282 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02202 191 990 1283 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02203 1579 1285 1284 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02204 1285 1284 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02205 192 990 1284 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02206 190 990 1285 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02207 1579 1287 1286 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02208 1287 1286 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02209 193 991 1286 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02210 191 991 1287 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02211 1579 1289 1288 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02212 1289 1288 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02213 192 991 1288 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02214 190 991 1289 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02215 1579 1291 1290 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02216 1291 1290 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02217 193 992 1290 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02218 191 992 1291 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02219 1579 1293 1292 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02220 1293 1292 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02221 192 992 1292 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02222 190 992 1293 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02223 1579 1295 1294 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02224 1295 1294 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02225 193 994 1294 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02226 191 994 1295 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02227 1579 1297 1296 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02228 1297 1296 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02229 192 994 1296 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02230 190 994 1297 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02231 190 1003 197 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02232 197 1004 191 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02233 192 1003 198 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02234 198 1004 193 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02235 1301 1036 1299 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02236 1306 1301 194 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02237 194 1573 1579 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02238 194 1299 1298 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02239 1579 1573 195 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02240 1300 198 195 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02241 195 197 1299 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02242 1301 198 196 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02243 196 1573 1579 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02244 196 197 1302 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02245 1580 1036 198 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02246 198 1036 1580 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02247 1580 1036 197 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02248 197 1036 1580 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02249 1303 1576 198 1579 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_02250 197 1576 1304 1579 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_02251 198 1036 197 1579 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_02252 1579 1583 1303 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_02253 1304 1305 1579 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_02254 1303 1583 1579 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_02255 1579 1305 1304 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_02256 1579 1583 1305 1579 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02257 1583 1307 1579 1579 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02258 1579 1307 1583 1579 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02259 1579 1576 1307 1579 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02260 1307 1306 1579 1579 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02261 1307 1573 1308 1579 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02262 202 742 200 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02263 202 742 1580 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02264 200 742 1580 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02265 201 742 199 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02266 1580 742 201 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02267 1580 742 199 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02268 1579 1310 1309 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02269 1310 1309 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02270 202 750 1309 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02271 200 750 1310 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02272 1579 1312 1311 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02273 1312 1311 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02274 201 750 1311 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02275 199 750 1312 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02276 1579 1314 1313 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02277 1314 1313 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02278 202 751 1313 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02279 200 751 1314 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02280 1579 1316 1315 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02281 1316 1315 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02282 201 751 1315 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02283 199 751 1316 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02284 1579 1318 1317 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02285 1318 1317 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02286 202 752 1317 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02287 200 752 1318 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02288 1579 1320 1319 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02289 1320 1319 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02290 201 752 1319 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02291 199 752 1320 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02292 1579 1322 1321 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02293 1322 1321 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02294 202 754 1321 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02295 200 754 1322 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02296 1579 1324 1323 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02297 1324 1323 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02298 201 754 1323 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02299 199 754 1324 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02300 1579 1326 1325 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02301 1326 1325 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02302 202 766 1325 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02303 200 766 1326 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02304 1579 1328 1327 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02305 1328 1327 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02306 201 766 1327 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02307 199 766 1328 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02308 1579 1330 1329 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02309 1330 1329 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02310 202 767 1329 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02311 200 767 1330 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02312 1579 1332 1331 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02313 1332 1331 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02314 201 767 1331 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02315 199 767 1332 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02316 1579 1334 1333 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02317 1334 1333 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02318 202 768 1333 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02319 200 768 1334 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02320 1579 1336 1335 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02321 1336 1335 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02322 201 768 1335 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02323 199 768 1336 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02324 1579 1338 1337 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02325 1338 1337 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02326 202 770 1337 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02327 200 770 1338 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02328 1579 1340 1339 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02329 1340 1339 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02330 201 770 1339 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02331 199 770 1340 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02332 1579 1342 1341 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02333 1342 1341 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02334 202 782 1341 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02335 200 782 1342 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02336 1579 1344 1343 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02337 1344 1343 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02338 201 782 1343 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02339 199 782 1344 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02340 1579 1346 1345 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02341 1346 1345 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02342 202 783 1345 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02343 200 783 1346 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02344 1579 1348 1347 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02345 1348 1347 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02346 201 783 1347 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02347 199 783 1348 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02348 1579 1350 1349 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02349 1350 1349 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02350 202 784 1349 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02351 200 784 1350 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02352 1579 1352 1351 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02353 1352 1351 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02354 201 784 1351 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02355 199 784 1352 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02356 1579 1354 1353 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02357 1354 1353 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02358 202 786 1353 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02359 200 786 1354 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02360 1579 1356 1355 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02361 1356 1355 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02362 201 786 1355 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02363 199 786 1356 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02364 1579 1358 1357 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02365 1358 1357 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02366 202 798 1357 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02367 200 798 1358 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02368 1579 1360 1359 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02369 1360 1359 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02370 201 798 1359 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02371 199 798 1360 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02372 1579 1362 1361 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02373 1362 1361 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02374 202 799 1361 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02375 200 799 1362 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02376 1579 1364 1363 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02377 1364 1363 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02378 201 799 1363 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02379 199 799 1364 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02380 1579 1366 1365 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02381 1366 1365 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02382 202 800 1365 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02383 200 800 1366 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02384 1579 1368 1367 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02385 1368 1367 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02386 201 800 1367 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02387 199 800 1368 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02388 1579 1370 1369 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02389 1370 1369 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02390 202 802 1369 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02391 200 802 1370 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02392 1579 1372 1371 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02393 1372 1371 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02394 201 802 1371 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02395 199 802 1372 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02396 1579 1374 1373 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02397 1374 1373 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02398 202 814 1373 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02399 200 814 1374 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02400 1579 1376 1375 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02401 1376 1375 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02402 201 814 1375 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02403 199 814 1376 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02404 1579 1378 1377 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02405 1378 1377 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02406 202 815 1377 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02407 200 815 1378 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02408 1579 1380 1379 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02409 1380 1379 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02410 201 815 1379 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02411 199 815 1380 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02412 1579 1382 1381 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02413 1382 1381 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02414 202 816 1381 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02415 200 816 1382 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02416 1579 1384 1383 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02417 1384 1383 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02418 201 816 1383 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02419 199 816 1384 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02420 1579 1386 1385 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02421 1386 1385 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02422 202 818 1385 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02423 200 818 1386 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02424 1579 1388 1387 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02425 1388 1387 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02426 201 818 1387 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02427 199 818 1388 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02428 1579 1390 1389 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02429 1390 1389 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02430 202 830 1389 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02431 200 830 1390 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02432 1579 1392 1391 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02433 1392 1391 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02434 201 830 1391 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02435 199 830 1392 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02436 1579 1394 1393 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02437 1394 1393 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02438 202 831 1393 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02439 200 831 1394 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02440 1579 1396 1395 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02441 1396 1395 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02442 201 831 1395 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02443 199 831 1396 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02444 1579 1398 1397 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02445 1398 1397 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02446 202 832 1397 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02447 200 832 1398 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02448 1579 1400 1399 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02449 1400 1399 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02450 201 832 1399 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02451 199 832 1400 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02452 1579 1402 1401 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02453 1402 1401 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02454 202 834 1401 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02455 200 834 1402 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02456 1579 1404 1403 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02457 1404 1403 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02458 201 834 1403 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02459 199 834 1404 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02460 1579 1406 1405 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02461 1406 1405 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02462 202 846 1405 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02463 200 846 1406 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02464 1579 1408 1407 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02465 1408 1407 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02466 201 846 1407 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02467 199 846 1408 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02468 1579 1410 1409 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02469 1410 1409 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02470 202 847 1409 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02471 200 847 1410 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02472 1579 1412 1411 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02473 1412 1411 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02474 201 847 1411 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02475 199 847 1412 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02476 1579 1414 1413 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02477 1414 1413 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02478 202 848 1413 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02479 200 848 1414 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02480 1579 1416 1415 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02481 1416 1415 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02482 201 848 1415 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02483 199 848 1416 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02484 1579 1418 1417 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02485 1418 1417 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02486 202 850 1417 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02487 200 850 1418 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02488 1579 1420 1419 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02489 1420 1419 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02490 201 850 1419 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02491 199 850 1420 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02492 1579 1422 1421 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02493 1422 1421 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02494 202 862 1421 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02495 200 862 1422 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02496 1579 1424 1423 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02497 1424 1423 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02498 201 862 1423 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02499 199 862 1424 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02500 1579 1426 1425 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02501 1426 1425 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02502 202 863 1425 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02503 200 863 1426 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02504 1579 1428 1427 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02505 1428 1427 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02506 201 863 1427 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02507 199 863 1428 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02508 1579 1430 1429 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02509 1430 1429 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02510 202 864 1429 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02511 200 864 1430 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02512 1579 1432 1431 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02513 1432 1431 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02514 201 864 1431 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02515 199 864 1432 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02516 1579 1434 1433 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02517 1434 1433 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02518 202 866 1433 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02519 200 866 1434 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02520 1579 1436 1435 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02521 1436 1435 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02522 201 866 1435 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02523 199 866 1436 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02524 1579 1438 1437 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02525 1438 1437 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02526 202 878 1437 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02527 200 878 1438 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02528 1579 1440 1439 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02529 1440 1439 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02530 201 878 1439 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02531 199 878 1440 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02532 1579 1442 1441 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02533 1442 1441 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02534 202 879 1441 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02535 200 879 1442 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02536 1579 1444 1443 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02537 1444 1443 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02538 201 879 1443 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02539 199 879 1444 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02540 1579 1446 1445 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02541 1446 1445 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02542 202 880 1445 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02543 200 880 1446 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02544 1579 1448 1447 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02545 1448 1447 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02546 201 880 1447 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02547 199 880 1448 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02548 1579 1450 1449 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02549 1450 1449 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02550 202 882 1449 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02551 200 882 1450 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02552 1579 1452 1451 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02553 1452 1451 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02554 201 882 1451 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02555 199 882 1452 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02556 1579 1454 1453 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02557 1454 1453 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02558 202 894 1453 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02559 200 894 1454 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02560 1579 1456 1455 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02561 1456 1455 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02562 201 894 1455 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02563 199 894 1456 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02564 1579 1458 1457 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02565 1458 1457 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02566 202 895 1457 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02567 200 895 1458 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02568 1579 1460 1459 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02569 1460 1459 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02570 201 895 1459 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02571 199 895 1460 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02572 1579 1462 1461 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02573 1462 1461 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02574 202 896 1461 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02575 200 896 1462 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02576 1579 1464 1463 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02577 1464 1463 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02578 201 896 1463 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02579 199 896 1464 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02580 1579 1466 1465 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02581 1466 1465 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02582 202 898 1465 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02583 200 898 1466 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02584 1579 1468 1467 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02585 1468 1467 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02586 201 898 1467 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02587 199 898 1468 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02588 1579 1470 1469 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02589 1470 1469 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02590 202 910 1469 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02591 200 910 1470 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02592 1579 1472 1471 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02593 1472 1471 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02594 201 910 1471 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02595 199 910 1472 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02596 1579 1474 1473 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02597 1474 1473 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02598 202 911 1473 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02599 200 911 1474 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02600 1579 1476 1475 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02601 1476 1475 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02602 201 911 1475 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02603 199 911 1476 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02604 1579 1478 1477 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02605 1478 1477 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02606 202 912 1477 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02607 200 912 1478 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02608 1579 1480 1479 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02609 1480 1479 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02610 201 912 1479 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02611 199 912 1480 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02612 1579 1482 1481 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02613 1482 1481 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02614 202 914 1481 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02615 200 914 1482 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02616 1579 1484 1483 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02617 1484 1483 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02618 201 914 1483 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02619 199 914 1484 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02620 1579 1486 1485 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02621 1486 1485 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02622 202 926 1485 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02623 200 926 1486 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02624 1579 1488 1487 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02625 1488 1487 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02626 201 926 1487 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02627 199 926 1488 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02628 1579 1490 1489 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02629 1490 1489 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02630 202 927 1489 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02631 200 927 1490 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02632 1579 1492 1491 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02633 1492 1491 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02634 201 927 1491 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02635 199 927 1492 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02636 1579 1494 1493 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02637 1494 1493 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02638 202 928 1493 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02639 200 928 1494 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02640 1579 1496 1495 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02641 1496 1495 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02642 201 928 1495 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02643 199 928 1496 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02644 1579 1498 1497 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02645 1498 1497 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02646 202 930 1497 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02647 200 930 1498 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02648 1579 1500 1499 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02649 1500 1499 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02650 201 930 1499 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02651 199 930 1500 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02652 1579 1502 1501 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02653 1502 1501 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02654 202 942 1501 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02655 200 942 1502 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02656 1579 1504 1503 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02657 1504 1503 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02658 201 942 1503 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02659 199 942 1504 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02660 1579 1506 1505 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02661 1506 1505 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02662 202 943 1505 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02663 200 943 1506 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02664 1579 1508 1507 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02665 1508 1507 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02666 201 943 1507 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02667 199 943 1508 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02668 1579 1510 1509 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02669 1510 1509 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02670 202 944 1509 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02671 200 944 1510 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02672 1579 1512 1511 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02673 1512 1511 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02674 201 944 1511 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02675 199 944 1512 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02676 1579 1514 1513 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02677 1514 1513 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02678 202 946 1513 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02679 200 946 1514 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02680 1579 1516 1515 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02681 1516 1515 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02682 201 946 1515 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02683 199 946 1516 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02684 1579 1518 1517 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02685 1518 1517 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02686 202 958 1517 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02687 200 958 1518 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02688 1579 1520 1519 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02689 1520 1519 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02690 201 958 1519 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02691 199 958 1520 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02692 1579 1522 1521 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02693 1522 1521 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02694 202 959 1521 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02695 200 959 1522 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02696 1579 1524 1523 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02697 1524 1523 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02698 201 959 1523 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02699 199 959 1524 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02700 1579 1526 1525 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02701 1526 1525 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02702 202 960 1525 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02703 200 960 1526 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02704 1579 1528 1527 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02705 1528 1527 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02706 201 960 1527 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02707 199 960 1528 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02708 1579 1530 1529 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02709 1530 1529 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02710 202 962 1529 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02711 200 962 1530 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02712 1579 1532 1531 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02713 1532 1531 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02714 201 962 1531 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02715 199 962 1532 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02716 1579 1534 1533 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02717 1534 1533 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02718 202 974 1533 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02719 200 974 1534 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02720 1579 1536 1535 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02721 1536 1535 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02722 201 974 1535 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02723 199 974 1536 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02724 1579 1538 1537 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02725 1538 1537 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02726 202 975 1537 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02727 200 975 1538 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02728 1579 1540 1539 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02729 1540 1539 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02730 201 975 1539 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02731 199 975 1540 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02732 1579 1542 1541 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02733 1542 1541 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02734 202 976 1541 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02735 200 976 1542 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02736 1579 1544 1543 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02737 1544 1543 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02738 201 976 1543 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02739 199 976 1544 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02740 1579 1546 1545 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02741 1546 1545 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02742 202 978 1545 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02743 200 978 1546 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02744 1579 1548 1547 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02745 1548 1547 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02746 201 978 1547 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02747 199 978 1548 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02748 1579 1550 1549 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02749 1550 1549 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02750 202 990 1549 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02751 200 990 1550 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02752 1579 1552 1551 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02753 1552 1551 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02754 201 990 1551 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02755 199 990 1552 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02756 1579 1554 1553 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02757 1554 1553 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02758 202 991 1553 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02759 200 991 1554 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02760 1579 1556 1555 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02761 1556 1555 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02762 201 991 1555 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02763 199 991 1556 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02764 1579 1558 1557 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02765 1558 1557 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02766 202 992 1557 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02767 200 992 1558 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02768 1579 1560 1559 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02769 1560 1559 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02770 201 992 1559 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02771 199 992 1560 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02772 1579 1562 1561 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02773 1562 1561 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02774 202 994 1561 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02775 200 994 1562 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02776 1579 1564 1563 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02777 1564 1563 1579 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02778 201 994 1563 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02779 199 994 1564 1579 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02780 199 1003 206 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02781 206 1004 200 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02782 201 1003 207 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02783 207 1004 202 1579 tn L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02784 1568 1036 1566 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02785 1574 1568 203 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02786 203 1573 1579 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02787 203 1566 1565 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02788 1579 1573 204 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02789 1567 207 204 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02790 204 206 1566 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02791 1568 207 205 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02792 205 1573 1579 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02793 205 206 1569 1579 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02794 1580 1036 207 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02795 207 1036 1580 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02796 1580 1036 206 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02797 206 1036 1580 1579 tn L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02798 1570 1576 207 1579 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_02799 206 1576 1571 1579 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_02800 207 1036 206 1579 tn L=1U W=22U AS=44P AD=44P PS=48U PD=48U 
Mtr_02801 1579 1582 1570 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_02802 1571 1572 1579 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_02803 1570 1582 1579 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_02804 1579 1572 1571 1579 tn L=1U W=27U AS=54P AD=54P PS=58U PD=58U 
Mtr_02805 1579 1582 1572 1579 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02806 1582 1575 1579 1579 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02807 1579 1575 1582 1579 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02808 1579 1576 1575 1579 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02809 1575 1574 1579 1579 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02810 1575 1573 1577 1579 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02811 209 208 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02812 1580 209 208 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02813 211 210 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02814 1580 211 210 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02815 213 212 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02816 1580 213 212 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02817 215 214 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02818 1580 215 214 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02819 217 216 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02820 1580 217 216 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02821 219 218 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02822 1580 219 218 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02823 221 220 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02824 1580 221 220 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02825 223 222 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02826 1580 223 222 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02827 225 224 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02828 1580 225 224 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02829 227 226 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02830 1580 227 226 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02831 229 228 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02832 1580 229 228 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02833 231 230 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02834 1580 231 230 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02835 233 232 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02836 1580 233 232 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02837 235 234 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02838 1580 235 234 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02839 237 236 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02840 1580 237 236 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02841 239 238 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02842 1580 239 238 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02843 241 240 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02844 1580 241 240 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02845 243 242 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02846 1580 243 242 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02847 245 244 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02848 1580 245 244 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02849 247 246 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02850 1580 247 246 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02851 249 248 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02852 1580 249 248 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02853 251 250 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02854 1580 251 250 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02855 253 252 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02856 1580 253 252 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02857 255 254 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02858 1580 255 254 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02859 257 256 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02860 1580 257 256 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02861 259 258 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02862 1580 259 258 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02863 261 260 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02864 1580 261 260 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02865 263 262 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02866 1580 263 262 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02867 265 264 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02868 1580 265 264 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02869 267 266 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02870 1580 267 266 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02871 269 268 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02872 1580 269 268 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02873 271 270 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02874 1580 271 270 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02875 273 272 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02876 1580 273 272 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02877 275 274 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02878 1580 275 274 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02879 277 276 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02880 1580 277 276 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02881 279 278 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02882 1580 279 278 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02883 281 280 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02884 1580 281 280 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02885 283 282 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02886 1580 283 282 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02887 285 284 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02888 1580 285 284 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02889 287 286 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02890 1580 287 286 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02891 289 288 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02892 1580 289 288 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02893 291 290 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02894 1580 291 290 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02895 293 292 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02896 1580 293 292 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02897 295 294 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02898 1580 295 294 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02899 297 296 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02900 1580 297 296 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02901 299 298 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02902 1580 299 298 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02903 301 300 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02904 1580 301 300 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02905 303 302 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02906 1580 303 302 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02907 305 304 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02908 1580 305 304 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02909 307 306 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02910 1580 307 306 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02911 309 308 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02912 1580 309 308 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02913 311 310 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02914 1580 311 310 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02915 313 312 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02916 1580 313 312 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02917 315 314 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02918 1580 315 314 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02919 317 316 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02920 1580 317 316 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02921 319 318 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02922 1580 319 318 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02923 321 320 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02924 1580 321 320 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02925 323 322 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02926 1580 323 322 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02927 325 324 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02928 1580 325 324 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02929 327 326 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02930 1580 327 326 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02931 329 328 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02932 1580 329 328 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02933 331 330 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02934 1580 331 330 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02935 333 332 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02936 1580 333 332 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02937 335 334 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02938 1580 335 334 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02939 337 336 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02940 1580 337 336 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02941 339 338 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02942 1580 339 338 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02943 341 340 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02944 1580 341 340 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02945 343 342 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02946 1580 343 342 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02947 345 344 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02948 1580 345 344 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02949 347 346 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02950 1580 347 346 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02951 349 348 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02952 1580 349 348 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02953 351 350 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02954 1580 351 350 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02955 353 352 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02956 1580 353 352 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02957 355 354 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02958 1580 355 354 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02959 357 356 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02960 1580 357 356 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02961 359 358 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02962 1580 359 358 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02963 361 360 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02964 1580 361 360 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02965 363 362 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02966 1580 363 362 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02967 365 364 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02968 1580 365 364 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02969 367 366 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02970 1580 367 366 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02971 369 368 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02972 1580 369 368 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02973 371 370 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02974 1580 371 370 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02975 373 372 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02976 1580 373 372 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02977 375 374 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02978 1580 375 374 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02979 377 376 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02980 1580 377 376 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02981 379 378 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02982 1580 379 378 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02983 381 380 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02984 1580 381 380 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02985 383 382 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02986 1580 383 382 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02987 385 384 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02988 1580 385 384 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02989 387 386 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02990 1580 387 386 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02991 389 388 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02992 1580 389 388 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02993 391 390 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02994 1580 391 390 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02995 393 392 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02996 1580 393 392 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02997 395 394 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02998 1580 395 394 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02999 397 396 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03000 1580 397 396 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03001 399 398 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03002 1580 399 398 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03003 401 400 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03004 1580 401 400 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03005 403 402 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03006 1580 403 402 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03007 405 404 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03008 1580 405 404 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03009 407 406 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03010 1580 407 406 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03011 409 408 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03012 1580 409 408 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03013 411 410 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03014 1580 411 410 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03015 413 412 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03016 1580 413 412 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03017 415 414 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03018 1580 415 414 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03019 417 416 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03020 1580 417 416 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03021 419 418 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03022 1580 419 418 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03023 421 420 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03024 1580 421 420 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03025 423 422 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03026 1580 423 422 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03027 425 424 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03028 1580 425 424 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03029 427 426 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03030 1580 427 426 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03031 429 428 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03032 1580 429 428 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03033 431 430 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03034 1580 431 430 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03035 433 432 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03036 1580 433 432 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03037 435 434 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03038 1580 435 434 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03039 437 436 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03040 1580 437 436 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03041 439 438 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03042 1580 439 438 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03043 441 440 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03044 1580 441 440 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03045 443 442 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03046 1580 443 442 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03047 445 444 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03048 1580 445 444 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03049 447 446 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03050 1580 447 446 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03051 449 448 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03052 1580 449 448 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03053 451 450 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03054 1580 451 450 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03055 453 452 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03056 1580 453 452 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03057 455 454 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03058 1580 455 454 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03059 457 456 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03060 1580 457 456 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03061 459 458 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03062 1580 459 458 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03063 461 460 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03064 1580 461 460 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03065 463 462 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03066 1580 463 462 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03067 472 464 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03068 1580 464 464 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03069 466 466 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03070 1580 466 465 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03071 467 468 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03072 1580 468 468 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03073 469 1585 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03074 1580 471 470 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03075 471 1585 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03076 1580 1585 471 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03077 1585 474 1580 1580 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03078 1580 474 1585 1580 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03079 1580 1029 474 1580 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_03080 474 472 1580 1580 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_03081 474 1032 473 1580 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_03082 476 475 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03083 1580 476 475 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03084 478 477 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03085 1580 478 477 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03086 480 479 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03087 1580 480 479 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03088 482 481 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03089 1580 482 481 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03090 484 483 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03091 1580 484 483 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03092 486 485 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03093 1580 486 485 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03094 488 487 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03095 1580 488 487 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03096 490 489 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03097 1580 490 489 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03098 492 491 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03099 1580 492 491 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03100 494 493 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03101 1580 494 493 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03102 496 495 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03103 1580 496 495 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03104 498 497 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03105 1580 498 497 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03106 500 499 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03107 1580 500 499 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03108 502 501 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03109 1580 502 501 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03110 504 503 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03111 1580 504 503 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03112 506 505 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03113 1580 506 505 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03114 508 507 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03115 1580 508 507 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03116 510 509 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03117 1580 510 509 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03118 512 511 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03119 1580 512 511 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03120 514 513 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03121 1580 514 513 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03122 516 515 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03123 1580 516 515 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03124 518 517 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03125 1580 518 517 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03126 520 519 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03127 1580 520 519 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03128 522 521 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03129 1580 522 521 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03130 524 523 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03131 1580 524 523 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03132 526 525 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03133 1580 526 525 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03134 528 527 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03135 1580 528 527 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03136 530 529 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03137 1580 530 529 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03138 532 531 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03139 1580 532 531 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03140 534 533 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03141 1580 534 533 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03142 536 535 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03143 1580 536 535 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03144 538 537 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03145 1580 538 537 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03146 540 539 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03147 1580 540 539 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03148 542 541 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03149 1580 542 541 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03150 544 543 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03151 1580 544 543 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03152 546 545 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03153 1580 546 545 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03154 548 547 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03155 1580 548 547 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03156 550 549 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03157 1580 550 549 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03158 552 551 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03159 1580 552 551 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03160 554 553 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03161 1580 554 553 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03162 556 555 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03163 1580 556 555 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03164 558 557 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03165 1580 558 557 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03166 560 559 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03167 1580 560 559 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03168 562 561 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03169 1580 562 561 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03170 564 563 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03171 1580 564 563 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03172 566 565 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03173 1580 566 565 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03174 568 567 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03175 1580 568 567 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03176 570 569 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03177 1580 570 569 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03178 572 571 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03179 1580 572 571 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03180 574 573 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03181 1580 574 573 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03182 576 575 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03183 1580 576 575 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03184 578 577 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03185 1580 578 577 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03186 580 579 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03187 1580 580 579 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03188 582 581 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03189 1580 582 581 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03190 584 583 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03191 1580 584 583 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03192 586 585 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03193 1580 586 585 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03194 588 587 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03195 1580 588 587 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03196 590 589 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03197 1580 590 589 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03198 592 591 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03199 1580 592 591 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03200 594 593 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03201 1580 594 593 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03202 596 595 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03203 1580 596 595 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03204 598 597 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03205 1580 598 597 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03206 600 599 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03207 1580 600 599 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03208 602 601 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03209 1580 602 601 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03210 604 603 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03211 1580 604 603 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03212 606 605 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03213 1580 606 605 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03214 608 607 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03215 1580 608 607 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03216 610 609 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03217 1580 610 609 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03218 612 611 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03219 1580 612 611 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03220 614 613 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03221 1580 614 613 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03222 616 615 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03223 1580 616 615 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03224 618 617 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03225 1580 618 617 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03226 620 619 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03227 1580 620 619 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03228 622 621 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03229 1580 622 621 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03230 624 623 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03231 1580 624 623 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03232 626 625 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03233 1580 626 625 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03234 628 627 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03235 1580 628 627 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03236 630 629 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03237 1580 630 629 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03238 632 631 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03239 1580 632 631 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03240 634 633 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03241 1580 634 633 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03242 636 635 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03243 1580 636 635 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03244 638 637 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03245 1580 638 637 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03246 640 639 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03247 1580 640 639 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03248 642 641 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03249 1580 642 641 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03250 644 643 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03251 1580 644 643 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03252 646 645 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03253 1580 646 645 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03254 648 647 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03255 1580 648 647 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03256 650 649 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03257 1580 650 649 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03258 652 651 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03259 1580 652 651 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03260 654 653 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03261 1580 654 653 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03262 656 655 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03263 1580 656 655 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03264 658 657 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03265 1580 658 657 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03266 660 659 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03267 1580 660 659 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03268 662 661 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03269 1580 662 661 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03270 664 663 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03271 1580 664 663 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03272 666 665 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03273 1580 666 665 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03274 668 667 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03275 1580 668 667 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03276 670 669 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03277 1580 670 669 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03278 672 671 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03279 1580 672 671 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03280 674 673 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03281 1580 674 673 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03282 676 675 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03283 1580 676 675 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03284 678 677 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03285 1580 678 677 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03286 680 679 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03287 1580 680 679 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03288 682 681 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03289 1580 682 681 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03290 684 683 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03291 1580 684 683 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03292 686 685 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03293 1580 686 685 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03294 688 687 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03295 1580 688 687 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03296 690 689 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03297 1580 690 689 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03298 692 691 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03299 1580 692 691 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03300 694 693 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03301 1580 694 693 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03302 696 695 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03303 1580 696 695 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03304 698 697 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03305 1580 698 697 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03306 700 699 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03307 1580 700 699 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03308 702 701 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03309 1580 702 701 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03310 704 703 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03311 1580 704 703 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03312 706 705 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03313 1580 706 705 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03314 708 707 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03315 1580 708 707 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03316 710 709 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03317 1580 710 709 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03318 712 711 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03319 1580 712 711 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03320 714 713 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03321 1580 714 713 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03322 716 715 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03323 1580 716 715 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03324 718 717 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03325 1580 718 717 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03326 720 719 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03327 1580 720 719 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03328 722 721 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03329 1580 722 721 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03330 724 723 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03331 1580 724 723 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03332 726 725 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03333 1580 726 725 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03334 728 727 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03335 1580 728 727 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03336 730 729 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03337 1580 730 729 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03338 739 731 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03339 1580 731 731 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03340 733 733 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03341 1580 733 732 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03342 734 735 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03343 1580 735 735 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03344 736 1584 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03345 1580 738 737 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03346 738 1584 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03347 1580 1584 738 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03348 1584 741 1580 1580 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03349 1580 741 1584 1580 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03350 1580 1029 741 1580 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_03351 741 739 1580 1580 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_03352 741 1032 740 1580 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_03353 742 744 1580 1580 tp L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_03354 1580 744 742 1580 tp L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_03355 742 744 1580 1580 tp L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_03356 1580 744 742 1580 tp L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_03357 743 746 1580 1580 tp L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_03358 1580 746 743 1580 tp L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_03359 743 746 1580 1580 tp L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_03360 1580 746 743 1580 tp L=1U W=62U AS=124P AD=124P PS=128U PD=128U 
Mtr_03361 745 1040 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03362 1580 745 744 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03363 744 1041 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03364 1580 745 746 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03365 746 1041 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03366 749 1006 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03367 1580 1009 749 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03368 1580 1015 747 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03369 747 1012 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03370 748 747 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03371 753 749 748 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03372 1580 762 750 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03373 752 758 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03374 751 756 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03375 754 760 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03376 750 762 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03377 1580 756 751 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03378 762 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03379 1580 1026 762 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03380 762 753 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03381 756 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03382 1580 1022 756 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03383 756 753 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03384 1580 758 752 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03385 1580 1040 758 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03386 758 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03387 1580 753 758 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03388 760 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03389 1580 753 760 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03390 1580 1040 760 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03391 1580 760 754 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03392 755 756 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03393 1580 756 755 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03394 757 758 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03395 1580 758 757 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03396 759 760 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03397 1580 760 759 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03398 761 762 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03399 1580 762 761 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03400 765 1005 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03401 1580 1009 765 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03402 1580 1015 763 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03403 763 1012 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03404 764 763 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03405 769 765 764 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03406 1580 778 766 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03407 768 774 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03408 767 772 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03409 770 776 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03410 766 778 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03411 1580 772 767 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03412 778 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03413 1580 1026 778 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03414 778 769 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03415 772 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03416 1580 1022 772 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03417 772 769 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03418 1580 774 768 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03419 1580 1040 774 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03420 774 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03421 1580 769 774 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03422 776 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03423 1580 769 776 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03424 1580 1040 776 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03425 1580 776 770 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03426 771 772 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03427 1580 772 771 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03428 773 774 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03429 1580 774 773 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03430 775 776 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03431 1580 776 775 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03432 777 778 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03433 1580 778 777 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03434 781 1006 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03435 1580 1008 781 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03436 1580 1015 779 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03437 779 1012 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03438 780 779 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03439 785 781 780 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03440 1580 794 782 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03441 784 790 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03442 783 788 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03443 786 792 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03444 782 794 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03445 1580 788 783 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03446 794 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03447 1580 1026 794 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03448 794 785 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03449 788 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03450 1580 1022 788 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03451 788 785 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03452 1580 790 784 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03453 1580 1040 790 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03454 790 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03455 1580 785 790 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03456 792 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03457 1580 785 792 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03458 1580 1040 792 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03459 1580 792 786 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03460 787 788 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03461 1580 788 787 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03462 789 790 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03463 1580 790 789 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03464 791 792 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03465 1580 792 791 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03466 793 794 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03467 1580 794 793 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03468 797 1005 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03469 1580 1008 797 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03470 1580 1015 795 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03471 795 1012 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03472 796 795 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03473 801 797 796 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03474 1580 810 798 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03475 800 806 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03476 799 804 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03477 802 808 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03478 798 810 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03479 1580 804 799 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03480 810 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03481 1580 1026 810 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03482 810 801 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03483 804 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03484 1580 1022 804 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03485 804 801 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03486 1580 806 800 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03487 1580 1040 806 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03488 806 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03489 1580 801 806 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03490 808 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03491 1580 801 808 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03492 1580 1040 808 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03493 1580 808 802 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03494 803 804 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03495 1580 804 803 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03496 805 806 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03497 1580 806 805 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03498 807 808 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03499 1580 808 807 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03500 809 810 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03501 1580 810 809 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03502 813 1006 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03503 1580 1009 813 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03504 1580 1015 811 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03505 811 1011 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03506 812 811 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03507 817 813 812 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03508 1580 826 814 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03509 816 822 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03510 815 820 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03511 818 824 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03512 814 826 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03513 1580 820 815 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03514 826 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03515 1580 1026 826 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03516 826 817 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03517 820 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03518 1580 1022 820 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03519 820 817 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03520 1580 822 816 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03521 1580 1040 822 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03522 822 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03523 1580 817 822 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03524 824 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03525 1580 817 824 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03526 1580 1040 824 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03527 1580 824 818 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03528 819 820 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03529 1580 820 819 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03530 821 822 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03531 1580 822 821 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03532 823 824 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03533 1580 824 823 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03534 825 826 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03535 1580 826 825 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03536 829 1005 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03537 1580 1009 829 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03538 1580 1015 827 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03539 827 1011 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03540 828 827 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03541 833 829 828 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03542 1580 842 830 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03543 832 838 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03544 831 836 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03545 834 840 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03546 830 842 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03547 1580 836 831 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03548 842 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03549 1580 1026 842 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03550 842 833 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03551 836 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03552 1580 1022 836 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03553 836 833 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03554 1580 838 832 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03555 1580 1040 838 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03556 838 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03557 1580 833 838 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03558 840 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03559 1580 833 840 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03560 1580 1040 840 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03561 1580 840 834 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03562 835 836 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03563 1580 836 835 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03564 837 838 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03565 1580 838 837 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03566 839 840 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03567 1580 840 839 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03568 841 842 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03569 1580 842 841 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03570 845 1006 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03571 1580 1008 845 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03572 1580 1015 843 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03573 843 1011 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03574 844 843 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03575 849 845 844 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03576 1580 858 846 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03577 848 854 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03578 847 852 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03579 850 856 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03580 846 858 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03581 1580 852 847 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03582 858 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03583 1580 1026 858 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03584 858 849 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03585 852 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03586 1580 1022 852 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03587 852 849 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03588 1580 854 848 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03589 1580 1040 854 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03590 854 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03591 1580 849 854 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03592 856 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03593 1580 849 856 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03594 1580 1040 856 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03595 1580 856 850 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03596 851 852 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03597 1580 852 851 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03598 853 854 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03599 1580 854 853 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03600 855 856 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03601 1580 856 855 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03602 857 858 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03603 1580 858 857 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03604 861 1005 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03605 1580 1008 861 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03606 1580 1015 859 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03607 859 1011 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03608 860 859 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03609 865 861 860 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03610 1580 874 862 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03611 864 870 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03612 863 868 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03613 866 872 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03614 862 874 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03615 1580 868 863 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03616 874 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03617 1580 1026 874 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03618 874 865 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03619 868 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03620 1580 1022 868 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03621 868 865 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03622 1580 870 864 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03623 1580 1040 870 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03624 870 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03625 1580 865 870 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03626 872 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03627 1580 865 872 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03628 1580 1040 872 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03629 1580 872 866 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03630 867 868 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03631 1580 868 867 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03632 869 870 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03633 1580 870 869 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03634 871 872 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03635 1580 872 871 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03636 873 874 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03637 1580 874 873 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03638 877 1006 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03639 1580 1009 877 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03640 1580 1014 875 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03641 875 1012 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03642 876 875 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03643 881 877 876 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03644 1580 890 878 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03645 880 886 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03646 879 884 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03647 882 888 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03648 878 890 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03649 1580 884 879 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03650 890 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03651 1580 1026 890 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03652 890 881 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03653 884 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03654 1580 1022 884 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03655 884 881 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03656 1580 886 880 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03657 1580 1040 886 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03658 886 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03659 1580 881 886 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03660 888 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03661 1580 881 888 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03662 1580 1040 888 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03663 1580 888 882 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03664 883 884 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03665 1580 884 883 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03666 885 886 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03667 1580 886 885 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03668 887 888 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03669 1580 888 887 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03670 889 890 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03671 1580 890 889 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03672 893 1005 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03673 1580 1009 893 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03674 1580 1014 891 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03675 891 1012 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03676 892 891 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03677 897 893 892 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03678 1580 906 894 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03679 896 902 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03680 895 900 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03681 898 904 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03682 894 906 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03683 1580 900 895 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03684 906 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03685 1580 1026 906 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03686 906 897 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03687 900 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03688 1580 1022 900 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03689 900 897 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03690 1580 902 896 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03691 1580 1040 902 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03692 902 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03693 1580 897 902 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03694 904 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03695 1580 897 904 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03696 1580 1040 904 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03697 1580 904 898 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03698 899 900 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03699 1580 900 899 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03700 901 902 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03701 1580 902 901 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03702 903 904 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03703 1580 904 903 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03704 905 906 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03705 1580 906 905 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03706 909 1006 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03707 1580 1008 909 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03708 1580 1014 907 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03709 907 1012 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03710 908 907 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03711 913 909 908 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03712 1580 922 910 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03713 912 918 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03714 911 916 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03715 914 920 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03716 910 922 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03717 1580 916 911 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03718 922 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03719 1580 1026 922 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03720 922 913 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03721 916 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03722 1580 1022 916 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03723 916 913 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03724 1580 918 912 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03725 1580 1040 918 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03726 918 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03727 1580 913 918 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03728 920 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03729 1580 913 920 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03730 1580 1040 920 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03731 1580 920 914 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03732 915 916 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03733 1580 916 915 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03734 917 918 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03735 1580 918 917 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03736 919 920 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03737 1580 920 919 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03738 921 922 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03739 1580 922 921 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03740 925 1005 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03741 1580 1008 925 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03742 1580 1014 923 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03743 923 1012 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03744 924 923 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03745 929 925 924 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03746 1580 938 926 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03747 928 934 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03748 927 932 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03749 930 936 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03750 926 938 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03751 1580 932 927 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03752 938 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03753 1580 1026 938 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03754 938 929 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03755 932 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03756 1580 1022 932 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03757 932 929 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03758 1580 934 928 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03759 1580 1040 934 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03760 934 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03761 1580 929 934 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03762 936 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03763 1580 929 936 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03764 1580 1040 936 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03765 1580 936 930 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03766 931 932 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03767 1580 932 931 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03768 933 934 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03769 1580 934 933 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03770 935 936 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03771 1580 936 935 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03772 937 938 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03773 1580 938 937 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03774 941 1006 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03775 1580 1009 941 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03776 1580 1014 939 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03777 939 1011 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03778 940 939 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03779 945 941 940 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03780 1580 954 942 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03781 944 950 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03782 943 948 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03783 946 952 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03784 942 954 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03785 1580 948 943 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03786 954 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03787 1580 1026 954 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03788 954 945 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03789 948 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03790 1580 1022 948 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03791 948 945 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03792 1580 950 944 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03793 1580 1040 950 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03794 950 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03795 1580 945 950 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03796 952 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03797 1580 945 952 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03798 1580 1040 952 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03799 1580 952 946 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03800 947 948 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03801 1580 948 947 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03802 949 950 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03803 1580 950 949 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03804 951 952 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03805 1580 952 951 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03806 953 954 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03807 1580 954 953 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03808 957 1005 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03809 1580 1009 957 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03810 1580 1014 955 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03811 955 1011 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03812 956 955 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03813 961 957 956 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03814 1580 970 958 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03815 960 966 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03816 959 964 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03817 962 968 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03818 958 970 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03819 1580 964 959 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03820 970 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03821 1580 1026 970 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03822 970 961 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03823 964 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03824 1580 1022 964 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03825 964 961 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03826 1580 966 960 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03827 1580 1040 966 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03828 966 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03829 1580 961 966 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03830 968 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03831 1580 961 968 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03832 1580 1040 968 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03833 1580 968 962 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03834 963 964 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03835 1580 964 963 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03836 965 966 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03837 1580 966 965 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03838 967 968 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03839 1580 968 967 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03840 969 970 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03841 1580 970 969 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03842 973 1006 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03843 1580 1008 973 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03844 1580 1014 971 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03845 971 1011 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03846 972 971 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03847 977 973 972 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03848 1580 986 974 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03849 976 982 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03850 975 980 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03851 978 984 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03852 974 986 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03853 1580 980 975 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03854 986 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03855 1580 1026 986 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03856 986 977 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03857 980 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03858 1580 1022 980 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03859 980 977 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03860 1580 982 976 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03861 1580 1040 982 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03862 982 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03863 1580 977 982 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03864 984 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03865 1580 977 984 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03866 1580 1040 984 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03867 1580 984 978 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03868 979 980 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03869 1580 980 979 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03870 981 982 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03871 1580 982 981 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03872 983 984 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03873 1580 984 983 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03874 985 986 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03875 1580 986 985 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03876 989 1005 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03877 1580 1008 989 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03878 1580 1014 987 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03879 987 1011 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03880 988 987 1580 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03881 993 989 988 1580 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_03882 1580 1002 990 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03883 992 998 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03884 991 996 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03885 994 1000 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03886 990 1002 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03887 1580 996 991 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03888 1002 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03889 1580 1026 1002 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03890 1002 993 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03891 996 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03892 1580 1022 996 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03893 996 993 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03894 1580 998 992 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03895 1580 1040 998 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03896 998 1023 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03897 1580 993 998 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03898 1000 1019 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03899 1580 993 1000 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03900 1580 1040 1000 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03901 1580 1000 994 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03902 995 996 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03903 1580 996 995 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03904 997 998 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03905 1580 998 997 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03906 999 1000 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03907 1580 1000 999 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03908 1001 1002 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03909 1580 1002 1001 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03910 1580 1027 1003 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03911 1004 1028 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03912 1005 1590 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03913 1580 1007 1006 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03914 1580 1590 1007 1580 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03915 1008 1589 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03916 1580 1010 1009 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03917 1580 1589 1010 1580 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03918 1011 1588 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03919 1580 1013 1012 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03920 1580 1588 1013 1580 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03921 1014 1587 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03922 1580 1016 1015 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03923 1580 1587 1016 1580 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03924 1580 1592 1017 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03925 1018 1591 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03926 1580 1592 1025 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03927 1025 1591 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03928 1580 1592 1024 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03929 1020 1018 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03930 1580 1017 1020 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03931 1021 1591 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03932 1580 1017 1021 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03933 1024 1018 1580 1580 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03934 1580 1020 1019 1580 tp L=1U W=38U AS=76P AD=76P PS=80U PD=80U 
Mtr_03935 1022 1021 1580 1580 tp L=1U W=38U AS=76P AD=76P PS=80U PD=80U 
Mtr_03936 1580 1024 1023 1580 tp L=1U W=38U AS=76P AD=76P PS=80U PD=80U 
Mtr_03937 1026 1025 1580 1580 tp L=1U W=38U AS=76P AD=76P PS=80U PD=80U 
Mtr_03938 1027 1028 1580 1580 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_03939 1580 1593 1028 1580 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_03940 1029 1030 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03941 1030 1033 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03942 1580 1030 1029 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03943 1573 1031 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03944 1031 1034 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03945 1580 1031 1573 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03946 1032 1033 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03947 1033 1578 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03948 1580 1040 1033 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03949 1580 1033 1032 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03950 1576 1034 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03951 1034 1578 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03952 1580 1040 1034 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03953 1580 1034 1576 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03954 1580 1035 1036 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03955 1580 1041 1035 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03956 1035 1039 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03957 1036 1035 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03958 1580 1037 1038 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03959 1580 1041 1037 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03960 1037 1039 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03961 1038 1037 1580 1580 tp L=1U W=39U AS=78P AD=78P PS=82U PD=82U 
Mtr_03962 1039 1040 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_03963 1580 1041 1040 1580 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_03964 1040 1041 1580 1580 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_03965 1580 1041 1040 1580 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_03966 1040 1041 1580 1580 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_03967 1041 1586 1580 1580 tp L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_03968 1580 1581 1041 1580 tp L=1U W=17U AS=34P AD=34P PS=38U PD=38U 
Mtr_03969 1043 1042 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03970 1580 1043 1042 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03971 1045 1044 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03972 1580 1045 1044 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03973 1047 1046 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03974 1580 1047 1046 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03975 1049 1048 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03976 1580 1049 1048 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03977 1051 1050 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03978 1580 1051 1050 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03979 1053 1052 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03980 1580 1053 1052 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03981 1055 1054 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03982 1580 1055 1054 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03983 1057 1056 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03984 1580 1057 1056 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03985 1059 1058 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03986 1580 1059 1058 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03987 1061 1060 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03988 1580 1061 1060 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03989 1063 1062 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03990 1580 1063 1062 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03991 1065 1064 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03992 1580 1065 1064 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03993 1067 1066 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03994 1580 1067 1066 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03995 1069 1068 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03996 1580 1069 1068 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03997 1071 1070 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03998 1580 1071 1070 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_03999 1073 1072 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04000 1580 1073 1072 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04001 1075 1074 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04002 1580 1075 1074 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04003 1077 1076 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04004 1580 1077 1076 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04005 1079 1078 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04006 1580 1079 1078 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04007 1081 1080 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04008 1580 1081 1080 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04009 1083 1082 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04010 1580 1083 1082 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04011 1085 1084 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04012 1580 1085 1084 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04013 1087 1086 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04014 1580 1087 1086 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04015 1089 1088 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04016 1580 1089 1088 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04017 1091 1090 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04018 1580 1091 1090 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04019 1093 1092 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04020 1580 1093 1092 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04021 1095 1094 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04022 1580 1095 1094 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04023 1097 1096 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04024 1580 1097 1096 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04025 1099 1098 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04026 1580 1099 1098 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04027 1101 1100 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04028 1580 1101 1100 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04029 1103 1102 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04030 1580 1103 1102 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04031 1105 1104 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04032 1580 1105 1104 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04033 1107 1106 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04034 1580 1107 1106 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04035 1109 1108 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04036 1580 1109 1108 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04037 1111 1110 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04038 1580 1111 1110 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04039 1113 1112 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04040 1580 1113 1112 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04041 1115 1114 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04042 1580 1115 1114 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04043 1117 1116 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04044 1580 1117 1116 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04045 1119 1118 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04046 1580 1119 1118 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04047 1121 1120 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04048 1580 1121 1120 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04049 1123 1122 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04050 1580 1123 1122 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04051 1125 1124 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04052 1580 1125 1124 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04053 1127 1126 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04054 1580 1127 1126 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04055 1129 1128 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04056 1580 1129 1128 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04057 1131 1130 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04058 1580 1131 1130 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04059 1133 1132 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04060 1580 1133 1132 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04061 1135 1134 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04062 1580 1135 1134 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04063 1137 1136 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04064 1580 1137 1136 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04065 1139 1138 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04066 1580 1139 1138 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04067 1141 1140 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04068 1580 1141 1140 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04069 1143 1142 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04070 1580 1143 1142 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04071 1145 1144 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04072 1580 1145 1144 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04073 1147 1146 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04074 1580 1147 1146 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04075 1149 1148 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04076 1580 1149 1148 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04077 1151 1150 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04078 1580 1151 1150 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04079 1153 1152 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04080 1580 1153 1152 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04081 1155 1154 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04082 1580 1155 1154 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04083 1157 1156 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04084 1580 1157 1156 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04085 1159 1158 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04086 1580 1159 1158 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04087 1161 1160 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04088 1580 1161 1160 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04089 1163 1162 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04090 1580 1163 1162 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04091 1165 1164 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04092 1580 1165 1164 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04093 1167 1166 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04094 1580 1167 1166 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04095 1169 1168 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04096 1580 1169 1168 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04097 1171 1170 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04098 1580 1171 1170 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04099 1173 1172 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04100 1580 1173 1172 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04101 1175 1174 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04102 1580 1175 1174 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04103 1177 1176 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04104 1580 1177 1176 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04105 1179 1178 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04106 1580 1179 1178 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04107 1181 1180 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04108 1580 1181 1180 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04109 1183 1182 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04110 1580 1183 1182 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04111 1185 1184 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04112 1580 1185 1184 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04113 1187 1186 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04114 1580 1187 1186 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04115 1189 1188 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04116 1580 1189 1188 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04117 1191 1190 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04118 1580 1191 1190 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04119 1193 1192 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04120 1580 1193 1192 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04121 1195 1194 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04122 1580 1195 1194 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04123 1197 1196 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04124 1580 1197 1196 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04125 1199 1198 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04126 1580 1199 1198 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04127 1201 1200 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04128 1580 1201 1200 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04129 1203 1202 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04130 1580 1203 1202 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04131 1205 1204 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04132 1580 1205 1204 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04133 1207 1206 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04134 1580 1207 1206 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04135 1209 1208 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04136 1580 1209 1208 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04137 1211 1210 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04138 1580 1211 1210 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04139 1213 1212 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04140 1580 1213 1212 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04141 1215 1214 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04142 1580 1215 1214 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04143 1217 1216 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04144 1580 1217 1216 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04145 1219 1218 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04146 1580 1219 1218 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04147 1221 1220 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04148 1580 1221 1220 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04149 1223 1222 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04150 1580 1223 1222 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04151 1225 1224 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04152 1580 1225 1224 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04153 1227 1226 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04154 1580 1227 1226 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04155 1229 1228 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04156 1580 1229 1228 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04157 1231 1230 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04158 1580 1231 1230 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04159 1233 1232 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04160 1580 1233 1232 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04161 1235 1234 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04162 1580 1235 1234 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04163 1237 1236 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04164 1580 1237 1236 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04165 1239 1238 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04166 1580 1239 1238 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04167 1241 1240 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04168 1580 1241 1240 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04169 1243 1242 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04170 1580 1243 1242 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04171 1245 1244 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04172 1580 1245 1244 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04173 1247 1246 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04174 1580 1247 1246 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04175 1249 1248 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04176 1580 1249 1248 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04177 1251 1250 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04178 1580 1251 1250 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04179 1253 1252 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04180 1580 1253 1252 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04181 1255 1254 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04182 1580 1255 1254 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04183 1257 1256 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04184 1580 1257 1256 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04185 1259 1258 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04186 1580 1259 1258 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04187 1261 1260 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04188 1580 1261 1260 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04189 1263 1262 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04190 1580 1263 1262 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04191 1265 1264 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04192 1580 1265 1264 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04193 1267 1266 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04194 1580 1267 1266 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04195 1269 1268 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04196 1580 1269 1268 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04197 1271 1270 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04198 1580 1271 1270 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04199 1273 1272 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04200 1580 1273 1272 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04201 1275 1274 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04202 1580 1275 1274 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04203 1277 1276 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04204 1580 1277 1276 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04205 1279 1278 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04206 1580 1279 1278 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04207 1281 1280 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04208 1580 1281 1280 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04209 1283 1282 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04210 1580 1283 1282 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04211 1285 1284 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04212 1580 1285 1284 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04213 1287 1286 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04214 1580 1287 1286 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04215 1289 1288 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04216 1580 1289 1288 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04217 1291 1290 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04218 1580 1291 1290 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04219 1293 1292 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04220 1580 1293 1292 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04221 1295 1294 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04222 1580 1295 1294 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04223 1297 1296 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04224 1580 1297 1296 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04225 1306 1298 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04226 1580 1298 1298 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04227 1300 1300 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04228 1580 1300 1299 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04229 1301 1302 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04230 1580 1302 1302 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04231 1303 1583 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04232 1580 1305 1304 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04233 1305 1583 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04234 1580 1583 1305 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04235 1583 1308 1580 1580 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04236 1580 1308 1583 1580 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04237 1580 1573 1308 1580 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_04238 1308 1306 1580 1580 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_04239 1308 1576 1307 1580 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_04240 1310 1309 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04241 1580 1310 1309 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04242 1312 1311 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04243 1580 1312 1311 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04244 1314 1313 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04245 1580 1314 1313 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04246 1316 1315 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04247 1580 1316 1315 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04248 1318 1317 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04249 1580 1318 1317 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04250 1320 1319 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04251 1580 1320 1319 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04252 1322 1321 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04253 1580 1322 1321 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04254 1324 1323 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04255 1580 1324 1323 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04256 1326 1325 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04257 1580 1326 1325 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04258 1328 1327 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04259 1580 1328 1327 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04260 1330 1329 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04261 1580 1330 1329 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04262 1332 1331 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04263 1580 1332 1331 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04264 1334 1333 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04265 1580 1334 1333 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04266 1336 1335 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04267 1580 1336 1335 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04268 1338 1337 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04269 1580 1338 1337 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04270 1340 1339 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04271 1580 1340 1339 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04272 1342 1341 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04273 1580 1342 1341 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04274 1344 1343 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04275 1580 1344 1343 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04276 1346 1345 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04277 1580 1346 1345 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04278 1348 1347 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04279 1580 1348 1347 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04280 1350 1349 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04281 1580 1350 1349 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04282 1352 1351 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04283 1580 1352 1351 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04284 1354 1353 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04285 1580 1354 1353 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04286 1356 1355 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04287 1580 1356 1355 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04288 1358 1357 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04289 1580 1358 1357 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04290 1360 1359 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04291 1580 1360 1359 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04292 1362 1361 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04293 1580 1362 1361 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04294 1364 1363 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04295 1580 1364 1363 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04296 1366 1365 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04297 1580 1366 1365 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04298 1368 1367 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04299 1580 1368 1367 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04300 1370 1369 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04301 1580 1370 1369 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04302 1372 1371 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04303 1580 1372 1371 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04304 1374 1373 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04305 1580 1374 1373 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04306 1376 1375 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04307 1580 1376 1375 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04308 1378 1377 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04309 1580 1378 1377 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04310 1380 1379 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04311 1580 1380 1379 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04312 1382 1381 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04313 1580 1382 1381 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04314 1384 1383 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04315 1580 1384 1383 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04316 1386 1385 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04317 1580 1386 1385 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04318 1388 1387 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04319 1580 1388 1387 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04320 1390 1389 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04321 1580 1390 1389 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04322 1392 1391 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04323 1580 1392 1391 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04324 1394 1393 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04325 1580 1394 1393 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04326 1396 1395 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04327 1580 1396 1395 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04328 1398 1397 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04329 1580 1398 1397 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04330 1400 1399 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04331 1580 1400 1399 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04332 1402 1401 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04333 1580 1402 1401 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04334 1404 1403 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04335 1580 1404 1403 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04336 1406 1405 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04337 1580 1406 1405 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04338 1408 1407 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04339 1580 1408 1407 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04340 1410 1409 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04341 1580 1410 1409 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04342 1412 1411 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04343 1580 1412 1411 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04344 1414 1413 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04345 1580 1414 1413 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04346 1416 1415 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04347 1580 1416 1415 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04348 1418 1417 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04349 1580 1418 1417 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04350 1420 1419 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04351 1580 1420 1419 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04352 1422 1421 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04353 1580 1422 1421 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04354 1424 1423 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04355 1580 1424 1423 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04356 1426 1425 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04357 1580 1426 1425 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04358 1428 1427 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04359 1580 1428 1427 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04360 1430 1429 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04361 1580 1430 1429 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04362 1432 1431 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04363 1580 1432 1431 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04364 1434 1433 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04365 1580 1434 1433 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04366 1436 1435 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04367 1580 1436 1435 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04368 1438 1437 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04369 1580 1438 1437 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04370 1440 1439 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04371 1580 1440 1439 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04372 1442 1441 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04373 1580 1442 1441 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04374 1444 1443 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04375 1580 1444 1443 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04376 1446 1445 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04377 1580 1446 1445 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04378 1448 1447 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04379 1580 1448 1447 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04380 1450 1449 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04381 1580 1450 1449 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04382 1452 1451 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04383 1580 1452 1451 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04384 1454 1453 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04385 1580 1454 1453 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04386 1456 1455 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04387 1580 1456 1455 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04388 1458 1457 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04389 1580 1458 1457 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04390 1460 1459 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04391 1580 1460 1459 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04392 1462 1461 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04393 1580 1462 1461 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04394 1464 1463 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04395 1580 1464 1463 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04396 1466 1465 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04397 1580 1466 1465 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04398 1468 1467 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04399 1580 1468 1467 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04400 1470 1469 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04401 1580 1470 1469 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04402 1472 1471 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04403 1580 1472 1471 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04404 1474 1473 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04405 1580 1474 1473 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04406 1476 1475 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04407 1580 1476 1475 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04408 1478 1477 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04409 1580 1478 1477 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04410 1480 1479 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04411 1580 1480 1479 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04412 1482 1481 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04413 1580 1482 1481 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04414 1484 1483 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04415 1580 1484 1483 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04416 1486 1485 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04417 1580 1486 1485 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04418 1488 1487 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04419 1580 1488 1487 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04420 1490 1489 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04421 1580 1490 1489 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04422 1492 1491 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04423 1580 1492 1491 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04424 1494 1493 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04425 1580 1494 1493 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04426 1496 1495 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04427 1580 1496 1495 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04428 1498 1497 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04429 1580 1498 1497 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04430 1500 1499 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04431 1580 1500 1499 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04432 1502 1501 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04433 1580 1502 1501 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04434 1504 1503 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04435 1580 1504 1503 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04436 1506 1505 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04437 1580 1506 1505 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04438 1508 1507 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04439 1580 1508 1507 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04440 1510 1509 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04441 1580 1510 1509 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04442 1512 1511 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04443 1580 1512 1511 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04444 1514 1513 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04445 1580 1514 1513 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04446 1516 1515 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04447 1580 1516 1515 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04448 1518 1517 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04449 1580 1518 1517 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04450 1520 1519 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04451 1580 1520 1519 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04452 1522 1521 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04453 1580 1522 1521 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04454 1524 1523 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04455 1580 1524 1523 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04456 1526 1525 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04457 1580 1526 1525 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04458 1528 1527 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04459 1580 1528 1527 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04460 1530 1529 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04461 1580 1530 1529 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04462 1532 1531 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04463 1580 1532 1531 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04464 1534 1533 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04465 1580 1534 1533 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04466 1536 1535 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04467 1580 1536 1535 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04468 1538 1537 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04469 1580 1538 1537 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04470 1540 1539 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04471 1580 1540 1539 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04472 1542 1541 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04473 1580 1542 1541 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04474 1544 1543 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04475 1580 1544 1543 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04476 1546 1545 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04477 1580 1546 1545 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04478 1548 1547 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04479 1580 1548 1547 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04480 1550 1549 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04481 1580 1550 1549 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04482 1552 1551 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04483 1580 1552 1551 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04484 1554 1553 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04485 1580 1554 1553 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04486 1556 1555 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04487 1580 1556 1555 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04488 1558 1557 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04489 1580 1558 1557 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04490 1560 1559 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04491 1580 1560 1559 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04492 1562 1561 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04493 1580 1562 1561 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04494 1564 1563 1580 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04495 1580 1564 1563 1580 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_04496 1574 1565 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04497 1580 1565 1565 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04498 1567 1567 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04499 1580 1567 1566 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04500 1568 1569 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04501 1580 1569 1569 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04502 1570 1582 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04503 1580 1572 1571 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04504 1572 1582 1580 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04505 1580 1582 1572 1580 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_04506 1582 1577 1580 1580 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04507 1580 1577 1582 1580 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04508 1580 1573 1577 1580 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_04509 1577 1574 1580 1580 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_04510 1577 1576 1575 1580 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
.ends ram4x128

