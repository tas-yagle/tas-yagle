* Spice description of r256x8_5
* Spice driver version 700
* Date ( dd/mm/yyyy hh:mm:ss ): 20/09/2002 at 17:50:04

* INTERF adr[0] adr[1] adr[2] adr[3] adr[4] adr[5] adr[6] adr[7] ck[0] ck[1] 
* INTERF f[0] f[1] f[2] f[3] f[4] f[5] f[6] f[7] vdd vss 


.subckt r256x8_5 308 302 303 304 296 297 298 294 210 1 326 323 321 319 
+ 317 315 313 311 324 327 
* NET 1 = ck[1] 
* NET 5 = rl/7.w1 
* NET 6 = rbl4/1/2.e0 
* NET 7 = rck.ckp 
* NET 13 = rl/7.e1 
* NET 14 = rl/7.tr_p 
* NET 15 = rl/7.w2 
* NET 16 = rl/7.w3 
* NET 17 = rl/7.w4 
* NET 18 = rbl4/1/2.e1 
* NET 19 = rbl4/1/2.e2 
* NET 20 = rbl4/1/2.e3 
* NET 26 = rl/6.e1 
* NET 27 = rl/6.tr_p 
* NET 28 = rl/6.w1 
* NET 29 = rl/6.w2 
* NET 30 = rl/6.w3 
* NET 31 = rl/6.w4 
* NET 32 = rbl4/1/2.e7 
* NET 33 = rbl4/1/2.e6 
* NET 34 = umf.e31 
* NET 35 = rbl4/1/2.e5 
* NET 40 = rl/5.w1 
* NET 41 = rl/5.w2 
* NET 42 = rl/5.w3 
* NET 43 = rbl4/1/2.e10 
* NET 44 = rbl4/1/2.e8 
* NET 45 = rbl4/1/2.e9 
* NET 50 = rl/5.e1 
* NET 51 = rl/5.tr_p 
* NET 52 = rl/5.w4 
* NET 53 = rl/4.w1 
* NET 54 = rl/4.w2 
* NET 55 = rbl4/1/2.e11 
* NET 56 = rbl4/1/2.e14 
* NET 57 = rbl4/1/2.e13 
* NET 58 = rbl4/1/2.e12 
* NET 63 = rl/4.e1 
* NET 64 = rl/4.tr_p 
* NET 65 = rl/4.w3 
* NET 66 = rl/4.w4 
* NET 67 = rl/3.w1 
* NET 68 = rl/3.w2 
* NET 69 = umf.e0 
* NET 70 = rbl4/1/2.e15 
* NET 71 = umf.e1 
* NET 77 = rl/3.e1 
* NET 78 = rl/3.tr_p 
* NET 79 = rl/3.w3 
* NET 80 = rl/3.w4 
* NET 81 = rl/2.w1 
* NET 82 = rl/2.w2 
* NET 83 = umf.e2 
* NET 84 = umf.e5 
* NET 85 = umf.e4 
* NET 86 = umf.e3 
* NET 92 = rl/2.e1 
* NET 93 = rl/2.tr_p 
* NET 94 = rl/2.w3 
* NET 95 = rl/2.w4 
* NET 96 = rl/1.w1 
* NET 97 = umf.e8 
* NET 98 = umf.e7 
* NET 99 = umf.e6 
* NET 103 = rl/1.e1 
* NET 104 = rl/1.tr_p 
* NET 105 = rl/1.w2 
* NET 106 = rl/1.w3 
* NET 107 = rl/1.w4 
* NET 108 = rl/0.w1 
* NET 109 = umf.e9 
* NET 110 = umf.e12 
* NET 111 = umf.e11 
* NET 112 = umf.e10 
* NET 115 = rck.ck_02 
* NET 119 = rl/0.e1 
* NET 120 = rl/0.tr_p 
* NET 121 = rck.ck_03 
* NET 122 = rl/0.w2 
* NET 123 = rl/0.w3 
* NET 124 = rl/0.w4 
* NET 125 = umf.e14 
* NET 126 = umf.e13 
* NET 127 = umf.e15 
* NET 128 = rw2.n1 
* NET 129 = rw3.n1 
* NET 130 = rw1.n1 
* NET 131 = rw0.n1 
* NET 132 = rc116.n2 
* NET 143 = rp4/15.s3 
* NET 144 = rmx4/15.bl0_p 
* NET 145 = rp4/14.s2 
* NET 146 = rp4/14.s1 
* NET 147 = rp4/15.s2 
* NET 148 = rp4/15.s1 
* NET 149 = rp4/14.s3 
* NET 150 = rmx4/14.bl0_p 
* NET 151 = rp4/13.s3 
* NET 152 = rmx4/13.bl0_p 
* NET 153 = rp4/12.s2 
* NET 154 = rp4/13.s2 
* NET 155 = rp4/12.s3 
* NET 156 = rp4/12.s1 
* NET 157 = rp4/13.s1 
* NET 158 = rp4/11.s3 
* NET 159 = rmx4/11.bl0_p 
* NET 160 = rp4/11.s2 
* NET 161 = rp4/11.s1 
* NET 162 = rmx4/12.bl0_p 
* NET 163 = rp4/10.s2 
* NET 164 = rp4/10.s3 
* NET 165 = rp4/10.s1 
* NET 166 = rmx4/10.bl0_p 
* NET 167 = rp4/9.s3 
* NET 168 = rmx4/9.bl0_p 
* NET 169 = rp4/9.s2 
* NET 170 = rp4/9.s1 
* NET 171 = rmx4/7.bl0_p 
* NET 172 = rp4/7.s3 
* NET 173 = rp4/8.s3 
* NET 174 = rmx4/8.bl0_p 
* NET 175 = rp4/8.s2 
* NET 176 = rp4/8.s1 
* NET 177 = rp4/6.s2 
* NET 178 = rp4/6.s1 
* NET 179 = rp4/7.s2 
* NET 180 = rp4/7.s1 
* NET 181 = rp4/5.s3 
* NET 182 = rmx4/5.bl0_p 
* NET 183 = rp4/6.s3 
* NET 184 = rmx4/6.bl0_p 
* NET 185 = rp4/4.s2 
* NET 186 = rp4/4.s1 
* NET 187 = rp4/5.s2 
* NET 188 = rp4/5.s1 
* NET 189 = rp4/3.s2 
* NET 190 = rp4/3.s3 
* NET 191 = rp4/3.s1 
* NET 192 = rmx4/3.bl0_p 
* NET 193 = rp4/4.s3 
* NET 194 = rmx4/4.bl0_p 
* NET 195 = rp4/2.s2 
* NET 196 = rp4/2.s3 
* NET 197 = rp4/2.s1 
* NET 198 = rmx4/2.bl0_p 
* NET 199 = rp4/1.s2 
* NET 200 = rp4/1.s3 
* NET 201 = rp4/1.s1 
* NET 202 = rmx4/1.bl0_p 
* NET 203 = x0.w2 
* NET 204 = x0.w1 
* NET 205 = x0.w0 
* NET 206 = rp4/0.s2 
* NET 207 = rp4/0.s3 
* NET 208 = rp4/0.s1 
* NET 209 = rmx4/0.bl0_p 
* NET 210 = ck[0] 
* NET 217 = rw1.inv 
* NET 220 = x2.ck_11 
* NET 222 = x1.w3 
* NET 223 = rmx4/15.bit_p 
* NET 224 = rmx4/14.bit_p 
* NET 225 = rmx4/13.bit_p 
* NET 226 = rmx4/12.bit_p 
* NET 227 = rmx4/11.bit_p 
* NET 228 = rmx4/10.bit_p 
* NET 229 = rmx4/9.bit_p 
* NET 230 = rmx4/8.bit_p 
* NET 231 = rmx4/7.bit_p 
* NET 232 = rmx4/6.bit_p 
* NET 233 = rmx4/5.bit_p 
* NET 234 = rmx4/4.bit_p 
* NET 235 = rmx4/3.bit_p 
* NET 236 = rmx4/2.bit_p 
* NET 237 = rmx4/1.bit_p 
* NET 238 = x1.ck_13 
* NET 239 = rmx4/0.bit_p 
* NET 242 = x2.n3b 
* NET 244 = rmx2/7.i1 
* NET 246 = rmx2/7.i0 
* NET 248 = rmx2/7.s_p 
* NET 252 = rmx2/6.s_p 
* NET 254 = rmx2/5.i1 
* NET 257 = rmx2/5.i0 
* NET 258 = rmx2/5.s_p 
* NET 260 = rmx2/3.i1 
* NET 265 = rmx2/4.s_p 
* NET 266 = rmx2/3.i0 
* NET 268 = rmx2/3.s_p 
* NET 273 = rmx2/1.i1 
* NET 274 = rmx2/2.s_p 
* NET 277 = rmx2/1.i0 
* NET 278 = rmx2/1.s_p 
* NET 281 = bf.e1 
* NET 282 = bf.e0 
* NET 284 = rmx2/0.s_p 
* NET 294 = adr[7] 
* NET 295 = rli/0.f 
* NET 296 = adr[4] 
* NET 297 = adr[5] 
* NET 298 = adr[6] 
* NET 299 = rw3.e1 
* NET 300 = rli/2.f 
* NET 301 = rli/1.f 
* NET 302 = adr[1] 
* NET 303 = adr[2] 
* NET 304 = adr[3] 
* NET 305 = x1.s5 
* NET 306 = x2.s0 
* NET 307 = rw3.e3 
* NET 308 = adr[0] 
* NET 309 = x0.s7 
* NET 310 = rob/7.vss1 
* NET 311 = f[7] 
* NET 312 = rob/6.vss1 
* NET 313 = f[6] 
* NET 314 = rob/5.vss1 
* NET 315 = f[5] 
* NET 316 = rob/4.vss1 
* NET 317 = f[4] 
* NET 318 = rob/3.vss1 
* NET 319 = f[3] 
* NET 320 = rob/2.vss1 
* NET 321 = f[2] 
* NET 322 = rob/1.vss1 
* NET 323 = f[1] 
* NET 324 = vdd 
* NET 325 = rob/0.vss1 
* NET 326 = f[0] 
* NET 327 = vss 
Mtr_02885 2 1 324 324 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02884 115 2 324 324 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02883 324 2 115 324 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02882 115 2 324 324 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02881 324 115 121 324 tp L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02880 324 121 3 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02879 324 3 4 324 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02878 7 4 324 324 tp L=1U W=54U AS=108P AD=108P PS=112U PD=112U 
Mtr_02877 11 294 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02876 324 11 9 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02875 11 297 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02874 8 327 13 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02873 9 115 8 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02872 324 298 11 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02871 14 121 324 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02870 324 5 6 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02869 18 15 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02868 18 15 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02867 324 6 5 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02866 15 18 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02865 324 121 5 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02864 15 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02863 324 16 19 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02862 20 17 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02861 324 16 19 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02860 20 17 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02859 324 121 16 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02858 17 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02857 17 20 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02856 324 19 16 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02855 324 5 6 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02854 25 294 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02853 324 25 22 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02852 25 300 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02851 21 327 26 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02850 22 115 21 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02849 324 298 25 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02848 27 121 324 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02847 324 28 34 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02846 35 29 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02845 35 29 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02844 324 34 28 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02843 29 35 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02842 324 121 28 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02841 29 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02840 324 30 33 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02839 32 31 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02838 324 30 33 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02837 32 31 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02836 324 121 30 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02835 31 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02834 31 32 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02833 324 33 30 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02832 324 28 34 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02831 49 294 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02830 324 49 37 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02829 49 297 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02828 36 327 50 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02827 37 115 36 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02826 324 301 49 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02825 51 121 324 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02824 324 40 44 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02823 45 41 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02822 45 41 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02821 324 44 40 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02820 41 45 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02819 324 121 40 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02818 41 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02817 324 42 43 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02816 55 52 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02815 324 42 43 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02814 55 52 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02813 324 121 42 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02812 52 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02811 52 55 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02810 324 43 42 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02809 324 40 44 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02808 61 294 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02807 324 61 47 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02806 61 300 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02805 46 327 63 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02804 47 115 46 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02803 324 301 61 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02802 64 121 324 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02801 324 53 58 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02800 57 54 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02799 57 54 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02798 324 58 53 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02797 54 57 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02796 324 121 53 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02795 54 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02794 324 65 56 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02793 70 66 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02792 324 65 56 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02791 70 66 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02790 324 121 65 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02789 66 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02788 66 70 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02787 324 56 65 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02786 324 53 58 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02785 74 295 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02784 324 74 60 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02783 74 297 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02782 59 327 77 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02781 60 115 59 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02780 324 298 74 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02779 78 121 324 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02778 324 67 69 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02777 71 68 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02776 71 68 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02775 324 69 67 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02774 68 71 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02773 324 121 67 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02772 68 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02771 324 79 83 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02770 86 80 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02769 324 79 83 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02768 86 80 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02767 324 121 79 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02766 80 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02765 80 86 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02764 324 83 79 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02763 324 67 69 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02762 89 295 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02761 324 89 72 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02760 89 300 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02759 73 327 92 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02758 72 115 73 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02757 324 298 89 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02756 93 121 324 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02755 324 81 85 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02754 84 82 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02753 84 82 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02752 324 85 81 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02751 82 84 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02750 324 121 81 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02749 82 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02748 324 94 99 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02747 98 95 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02746 324 94 99 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02745 98 95 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02744 324 121 94 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02743 95 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02742 95 98 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02741 324 99 94 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02740 324 81 85 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02739 100 295 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02738 324 100 87 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02737 100 297 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02736 88 327 103 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02735 87 115 88 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02734 324 301 100 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02733 104 121 324 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02732 324 96 97 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02731 109 105 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02730 109 105 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02729 324 97 96 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02728 105 109 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02727 324 121 96 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02726 105 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02725 324 106 112 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02724 111 107 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02723 324 106 112 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02722 111 107 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02721 324 121 106 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02720 107 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02719 107 111 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02718 324 112 106 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02717 324 96 97 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02716 118 295 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02715 324 118 114 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02714 118 300 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02713 113 327 119 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02712 114 115 113 324 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_02711 324 301 118 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02710 120 121 324 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02709 324 108 110 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02708 126 122 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02707 126 122 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02706 324 110 108 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02705 122 126 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02704 324 121 108 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02703 122 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02702 324 123 125 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02701 127 124 324 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02700 324 123 125 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02699 127 124 324 324 tp L=1U W=45U AS=90P AD=90P PS=94U PD=94U 
Mtr_02698 324 121 123 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02697 124 121 324 324 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02696 124 127 324 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02695 324 125 123 324 tp L=2U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02694 324 108 110 324 tp L=1U W=46U AS=92P AD=92P PS=96U PD=96U 
Mtr_02693 220 210 324 324 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02692 324 212 129 324 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02691 129 212 324 324 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02690 212 296 324 324 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02689 324 304 212 324 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02688 324 213 128 324 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02687 128 213 324 324 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02686 324 296 213 324 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02685 213 307 324 324 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02684 324 217 130 324 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02683 130 217 324 324 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02682 217 299 324 324 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02681 324 304 217 324 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02680 324 218 131 324 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02679 131 218 324 324 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_02678 324 299 218 324 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02677 218 307 324 324 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02676 324 220 132 324 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02675 238 132 324 324 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02674 324 132 238 324 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02673 238 132 324 324 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02672 324 132 238 324 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02671 324 142 205 324 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02670 204 141 324 324 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02669 324 220 141 324 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02668 141 309 324 324 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02667 324 302 141 324 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02666 142 308 324 324 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02665 324 302 142 324 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02664 324 220 142 324 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02663 324 219 203 324 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02662 222 221 324 324 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02661 219 220 324 324 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02660 219 308 324 324 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02659 221 220 324 324 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02658 324 305 221 324 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02657 221 309 324 324 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02656 324 305 219 324 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02655 324 306 242 324 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02654 242 220 324 324 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02653 324 303 243 324 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02652 243 220 324 324 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02651 282 242 324 324 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02650 324 243 281 324 tp L=1U W=34U AS=68P AD=68P PS=72U PD=72U 
Mtr_02649 223 244 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02648 324 238 223 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02647 324 223 244 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02646 224 246 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02645 324 238 224 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02644 324 224 246 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02643 225 249 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02642 324 238 225 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02641 324 225 249 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02640 226 250 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02639 324 238 226 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02638 324 226 250 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02637 227 254 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02636 324 238 227 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02635 324 227 254 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02634 228 257 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02633 324 238 228 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02632 324 228 257 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02631 229 259 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02630 324 238 229 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02629 324 229 259 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02628 230 261 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02627 324 238 230 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02626 324 230 261 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02625 231 260 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02624 324 238 231 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02623 324 231 260 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02622 232 266 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02621 324 238 232 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02620 324 232 266 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02619 233 269 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02618 324 238 233 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02617 324 233 269 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02616 234 270 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02615 324 238 234 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02614 324 234 270 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02613 235 273 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02612 324 238 235 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02611 324 235 273 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02610 236 277 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02609 324 238 236 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02608 324 236 277 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02607 237 279 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02606 324 238 237 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02605 324 237 279 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02604 239 280 324 324 tp L=4U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02603 324 238 239 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02602 324 239 280 324 tp L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02601 324 294 295 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02600 295 294 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02599 295 294 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02598 324 294 295 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02597 295 294 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02596 295 294 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02595 324 298 301 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02594 301 298 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02593 301 298 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02592 324 298 301 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02591 301 298 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02590 301 298 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02589 324 297 300 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02588 300 297 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02587 300 297 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02586 324 297 300 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02585 300 297 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02584 300 297 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02583 324 296 299 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02582 299 296 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02581 299 296 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02580 324 296 299 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02579 299 296 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02578 299 296 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02577 324 304 307 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02576 307 304 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02575 307 304 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02574 324 304 307 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02573 307 304 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02572 307 304 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02571 324 303 306 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02570 306 303 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02569 306 303 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02568 324 303 306 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02567 306 303 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02566 306 303 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02565 324 302 305 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02564 305 302 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02563 305 302 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02562 324 302 305 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02561 305 302 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02560 305 302 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02559 324 308 309 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02558 309 308 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02557 309 308 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02556 324 308 309 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02555 309 308 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02554 309 308 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02553 248 238 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02552 248 286 324 324 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02551 286 248 324 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02550 324 248 286 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02549 324 310 311 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02548 311 310 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02547 324 310 311 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02546 324 310 311 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02545 311 310 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02544 324 310 311 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02543 324 286 310 324 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02542 252 238 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02541 252 287 324 324 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02540 287 252 324 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02539 324 252 287 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02538 324 312 313 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02537 313 312 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02536 324 312 313 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02535 324 312 313 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02534 313 312 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02533 324 312 313 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02532 324 287 312 324 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02531 258 238 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02530 258 288 324 324 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02529 288 258 324 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02528 324 258 288 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02527 324 314 315 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02526 315 314 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02525 324 314 315 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02524 324 314 315 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02523 315 314 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02522 324 314 315 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02521 324 288 314 324 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02520 265 238 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02519 265 289 324 324 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02518 289 265 324 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02517 324 265 289 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02516 324 316 317 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02515 317 316 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02514 324 316 317 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02513 324 316 317 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02512 317 316 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02511 324 316 317 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02510 324 289 316 324 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02509 268 238 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02508 268 290 324 324 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02507 290 268 324 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02506 324 268 290 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02505 324 318 319 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02504 319 318 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02503 324 318 319 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02502 324 318 319 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02501 319 318 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02500 324 318 319 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02499 324 290 318 324 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02498 274 238 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02497 274 291 324 324 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02496 291 274 324 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02495 324 274 291 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02494 324 320 321 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02493 321 320 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02492 324 320 321 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02491 324 320 321 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02490 321 320 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02489 324 320 321 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02488 324 291 320 324 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02487 278 238 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02486 278 292 324 324 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02485 292 278 324 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02484 324 278 292 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02483 324 322 323 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02482 323 322 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02481 324 322 323 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02480 324 322 323 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02479 323 322 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02478 324 322 323 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02477 324 292 322 324 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02476 284 238 324 324 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02475 284 293 324 324 tp L=3U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_02474 293 284 324 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02473 324 284 293 324 tp L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02472 324 325 326 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02471 326 325 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02470 324 325 326 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02469 324 325 326 324 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02468 326 325 324 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02467 324 325 326 324 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02466 324 293 325 324 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02465 2 1 327 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02464 115 2 327 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02463 327 2 115 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02462 327 121 3 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02461 121 115 327 327 tn L=1U W=18U AS=36P AD=36P PS=40U PD=40U 
Mtr_02460 327 3 4 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02459 7 4 327 327 tn L=1U W=28U AS=56P AD=56P PS=60U PD=60U 
Mtr_02458 327 327 13 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02457 11 297 10 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02456 10 298 12 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02455 12 294 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02454 327 11 13 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02453 13 115 327 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02452 14 129 5 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02451 15 128 14 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02450 14 130 16 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02449 17 131 14 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02448 327 13 14 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02447 14 13 327 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02446 327 5 6 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02445 18 15 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02444 327 16 19 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02443 20 17 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02442 327 327 26 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02441 25 300 23 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02440 23 298 24 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02439 24 294 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02438 327 25 26 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02437 26 115 327 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02436 27 129 28 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02435 29 128 27 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02434 27 130 30 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02433 31 131 27 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02432 327 26 27 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02431 27 26 327 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02430 327 28 34 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02429 35 29 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02428 327 30 33 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02427 32 31 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02426 327 327 50 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02425 49 297 39 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02424 39 301 38 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02423 38 294 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02422 327 49 50 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02421 50 115 327 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02420 51 129 40 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02419 41 128 51 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02418 51 130 42 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02417 52 131 51 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02416 327 50 51 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02415 51 50 327 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02414 327 40 44 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02413 45 41 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02412 327 42 43 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02411 55 52 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02410 327 327 63 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02409 61 300 62 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02408 62 301 48 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02407 48 294 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02406 327 61 63 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02405 63 115 327 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02404 64 129 53 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02403 54 128 64 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02402 64 130 65 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02401 66 131 64 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02400 327 63 64 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02399 64 63 327 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02398 327 53 58 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02397 57 54 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02396 327 65 56 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02395 70 66 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02394 327 327 77 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02393 74 297 75 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02392 75 298 76 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02391 76 295 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02390 327 74 77 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02389 77 115 327 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02388 78 129 67 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02387 68 128 78 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02386 78 130 79 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02385 80 131 78 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02384 327 77 78 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02383 78 77 327 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02382 327 67 69 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02381 71 68 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02380 327 79 83 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02379 86 80 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02378 327 327 92 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02377 89 300 91 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02376 91 298 90 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02375 90 295 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02374 327 89 92 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02373 92 115 327 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02372 93 129 81 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02371 82 128 93 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02370 93 130 94 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02369 95 131 93 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02368 327 92 93 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02367 93 92 327 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02366 327 81 85 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02365 84 82 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02364 327 94 99 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02363 98 95 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02362 327 327 103 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02361 100 297 101 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02360 101 301 102 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02359 102 295 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02358 327 100 103 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02357 103 115 327 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02356 104 129 96 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02355 105 128 104 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02354 104 130 106 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02353 107 131 104 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02352 327 103 104 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02351 104 103 327 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02350 327 96 97 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02349 109 105 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02348 327 106 112 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02347 111 107 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02346 327 327 119 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02345 118 300 116 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02344 116 301 117 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02343 117 295 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02342 327 118 119 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02341 119 115 327 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02340 120 129 108 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02339 122 128 120 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02338 120 130 123 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02337 124 131 120 327 tn L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02336 327 119 120 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02335 120 119 327 327 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02334 327 108 110 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02333 126 122 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02332 327 123 125 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02331 127 124 327 327 tn L=1U W=36U AS=72P AD=72P PS=76U PD=76U 
Mtr_02330 327 210 220 327 tn L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_02329 129 212 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02328 327 212 129 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02327 212 304 211 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02326 211 296 327 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02325 128 213 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02324 327 213 128 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02323 214 307 213 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02322 327 296 214 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02321 130 217 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02320 327 217 130 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02319 216 299 327 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02318 217 304 216 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02317 327 218 131 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02316 215 307 218 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02315 327 299 215 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02314 131 218 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02313 132 220 327 327 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02312 327 132 238 327 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_02311 238 132 327 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02310 139 220 141 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02309 140 309 139 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02308 327 302 140 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02307 204 141 327 327 tn L=1U W=26U AS=52P AD=52P PS=56U PD=56U 
Mtr_02306 137 220 142 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02305 138 308 137 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02304 327 302 138 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02303 327 142 205 327 tn L=1U W=26U AS=52P AD=52P PS=56U PD=56U 
Mtr_02302 135 220 327 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02301 136 305 135 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02300 219 308 136 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02299 327 219 203 327 tn L=1U W=26U AS=52P AD=52P PS=56U PD=56U 
Mtr_02298 222 221 327 327 tn L=1U W=26U AS=52P AD=52P PS=56U PD=56U 
Mtr_02297 133 220 327 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02296 134 305 133 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02295 221 309 134 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02294 242 306 240 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02293 240 220 327 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02292 282 242 327 327 tn L=1U W=18U AS=36P AD=36P PS=40U PD=40U 
Mtr_02291 327 243 281 327 tn L=1U W=18U AS=36P AD=36P PS=40U PD=40U 
Mtr_02290 243 303 241 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02289 241 220 327 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02288 144 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02287 143 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02286 147 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02285 148 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02284 148 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02283 147 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02282 327 34 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02281 327 34 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02280 148 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02279 147 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02278 327 19 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02277 327 19 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02276 327 6 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02275 327 6 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02274 148 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02273 147 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02272 143 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02271 327 34 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02270 143 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02269 327 19 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02268 143 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02267 327 6 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02266 144 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02265 327 34 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02264 144 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02263 327 19 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02262 144 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02261 327 6 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02260 148 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02259 147 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02258 327 44 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02257 327 44 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02256 147 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02255 148 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02254 327 33 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02253 327 33 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02252 327 33 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02251 143 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02250 327 44 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02249 143 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02248 327 33 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02247 144 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02246 327 44 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02245 144 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02244 327 43 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02243 327 43 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02242 148 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02241 147 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02240 327 43 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02239 327 43 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02238 143 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02237 144 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02236 327 58 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02235 327 58 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02234 327 58 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02233 327 58 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02232 148 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02231 147 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02230 143 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02229 144 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02228 148 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02227 327 56 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02226 147 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02225 327 56 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02224 143 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02223 327 56 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02222 327 56 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02221 144 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02220 148 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02219 147 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02218 327 85 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02217 327 85 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02216 148 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02215 147 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02214 327 83 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02213 327 83 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02212 327 69 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02211 327 69 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02210 148 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02209 147 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02208 143 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02207 327 85 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02206 143 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02205 327 83 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02204 143 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02203 327 69 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02202 144 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02201 327 85 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02200 144 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02199 327 83 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02198 144 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02197 327 69 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02196 148 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02195 147 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02194 327 97 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02193 327 97 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02192 147 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02191 148 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02190 327 99 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02189 327 99 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02188 327 99 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02187 143 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02186 327 97 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02185 143 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02184 327 99 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02183 144 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02182 327 97 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02181 144 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02180 327 112 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02179 327 112 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02178 148 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02177 147 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02176 327 112 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02175 327 112 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02174 143 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02173 144 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02172 327 110 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02171 327 110 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02170 327 110 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02169 327 110 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02168 148 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02167 147 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02166 143 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02165 144 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02164 148 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02163 327 125 148 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02162 147 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02161 327 125 147 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02160 143 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02159 327 125 143 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02158 327 125 144 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02157 144 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02156 223 205 144 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02155 327 223 244 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02154 147 203 223 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02153 223 222 148 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02152 223 204 143 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02151 150 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02150 149 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02149 145 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02148 146 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02147 146 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02146 145 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02145 327 34 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02144 327 34 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02143 146 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02142 145 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02141 327 19 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02140 327 19 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02139 327 6 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02138 327 6 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02137 146 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02136 145 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02135 149 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02134 327 34 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02133 149 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02132 327 19 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02131 149 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02130 327 6 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02129 150 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02128 327 34 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02127 150 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02126 327 19 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02125 150 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02124 327 6 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02123 146 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02122 145 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02121 327 44 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02120 327 44 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02119 145 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02118 146 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02117 327 33 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02116 327 33 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02115 327 33 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02114 149 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02113 327 44 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02112 149 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02111 327 33 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02110 150 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02109 327 44 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02108 150 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02107 327 43 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02106 327 43 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02105 146 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02104 145 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02103 327 43 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02102 327 43 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02101 149 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02100 150 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02099 327 58 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02098 327 58 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02097 327 58 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02096 327 58 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02095 146 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02094 145 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02093 149 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02092 150 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02091 146 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02090 327 56 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02089 145 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02088 327 56 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02087 149 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02086 327 56 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02085 327 56 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02084 150 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02083 146 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02082 145 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02081 327 85 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02080 327 85 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02079 146 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02078 145 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02077 327 83 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02076 327 83 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02075 327 69 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02074 327 69 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02073 146 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02072 145 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02071 149 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02070 327 85 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02069 149 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02068 327 83 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02067 149 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02066 327 69 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02065 150 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02064 327 85 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02063 150 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02062 327 83 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02061 150 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02060 327 69 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02059 146 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02058 145 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02057 327 97 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02056 327 97 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02055 145 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02054 146 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02053 327 99 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02052 327 99 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02051 327 99 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02050 149 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02049 327 97 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02048 149 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02047 327 99 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02046 150 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02045 327 97 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02044 150 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02043 327 112 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02042 327 112 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02041 146 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02040 145 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02039 327 112 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02038 327 112 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02037 149 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02036 150 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02035 327 110 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02034 327 110 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02033 327 110 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02032 327 110 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02031 146 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02030 145 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02029 149 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02028 150 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02027 146 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02026 327 125 146 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02025 145 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02024 327 125 145 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02023 149 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02022 327 125 149 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02021 327 125 150 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02020 150 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02019 224 205 150 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02018 327 224 246 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_02017 145 203 224 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02016 224 222 146 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02015 224 204 149 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02014 152 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02013 151 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02012 154 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02011 157 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02010 157 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02009 154 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02008 327 34 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02007 327 34 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02006 157 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02005 154 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02004 327 19 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02003 327 19 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02002 327 6 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02001 327 6 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02000 157 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01999 154 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01998 151 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01997 327 34 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01996 151 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01995 327 19 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01994 151 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01993 327 6 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01992 152 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01991 327 34 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01990 152 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01989 327 19 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01988 152 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01987 327 6 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01986 157 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01985 154 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01984 327 44 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01983 327 44 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01982 154 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01981 157 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01980 327 33 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01979 327 33 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01978 327 33 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01977 151 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01976 327 44 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01975 151 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01974 327 33 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01973 152 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01972 327 44 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01971 152 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01970 327 43 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01969 327 43 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01968 157 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01967 154 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01966 327 43 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01965 327 43 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01964 151 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01963 152 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01962 327 58 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01961 327 58 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01960 327 58 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01959 327 58 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01958 157 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01957 154 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01956 151 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01955 152 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01954 157 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01953 327 56 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01952 154 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01951 327 56 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01950 151 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01949 327 56 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01948 327 56 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01947 152 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01946 157 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01945 154 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01944 327 85 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01943 327 85 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01942 157 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01941 154 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01940 327 83 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01939 327 83 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01938 327 69 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01937 327 69 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01936 157 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01935 154 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01934 151 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01933 327 85 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01932 151 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01931 327 83 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01930 151 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01929 327 69 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01928 152 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01927 327 85 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01926 152 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01925 327 83 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01924 152 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01923 327 69 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01922 157 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01921 154 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01920 327 97 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01919 327 97 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01918 154 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01917 157 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01916 327 99 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01915 327 99 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01914 327 99 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01913 151 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01912 327 97 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01911 151 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01910 327 99 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01909 152 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01908 327 97 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01907 152 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01906 327 112 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01905 327 112 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01904 157 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01903 154 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01902 327 112 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01901 327 112 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01900 151 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01899 152 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01898 327 110 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01897 327 110 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01896 327 110 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01895 327 110 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01894 157 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01893 154 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01892 151 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01891 152 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01890 157 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01889 327 125 157 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01888 154 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01887 327 125 154 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01886 151 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01885 327 125 151 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01884 327 125 152 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01883 152 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01882 225 205 152 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01881 327 225 249 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01880 154 203 225 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01879 225 222 157 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01878 225 204 151 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01877 162 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01876 155 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01875 153 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01874 156 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01873 156 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01872 153 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01871 327 34 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01870 327 34 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01869 156 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01868 153 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01867 327 19 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01866 327 19 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01865 327 6 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01864 327 6 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01863 156 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01862 153 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01861 155 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01860 327 34 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01859 155 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01858 327 19 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01857 155 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01856 327 6 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01855 162 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01854 327 34 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01853 162 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01852 327 19 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01851 162 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01850 327 6 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01849 156 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01848 153 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01847 327 44 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01846 327 44 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01845 153 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01844 156 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01843 327 33 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01842 327 33 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01841 327 33 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01840 155 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01839 327 44 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01838 155 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01837 327 33 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01836 162 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01835 327 44 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01834 162 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01833 327 43 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01832 327 43 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01831 156 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01830 153 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01829 327 43 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01828 327 43 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01827 155 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01826 162 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01825 327 58 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01824 327 58 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01823 327 58 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01822 327 58 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01821 156 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01820 153 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01819 155 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01818 162 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01817 156 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01816 327 56 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01815 153 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01814 327 56 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01813 155 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01812 327 56 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01811 327 56 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01810 162 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01809 156 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01808 153 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01807 327 85 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01806 327 85 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01805 156 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01804 153 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01803 327 83 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01802 327 83 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01801 327 69 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01800 327 69 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01799 156 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01798 153 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01797 155 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01796 327 85 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01795 155 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01794 327 83 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01793 155 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01792 327 69 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01791 162 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01790 327 85 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01789 162 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01788 327 83 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01787 162 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01786 327 69 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01785 156 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01784 153 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01783 327 97 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01782 327 97 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01781 153 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01780 156 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01779 327 99 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01778 327 99 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01777 327 99 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01776 155 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01775 327 97 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01774 155 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01773 327 99 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01772 162 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01771 327 97 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01770 162 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01769 327 112 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01768 327 112 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01767 156 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01766 153 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01765 327 112 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01764 327 112 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01763 155 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01762 162 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01761 327 110 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01760 327 110 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01759 327 110 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01758 327 110 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01757 156 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01756 153 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01755 155 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01754 162 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01753 156 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01752 327 125 156 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01751 153 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01750 327 125 153 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01749 155 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01748 327 125 155 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01747 327 125 162 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01746 162 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01745 226 205 162 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01744 327 226 250 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01743 153 203 226 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01742 226 222 156 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01741 226 204 155 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01740 159 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01739 158 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01738 160 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01737 161 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01736 161 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01735 160 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01734 327 34 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01733 327 34 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01732 161 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01731 160 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01730 327 19 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01729 327 19 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01728 327 6 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01727 327 6 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01726 161 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01725 160 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01724 158 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01723 327 34 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01722 158 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01721 327 19 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01720 158 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01719 327 6 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01718 159 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01717 327 34 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01716 159 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01715 327 19 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01714 159 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01713 327 6 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01712 161 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01711 160 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01710 327 44 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01709 327 44 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01708 160 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01707 161 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01706 327 33 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01705 327 33 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01704 327 33 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01703 158 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01702 327 44 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01701 158 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01700 327 33 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01699 159 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01698 327 44 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01697 159 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01696 327 43 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01695 327 43 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01694 161 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01693 160 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01692 327 43 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01691 327 43 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01690 158 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01689 159 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01688 327 58 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01687 327 58 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01686 327 58 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01685 327 58 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01684 161 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01683 160 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01682 158 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01681 159 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01680 161 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01679 327 56 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01678 160 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01677 327 56 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01676 158 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01675 327 56 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01674 327 56 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01673 159 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01672 161 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01671 160 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01670 327 85 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01669 327 85 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01668 161 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01667 160 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01666 327 83 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01665 327 83 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01664 327 69 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01663 327 69 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01662 161 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01661 160 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01660 158 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01659 327 85 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01658 158 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01657 327 83 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01656 158 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01655 327 69 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01654 159 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01653 327 85 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01652 159 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01651 327 83 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01650 159 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01649 327 69 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01648 161 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01647 160 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01646 327 97 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01645 327 97 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01644 160 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01643 161 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01642 327 99 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01641 327 99 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01640 327 99 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01639 158 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01638 327 97 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01637 158 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01636 327 99 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01635 159 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01634 327 97 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01633 159 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01632 327 112 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01631 327 112 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01630 161 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01629 160 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01628 327 112 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01627 327 112 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01626 158 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01625 159 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01624 327 110 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01623 327 110 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01622 327 110 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01621 327 110 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01620 161 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01619 160 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01618 158 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01617 159 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01616 161 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01615 327 125 161 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01614 160 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01613 327 125 160 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01612 158 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01611 327 125 158 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01610 327 125 159 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01609 159 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01608 227 205 159 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01607 327 227 254 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01606 160 203 227 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01605 227 222 161 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01604 227 204 158 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01603 166 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01602 164 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01601 163 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01600 165 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01599 165 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01598 163 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01597 327 34 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01596 327 34 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01595 165 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01594 163 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01593 327 19 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01592 327 19 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01591 327 6 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01590 327 6 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01589 165 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01588 163 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01587 164 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01586 327 34 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01585 164 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01584 327 19 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01583 164 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01582 327 6 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01581 166 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01580 327 34 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01579 166 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01578 327 19 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01577 166 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01576 327 6 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01575 165 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01574 163 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01573 327 44 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01572 327 44 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01571 163 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01570 165 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01569 327 33 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01568 327 33 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01567 327 33 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01566 164 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01565 327 44 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01564 164 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01563 327 33 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01562 166 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01561 327 44 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01560 166 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01559 327 43 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01558 327 43 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01557 165 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01556 163 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01555 327 43 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01554 327 43 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01553 164 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01552 166 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01551 327 58 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01550 327 58 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01549 327 58 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01548 327 58 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01547 165 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01546 163 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01545 164 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01544 166 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01543 165 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01542 327 56 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01541 163 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01540 327 56 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01539 164 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01538 327 56 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01537 327 56 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01536 166 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01535 165 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01534 163 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01533 327 85 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01532 327 85 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01531 165 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01530 163 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01529 327 83 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01528 327 83 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01527 327 69 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01526 327 69 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01525 165 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01524 163 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01523 164 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01522 327 85 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01521 164 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01520 327 83 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01519 164 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01518 327 69 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01517 166 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01516 327 85 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01515 166 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01514 327 83 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01513 166 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01512 327 69 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01511 165 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01510 163 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01509 327 97 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01508 327 97 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01507 163 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01506 165 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01505 327 99 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01504 327 99 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01503 327 99 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01502 164 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01501 327 97 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01500 164 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01499 327 99 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01498 166 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01497 327 97 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01496 166 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01495 327 112 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01494 327 112 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01493 165 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01492 163 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01491 327 112 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01490 327 112 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01489 164 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01488 166 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01487 327 110 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01486 327 110 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01485 327 110 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01484 327 110 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01483 165 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01482 163 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01481 164 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01480 166 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01479 165 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01478 327 125 165 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01477 163 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01476 327 125 163 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01475 164 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01474 327 125 164 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01473 327 125 166 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01472 166 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01471 228 205 166 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01470 327 228 257 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01469 163 203 228 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01468 228 222 165 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01467 228 204 164 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01466 168 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01465 167 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01464 169 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01463 170 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01462 170 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01461 169 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01460 327 34 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01459 327 34 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01458 170 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01457 169 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01456 327 19 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01455 327 19 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01454 327 6 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01453 327 6 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01452 170 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01451 169 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01450 167 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01449 327 34 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01448 167 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01447 327 19 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01446 167 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01445 327 6 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01444 168 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01443 327 34 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01442 168 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01441 327 19 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01440 168 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01439 327 6 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01438 170 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01437 169 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01436 327 44 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01435 327 44 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01434 169 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01433 170 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01432 327 33 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01431 327 33 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01430 327 33 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01429 167 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01428 327 44 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01427 167 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01426 327 33 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01425 168 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01424 327 44 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01423 168 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01422 327 43 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01421 327 43 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01420 170 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01419 169 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01418 327 43 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01417 327 43 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01416 167 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01415 168 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01414 327 58 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01413 327 58 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01412 327 58 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01411 327 58 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01410 170 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01409 169 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01408 167 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01407 168 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01406 170 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01405 327 56 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01404 169 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01403 327 56 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01402 167 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01401 327 56 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01400 327 56 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01399 168 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01398 170 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01397 169 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01396 327 85 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01395 327 85 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01394 170 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01393 169 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01392 327 83 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01391 327 83 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01390 327 69 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01389 327 69 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01388 170 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01387 169 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01386 167 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01385 327 85 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01384 167 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01383 327 83 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01382 167 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01381 327 69 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01380 168 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01379 327 85 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01378 168 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01377 327 83 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01376 168 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01375 327 69 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01374 170 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01373 169 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01372 327 97 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01371 327 97 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01370 169 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01369 170 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01368 327 99 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01367 327 99 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01366 327 99 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01365 167 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01364 327 97 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01363 167 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01362 327 99 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01361 168 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01360 327 97 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01359 168 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01358 327 112 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01357 327 112 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01356 170 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01355 169 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01354 327 112 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01353 327 112 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01352 167 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01351 168 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01350 327 110 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01349 327 110 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01348 327 110 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01347 327 110 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01346 170 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01345 169 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01344 167 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01343 168 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01342 170 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01341 327 125 170 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01340 169 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01339 327 125 169 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01338 167 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01337 327 125 167 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01336 327 125 168 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01335 168 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01334 229 205 168 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01333 327 229 259 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01332 169 203 229 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01331 229 222 170 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01330 229 204 167 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01329 174 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01328 173 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01327 175 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01326 176 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01325 176 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01324 175 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01323 327 34 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01322 327 34 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01321 176 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01320 175 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01319 327 19 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01318 327 19 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01317 327 6 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01316 327 6 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01315 176 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01314 175 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01313 173 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01312 327 34 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01311 173 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01310 327 19 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01309 173 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01308 327 6 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01307 174 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01306 327 34 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01305 174 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01304 327 19 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01303 174 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01302 327 6 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01301 176 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01300 175 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01299 327 44 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01298 327 44 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01297 175 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01296 176 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01295 327 33 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01294 327 33 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01293 327 33 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01292 173 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01291 327 44 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01290 173 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01289 327 33 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01288 174 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01287 327 44 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01286 174 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01285 327 43 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01284 327 43 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01283 176 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01282 175 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01281 327 43 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01280 327 43 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01279 173 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01278 174 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01277 327 58 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01276 327 58 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01275 327 58 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01274 327 58 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01273 176 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01272 175 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01271 173 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01270 174 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01269 176 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01268 327 56 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01267 175 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01266 327 56 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01265 173 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01264 327 56 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01263 327 56 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01262 174 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01261 176 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01260 175 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01259 327 85 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01258 327 85 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01257 176 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01256 175 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01255 327 83 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01254 327 83 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01253 327 69 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01252 327 69 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01251 176 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01250 175 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01249 173 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01248 327 85 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01247 173 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01246 327 83 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01245 173 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01244 327 69 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01243 174 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01242 327 85 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01241 174 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01240 327 83 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01239 174 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01238 327 69 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01237 176 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01236 175 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01235 327 97 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01234 327 97 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01233 175 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01232 176 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01231 327 99 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01230 327 99 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01229 327 99 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01228 173 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01227 327 97 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01226 173 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01225 327 99 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01224 174 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01223 327 97 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01222 174 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01221 327 112 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01220 327 112 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01219 176 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01218 175 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01217 327 112 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01216 327 112 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01215 173 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01214 174 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01213 327 110 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01212 327 110 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01211 327 110 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01210 327 110 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01209 176 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01208 175 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01207 173 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01206 174 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01205 176 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01204 327 125 176 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01203 175 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01202 327 125 175 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01201 173 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01200 327 125 173 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01199 327 125 174 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01198 174 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01197 230 205 174 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01196 327 230 261 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01195 175 203 230 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01194 230 222 176 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01193 230 204 173 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01192 171 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01191 172 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01190 179 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01189 180 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01188 180 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01187 179 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01186 327 34 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01185 327 34 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01184 180 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01183 179 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01182 327 19 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01181 327 19 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01180 327 6 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01179 327 6 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01178 180 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01177 179 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01176 172 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01175 327 34 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01174 172 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01173 327 19 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01172 172 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01171 327 6 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01170 171 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01169 327 34 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01168 171 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01167 327 19 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01166 171 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01165 327 6 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01164 180 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01163 179 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01162 327 44 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01161 327 44 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01160 179 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01159 180 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01158 327 33 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01157 327 33 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01156 327 33 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01155 172 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01154 327 44 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01153 172 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01152 327 33 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01151 171 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01150 327 44 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01149 171 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01148 327 43 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01147 327 43 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01146 180 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01145 179 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01144 327 43 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01143 327 43 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01142 172 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01141 171 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01140 327 58 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01139 327 58 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01138 327 58 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01137 327 58 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01136 180 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01135 179 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01134 172 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01133 171 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01132 180 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01131 327 56 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01130 179 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01129 327 56 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01128 172 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01127 327 56 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01126 327 56 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01125 171 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01124 180 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01123 179 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01122 327 85 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01121 327 85 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01120 180 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01119 179 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01118 327 83 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01117 327 83 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01116 327 69 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01115 327 69 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01114 180 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01113 179 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01112 172 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01111 327 85 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01110 172 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01109 327 83 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01108 172 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01107 327 69 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01106 171 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01105 327 85 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01104 171 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01103 327 83 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01102 171 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01101 327 69 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01100 180 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01099 179 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01098 327 97 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01097 327 97 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01096 179 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01095 180 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01094 327 99 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01093 327 99 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01092 327 99 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01091 172 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01090 327 97 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01089 172 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01088 327 99 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01087 171 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01086 327 97 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01085 171 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01084 327 112 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01083 327 112 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01082 180 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01081 179 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01080 327 112 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01079 327 112 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01078 172 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01077 171 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01076 327 110 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01075 327 110 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01074 327 110 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01073 327 110 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01072 180 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01071 179 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01070 172 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01069 171 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01068 180 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01067 327 125 180 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01066 179 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01065 327 125 179 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01064 172 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01063 327 125 172 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01062 327 125 171 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01061 171 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01060 231 205 171 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01059 327 231 260 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01058 179 203 231 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01057 231 222 180 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01056 231 204 172 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01055 184 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01054 183 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01053 177 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01052 178 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01051 178 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01050 177 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01049 327 34 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01048 327 34 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01047 178 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01046 177 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01045 327 19 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01044 327 19 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01043 327 6 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01042 327 6 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01041 178 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01040 177 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01039 183 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01038 327 34 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01037 183 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01036 327 19 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01035 183 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01034 327 6 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01033 184 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01032 327 34 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01031 184 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01030 327 19 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01029 184 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01028 327 6 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01027 178 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01026 177 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01025 327 44 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01024 327 44 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01023 177 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01022 178 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01021 327 33 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01020 327 33 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01019 327 33 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01018 183 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01017 327 44 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01016 183 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01015 327 33 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01014 184 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01013 327 44 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01012 184 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01011 327 43 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01010 327 43 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01009 178 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01008 177 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01007 327 43 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01006 327 43 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01005 183 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01004 184 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01003 327 58 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01002 327 58 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01001 327 58 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01000 327 58 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00999 178 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00998 177 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00997 183 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00996 184 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00995 178 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00994 327 56 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00993 177 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00992 327 56 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00991 183 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00990 327 56 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00989 327 56 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00988 184 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00987 178 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00986 177 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00985 327 85 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00984 327 85 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00983 178 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00982 177 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00981 327 83 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00980 327 83 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00979 327 69 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00978 327 69 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00977 178 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00976 177 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00975 183 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00974 327 85 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00973 183 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00972 327 83 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00971 183 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00970 327 69 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00969 184 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00968 327 85 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00967 184 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00966 327 83 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00965 184 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00964 327 69 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00963 178 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00962 177 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00961 327 97 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00960 327 97 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00959 177 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00958 178 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00957 327 99 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00956 327 99 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00955 327 99 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00954 183 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00953 327 97 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00952 183 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00951 327 99 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00950 184 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00949 327 97 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00948 184 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00947 327 112 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00946 327 112 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00945 178 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00944 177 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00943 327 112 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00942 327 112 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00941 183 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00940 184 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00939 327 110 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00938 327 110 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00937 327 110 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00936 327 110 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00935 178 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00934 177 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00933 183 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00932 184 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00931 178 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00930 327 125 178 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00929 177 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00928 327 125 177 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00927 183 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00926 327 125 183 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00925 327 125 184 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00924 184 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00923 232 205 184 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00922 327 232 266 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00921 177 203 232 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00920 232 222 178 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00919 232 204 183 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00918 182 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00917 181 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00916 187 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00915 188 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00914 188 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00913 187 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00912 327 34 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00911 327 34 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00910 188 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00909 187 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00908 327 19 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00907 327 19 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00906 327 6 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00905 327 6 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00904 188 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00903 187 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00902 181 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00901 327 34 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00900 181 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00899 327 19 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00898 181 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00897 327 6 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00896 182 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00895 327 34 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00894 182 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00893 327 19 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00892 182 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00891 327 6 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00890 188 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00889 187 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00888 327 44 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00887 327 44 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00886 187 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00885 188 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00884 327 33 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00883 327 33 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00882 327 33 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00881 181 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00880 327 44 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00879 181 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00878 327 33 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00877 182 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00876 327 44 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00875 182 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00874 327 43 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00873 327 43 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00872 188 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00871 187 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00870 327 43 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00869 327 43 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00868 181 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00867 182 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00866 327 58 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00865 327 58 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00864 327 58 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00863 327 58 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00862 188 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00861 187 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00860 181 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00859 182 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00858 188 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00857 327 56 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00856 187 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00855 327 56 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00854 181 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00853 327 56 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00852 327 56 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00851 182 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00850 188 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00849 187 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00848 327 85 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00847 327 85 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00846 188 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00845 187 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00844 327 83 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00843 327 83 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00842 327 69 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00841 327 69 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00840 188 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00839 187 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00838 181 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00837 327 85 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00836 181 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00835 327 83 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00834 181 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00833 327 69 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00832 182 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00831 327 85 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00830 182 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00829 327 83 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00828 182 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00827 327 69 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00826 188 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00825 187 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00824 327 97 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00823 327 97 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00822 187 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00821 188 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00820 327 99 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00819 327 99 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00818 327 99 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00817 181 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00816 327 97 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00815 181 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00814 327 99 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00813 182 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00812 327 97 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00811 182 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00810 327 112 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00809 327 112 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00808 188 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00807 187 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00806 327 112 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00805 327 112 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00804 181 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00803 182 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00802 327 110 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00801 327 110 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00800 327 110 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00799 327 110 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00798 188 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00797 187 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00796 181 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00795 182 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00794 188 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00793 327 125 188 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00792 187 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00791 327 125 187 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00790 181 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00789 327 125 181 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00788 327 125 182 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00787 182 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00786 233 205 182 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00785 327 233 269 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00784 187 203 233 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00783 233 222 188 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00782 233 204 181 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00781 194 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00780 193 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00779 185 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00778 186 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00777 186 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00776 185 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00775 327 34 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00774 327 34 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00773 186 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00772 185 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00771 327 19 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00770 327 19 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00769 327 6 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00768 327 6 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00767 186 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00766 185 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00765 193 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00764 327 34 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00763 193 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00762 327 19 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00761 193 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00760 327 6 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00759 194 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00758 327 34 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00757 194 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00756 327 19 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00755 194 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00754 327 6 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00753 186 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00752 185 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00751 327 44 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00750 327 44 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00749 185 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00748 186 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00747 327 33 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00746 327 33 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00745 327 33 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00744 193 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00743 327 44 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00742 193 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00741 327 33 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00740 194 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00739 327 44 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00738 194 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00737 327 43 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00736 327 43 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00735 186 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00734 185 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00733 327 43 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00732 327 43 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00731 193 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00730 194 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00729 327 58 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00728 327 58 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00727 327 58 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00726 327 58 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00725 186 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00724 185 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00723 193 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00722 194 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00721 186 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00720 327 56 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00719 185 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00718 327 56 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00717 193 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00716 327 56 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00715 327 56 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00714 194 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00713 186 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00712 185 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00711 327 85 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00710 327 85 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00709 186 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00708 185 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00707 327 83 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00706 327 83 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00705 327 69 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00704 327 69 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00703 186 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00702 185 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00701 193 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00700 327 85 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00699 193 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00698 327 83 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00697 193 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00696 327 69 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00695 194 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00694 327 85 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00693 194 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00692 327 83 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00691 194 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00690 327 69 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00689 186 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00688 185 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00687 327 97 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00686 327 97 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00685 185 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00684 186 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00683 327 99 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00682 327 99 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00681 327 99 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00680 193 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00679 327 97 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00678 193 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00677 327 99 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00676 194 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00675 327 97 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00674 194 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00673 327 112 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00672 327 112 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00671 186 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00670 185 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00669 327 112 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00668 327 112 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00667 193 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00666 194 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00665 327 110 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00664 327 110 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00663 327 110 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00662 327 110 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00661 186 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00660 185 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00659 193 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00658 194 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00657 186 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00656 327 125 186 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00655 185 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00654 327 125 185 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00653 193 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00652 327 125 193 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00651 327 125 194 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00650 194 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00649 234 205 194 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00648 327 234 270 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00647 185 203 234 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00646 234 222 186 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00645 234 204 193 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00644 192 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00643 190 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00642 189 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00641 191 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00640 191 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00639 189 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00638 327 34 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00637 327 34 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00636 191 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00635 189 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00634 327 19 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00633 327 19 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00632 327 6 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00631 327 6 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00630 191 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00629 189 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00628 190 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00627 327 34 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00626 190 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00625 327 19 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00624 190 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00623 327 6 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00622 192 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00621 327 34 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00620 192 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00619 327 19 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00618 192 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00617 327 6 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00616 191 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00615 189 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00614 327 44 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00613 327 44 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00612 189 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00611 191 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00610 327 33 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00609 327 33 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00608 327 33 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00607 190 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00606 327 44 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00605 190 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00604 327 33 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00603 192 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00602 327 44 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00601 192 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00600 327 43 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00599 327 43 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00598 191 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00597 189 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00596 327 43 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00595 327 43 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00594 190 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00593 192 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00592 327 58 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00591 327 58 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00590 327 58 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00589 327 58 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00588 191 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00587 189 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00586 190 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00585 192 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00584 191 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00583 327 56 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00582 189 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00581 327 56 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00580 190 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00579 327 56 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00578 327 56 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00577 192 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00576 191 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00575 189 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00574 327 85 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00573 327 85 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00572 191 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00571 189 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00570 327 83 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00569 327 83 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00568 327 69 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00567 327 69 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00566 191 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00565 189 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00564 190 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00563 327 85 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00562 190 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00561 327 83 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00560 190 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00559 327 69 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00558 192 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00557 327 85 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00556 192 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00555 327 83 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00554 192 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00553 327 69 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00552 191 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00551 189 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00550 327 97 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00549 327 97 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00548 189 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00547 191 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00546 327 99 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00545 327 99 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00544 327 99 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00543 190 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00542 327 97 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00541 190 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00540 327 99 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00539 192 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00538 327 97 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00537 192 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00536 327 112 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00535 327 112 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00534 191 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00533 189 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00532 327 112 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00531 327 112 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00530 190 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00529 192 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00528 327 110 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00527 327 110 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00526 327 110 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00525 327 110 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00524 191 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00523 189 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00522 190 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00521 192 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00520 191 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00519 327 125 191 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00518 189 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00517 327 125 189 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00516 190 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00515 327 125 190 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00514 327 125 192 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00513 192 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00512 235 205 192 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00511 327 235 273 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00510 189 203 235 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00509 235 222 191 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00508 235 204 190 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00507 198 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00506 196 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00505 195 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00504 197 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00503 197 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00502 195 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00501 327 34 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00500 327 34 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00499 197 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00498 195 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00497 327 19 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00496 327 19 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00495 327 6 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00494 327 6 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00493 197 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00492 195 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00491 196 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00490 327 34 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00489 196 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00488 327 19 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00487 196 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00486 327 6 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00485 198 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00484 327 34 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00483 198 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00482 327 19 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00481 198 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00480 327 6 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00479 197 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00478 195 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00477 327 44 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00476 327 44 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00475 195 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00474 197 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00473 327 33 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00472 327 33 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00471 327 33 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00470 196 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00469 327 44 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00468 196 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00467 327 33 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00466 198 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00465 327 44 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00464 198 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00463 327 43 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00462 327 43 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00461 197 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00460 195 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00459 327 43 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00458 327 43 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00457 196 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00456 198 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00455 327 58 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00454 327 58 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00453 327 58 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00452 327 58 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00451 197 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00450 195 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00449 196 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00448 198 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00447 197 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00446 327 56 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00445 195 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00444 327 56 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00443 196 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00442 327 56 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00441 327 56 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00440 198 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00439 197 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00438 195 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00437 327 85 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00436 327 85 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00435 197 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00434 195 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00433 327 83 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00432 327 83 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00431 327 69 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00430 327 69 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00429 197 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00428 195 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00427 196 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00426 327 85 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00425 196 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00424 327 83 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00423 196 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00422 327 69 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00421 198 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00420 327 85 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00419 198 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00418 327 83 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00417 198 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00416 327 69 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00415 197 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00414 195 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00413 327 97 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00412 327 97 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00411 195 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00410 197 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00409 327 99 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00408 327 99 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00407 327 99 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00406 196 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00405 327 97 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00404 196 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00403 327 99 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00402 198 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00401 327 97 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00400 198 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00399 327 112 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00398 327 112 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00397 197 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00396 195 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00395 327 112 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00394 327 112 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00393 196 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00392 198 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00391 327 110 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00390 327 110 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00389 327 110 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00388 327 110 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00387 197 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00386 195 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00385 196 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00384 198 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00383 197 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00382 327 125 197 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00381 195 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00380 327 125 195 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00379 196 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00378 327 125 196 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00377 327 125 198 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00376 198 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00375 236 205 198 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00374 327 236 277 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00373 195 203 236 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00372 236 222 197 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00371 236 204 196 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00370 202 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00369 200 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00368 199 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00367 201 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00366 201 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00365 199 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00364 327 34 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00363 327 34 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00362 201 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00361 199 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00360 327 19 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00359 327 19 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00358 327 6 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00357 327 6 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00356 201 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00355 199 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00354 200 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00353 327 34 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00352 200 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00351 327 19 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00350 200 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00349 327 6 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00348 202 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00347 327 34 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00346 202 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00345 327 19 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00344 202 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00343 327 6 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00342 201 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00341 199 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00340 327 44 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00339 327 44 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00338 199 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00337 201 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00336 327 33 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00335 327 33 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00334 327 33 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00333 200 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00332 327 44 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00331 200 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00330 327 33 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00329 202 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00328 327 44 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00327 202 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00326 327 43 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00325 327 43 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00324 201 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00323 199 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00322 327 43 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00321 327 43 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00320 200 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00319 202 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00318 327 58 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00317 327 58 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00316 327 58 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00315 327 58 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00314 201 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00313 199 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00312 200 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00311 202 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00310 201 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00309 327 56 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00308 199 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00307 327 56 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00306 200 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00305 327 56 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00304 327 56 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00303 202 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00302 201 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00301 199 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00300 327 85 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00299 327 85 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00298 201 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00297 199 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00296 327 83 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00295 327 83 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00294 327 69 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00293 327 69 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00292 201 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00291 199 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00290 200 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00289 327 85 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00288 200 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00287 327 83 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00286 200 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00285 327 69 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00284 202 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00283 327 85 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00282 202 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00281 327 83 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00280 202 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00279 327 69 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00278 201 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00277 199 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00276 327 97 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00275 327 97 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00274 199 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00273 201 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00272 327 99 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00271 327 99 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00270 327 99 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00269 200 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00268 327 97 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00267 200 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00266 327 99 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00265 202 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00264 327 97 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00263 202 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00262 327 112 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00261 327 112 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00260 201 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00259 199 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00258 327 112 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00257 327 112 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00256 200 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00255 202 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00254 327 110 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00253 327 110 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00252 327 110 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00251 327 110 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00250 201 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00249 199 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00248 200 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00247 202 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00246 201 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00245 327 125 201 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00244 199 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00243 327 125 199 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00242 200 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00241 327 125 200 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00240 327 125 202 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00239 202 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00238 237 205 202 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00237 327 237 279 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00236 199 203 237 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00235 237 222 201 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00234 237 204 200 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00233 209 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00232 207 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00231 206 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00230 208 7 324 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00229 208 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00228 206 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00227 327 34 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00226 327 34 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00225 208 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00224 206 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00223 327 19 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00222 327 19 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00221 327 6 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00220 327 6 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00219 208 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00218 206 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00217 207 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00216 327 34 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00215 207 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00214 327 19 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00213 207 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00212 327 6 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00211 209 35 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00210 327 34 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00209 209 20 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00208 327 19 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00207 209 18 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00206 327 6 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00205 208 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00204 206 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00203 327 44 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00202 327 44 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00201 206 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00200 208 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00199 327 33 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00198 327 33 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00197 327 33 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00196 207 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00195 327 44 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00194 207 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00193 327 33 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00192 209 32 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00191 327 44 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00190 209 45 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00189 327 43 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00188 327 43 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00187 208 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00186 206 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00185 327 43 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00184 327 43 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00183 207 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00182 209 55 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00181 327 58 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00180 327 58 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00179 327 58 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00178 327 58 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00177 208 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00176 206 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00175 207 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00174 209 57 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00173 208 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00172 327 56 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00171 206 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00170 327 56 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00169 207 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00168 327 56 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00167 327 56 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00166 209 70 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00165 208 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00164 206 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00163 327 85 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00162 327 85 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00161 208 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00160 206 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00159 327 83 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00158 327 83 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00157 327 69 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00156 327 69 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00155 208 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00154 206 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00153 207 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00152 327 85 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00151 207 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00150 327 83 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00149 207 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00148 327 69 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00147 209 84 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00146 327 85 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00145 209 86 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00144 327 83 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00143 209 71 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00142 327 69 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00141 208 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00140 206 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00139 327 97 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00138 327 97 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00137 206 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00136 208 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00135 327 99 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00134 327 99 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00133 327 99 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00132 207 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00131 327 97 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00130 207 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00129 327 99 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00128 209 98 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00127 327 97 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00126 209 109 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00125 327 112 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00124 327 112 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00123 208 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00122 206 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00121 327 112 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00120 327 112 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00119 207 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00118 209 111 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00117 327 110 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00116 327 110 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00115 327 110 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00114 327 110 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00113 208 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00112 206 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00111 207 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00110 209 126 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00109 208 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00108 327 125 208 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00107 206 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00106 327 125 206 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00105 207 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00104 327 125 207 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00103 327 125 209 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00102 209 127 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00101 239 205 209 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00100 327 239 280 327 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00099 206 203 239 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00098 239 222 208 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00097 239 204 207 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00096 327 294 295 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00095 295 294 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00094 295 294 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00093 327 298 301 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00092 301 298 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00091 301 298 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00090 327 297 300 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00089 300 297 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00088 300 297 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00087 327 296 299 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00086 299 296 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00085 299 296 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00084 327 304 307 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00083 307 304 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00082 307 304 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00081 327 303 306 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00080 306 303 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00079 306 303 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00078 327 302 305 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00077 305 302 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00076 305 302 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00075 327 308 309 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00074 309 308 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00073 309 308 327 327 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00072 327 246 247 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00071 247 281 248 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00070 248 282 245 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00069 245 244 327 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00068 286 248 327 327 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00067 311 310 327 327 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00066 327 310 311 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00065 327 286 310 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00064 311 310 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00063 327 250 253 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00062 253 281 252 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00061 252 282 251 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00060 251 249 327 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00059 287 252 327 327 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00058 313 312 327 327 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00057 327 312 313 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00056 327 287 312 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00055 313 312 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00054 327 257 256 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00053 256 281 258 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00052 258 282 255 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00051 255 254 327 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00050 288 258 327 327 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00049 315 314 327 327 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00048 327 314 315 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00047 327 288 314 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00046 315 314 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00045 327 261 264 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00044 264 281 265 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00043 265 282 263 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00042 263 259 327 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00041 289 265 327 327 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00040 317 316 327 327 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00039 327 316 317 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00038 327 289 316 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00037 317 316 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00036 327 266 267 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00035 267 281 268 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00034 268 282 262 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00033 262 260 327 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00032 290 268 327 327 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00031 319 318 327 327 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00030 327 318 319 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00029 327 290 318 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00028 319 318 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00027 327 270 272 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00026 272 281 274 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00025 274 282 271 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00024 271 269 327 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00023 291 274 327 327 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00022 321 320 327 327 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00021 327 320 321 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00020 327 291 320 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00019 321 320 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00018 327 277 275 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00017 275 281 278 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00016 278 282 276 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00015 276 273 327 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00014 292 278 327 327 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00013 323 322 327 327 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00012 327 322 323 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 327 292 322 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00010 323 322 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 327 280 285 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00008 285 281 284 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00007 284 282 283 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00006 283 279 327 327 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00005 293 284 327 327 tn L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00004 326 325 327 327 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00003 327 325 326 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 327 293 325 327 tn L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00001 326 325 327 327 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
.ends r256x8_5

